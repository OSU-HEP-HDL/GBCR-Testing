

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U7hExZJod/vUi3z5N4RSr1wa48P7uP/A8O0jgaKOZBD7WNfzo6GmQd7doggkH00XJgs7nLyNvPm0
0zWCfXninQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k253ey4kkVql4FDzRxE0SZp0nnUl5fXV3ls/4mgbh/6ghGRjfZ71MsiTZ71s3tpy77tZHD0rpNoh
xUysBr1hFwWkTjAISVTsWyokKm82DELzMzaI0lqt04f7kevY+q4XugjttAECZCOOrrnUQb5ODPuL
TN/5/7rekkgE3das7WY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WoA52aV8kh0bkIXA7aISXPgNn7kpio3O4wNzPv7z4wZK/v9qsQ4Fa+1FXV0tZ0D+Si1URd5Yt8PQ
TB8Mp2LGBm7aAfzTAAqLpPZr3KRYlBsnuQptgQwkquHJi1BcDR3dhZHYw2oUKeYXBoZJ80Dg1iyE
mKNc2EAX8dBe7hH745fnWjhDqr0z4schwVFz8IHUPGI/WDdrXtDdyYzuiWdux2vjC9Gao0MkqalL
zCFAkEPTT0xtWcvaccmMU2ICHf+NVjiwhEmFT/vt1jXBw7quncqpEDMuzTHteQFztMFqsgBfXXAR
/Q4rfhaHiuQ7xUCcTEngpAsL2ypgKweMgL0LDw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yb4xLqu3x9ghRLjHN7QkYl0tDMsZMeJQgGEQuxDwwPb+acIMCaRAm0LVh6gbF0arOSlfOKBs+X6I
1sCY01AUXvqPtXEUt+RvllN5odbTYkY9f5RujZ5aQ9olezUe3+JLEML7oIeJ23v82E3q5lEn2hpd
Yirga3+XXZGIeEC2Q5F3LdU1PK/hOr/QQAn7r3cfSPSRAYJBv2q0KFRrpHEdaRVBAVRTnMADnWqM
+83djfdVuwjO+GhXELQ+rhNH9dkL0cqvHYfgIcRG0rYfPORpbXH4Uiizi44H6tpqRpTeCgmUfW/1
kW3FxovGX7M2+iedny4BJan5eJXy8iA1/NmnQw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pj6m4D23BtF6RtOvVlnmIzux1ocpf3A3ahzdQxUHuwpW9nlstiQd0oSmGGaiF66UD31sHUT6dfQd
yKhb6vxivgHto8LAAEiyTiUmNTH/c41wB3zGzcZFasAPOJZMvUysBGURofn88ip4eLF52/qIKVON
l8AKPEa6atmUOWXPGRix1yyvpjUnvxZ+wFAbBvP0ZsReS6AW7b6zRE+vUOJaMz0EaWEMMRdw3vLT
W/hp9Ruis3IsgHsdn6M611ZJnxSa2tuwXuWdXURUJzFjnTsi2R7EoD0bDJINDuh7T6iiDjBFdO8L
a4ER9/C3EG6IOxU+oP2sYgSHnI7dLthCIjJ+rw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B2bb9hbJCVaDRqGS393PhTqcBLIIS3eowUvDjLX1RVvD9vYwfdlG9rjfAUVzitJwz5TOhOabACyb
mMpxy7hxgVO56ex26Ce3uZlntRRrSfXZFQT0ENioLNV+BxEHrr7uipCant7HxRFrLFt9nR5wi4m9
ZZq5zS207DucLy0jTX0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eqzUQVv3z3gvc1IAF6D1gFpnG3jJXG9SSewyb0B7YFlkq+2WoV55oUnb7Smo54ZcwqBR15BnF2xS
jlkL+wI6xvjzAFZaDFixez8MkTdRnrNZscyGLFWOHz7RNKwEpAxAm7RSsBEcZUaS6x+lEu8Fai/i
gBi8OQLkjYbSnKt8sfNmpRhCWxhkRR0QylraXCBqvJVR8s/2S9YSm3zj5TqvYxlJahDh9O3V0iE2
aVTZ//VjzAQrgKQboTMB5R+3O0GmOfi7O8vgrOvK/PiOq6kVyAYEvce5/1FU9VRi8AQk3Hi7BRZM
1pWTxx+bC6qDX+NQvgu8HPGpHmqeqS/CQlftQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
vKbT7ICuGzWbXWktmfkEsf1KxlMboJ4t5VRrre71Y5k+tB+BzkQ7a2y1gOcKIAp7dzsPwNShBdhS
1ThVHFnFRYtN9Uy38/CrXWxXN1mIFIIB3wyW0UHeXStHU8f0lOiSDvO9nKhINFxMj9qjFFS2W2Hw
bb4Q/BPJEu8M/bE9DZvR33bIesEjE8ong3gTZS+opulPKNHJrzsw7fwpliQDnjQX9Q3u6biziqx3
2znImsgEeNhjW13voMKtEHQf8JNjnIyzotOB9b7rAn7yk2JKE+1lotanCbfEVMTpRxFusQv2W4dz
eJJ3+cKwQ1hXRndh+i3Yqi4bS0vo2n/X4+sX5UB+IF9m5Zzc9JYZS53X+Mrzpr9ZNy9cCCZJtl3c
f83hW+b9ox7MZeLz3cwdh91LRjU9RhiyZSDIbX66sdsekBMAiR2GSBleC/amA4PytT/4IBZ/N3RU
N4NMR8VUqpcyQbkso9b5Lgi8c2DjayRmxIGCGCh+IeR+1DLZxhxAEWQP3uJGwW3d2RE5GilM4H6j
E8ETbV2Mx5I22W6ceI8qPjuyQx4Et/ltFvUUJ1RaMDYFDcrJzb5q2/FGkXRLog386+Qx9ijVpXXH
pbm6dLffsbjzI6DX8JVKczYEIy5qXM5NTJm45pMvVbCT/SGIegLZm/T2JAhU0Q/1QtIsbhoQsBkH
CJGXPDoTtIGTbxyjC+rAKPaiEFKjJK/KvZOOtZtjws+E2rq80XjUJ9IOpXYi5NICJCpYR84+Cyf/
bPUY4gB1/OdUrfA1k6otAEX1Sxxvfw3Sp+I+md8LAG1QBTCeBlpYmDDvoIeO3OmtFhc2wVfMLseI
DPC072hpO0DDQbOaizhLWJ4qqm/yLFVLdKp5vdLVc6FPD/hb4sM4tOAgMjCF/3NvPKzfqIj4WfjF
d6DIwsI3KQBp3KCnsGoUK9Pa7qD005mn5IYEtSU30+n+dCmZ4NnDsWNhHBcGjDZbqYMpCkHg9aMh
jlRl53FXqPkZwpkiRR4hKDtpZQW+wFzQqwk+NmWEzV937s+1BC7BVIVycCErmymlLyBXWidCw51z
XfkWLJC65Scu5Yvnjz+foDFqvYaMrY0Pqq8NnrOVb2l6t+463Z6H57AJ2TqOxOTX6iGb40dgio5i
H3Lo6eJRdmy77UCrcP3gnMMd6NuuD0jd6uMZt+8wx5CHjAVLMgFBzP1+MYNSbReoWHuQpFWq0+7w
annAwiIryKJcXCMdi2eIMSJuOPhh0OTV2+a722YSN7ZHHP2/Fzjpgr5yw0C8nC8OQwRfJwnrUWcf
m2y0TWRyahC1x7Sk4y54DKvDZhwAtxic96j/gxC5xo6LeWOqkj6OTamU+XWUEUDMrACpMpySdQGw
0Rz/92c3q+nNRYvBjX8H9HUJmuRIjtyoYVEU2YWMUmyWfh/ZPcHaJwggmyfHZOluIK4uDf28pdZz
J4Ulg4RVLhbmn5z9sOeHRFbNkDOHkaCYaOAOY3BIIhAw0UF5BjqJL5Vov0bWvbcIQn+0B856kGBE
7hrOXbPxrM+WiXc2m7exvfnRL0Elmjz+oUlpv/f3unvGkwsKzBnn43cC+mnHQr3RBUWKmmYrjTkM
zwszqwwgOWwgjfvWQtlo243cpu7TRGGhgfe6Qet5oelVVLoLR5SwFanstEF8adtAQBXlR865Alfw
J5ELQnT2R9vZFhX0Yb/bgb5SXRFwOchmWf/x+zeVmb+WC6A7dkWaBpYvzrFSLe/OYwfS7CqveG6m
lOuIsTUdiCfjF/BJloCRLflnY8GOMBOOLVtc/ZlN+Ikf03GA70fYoOVuwvHlHNeUlwZxpPoPp89L
C1G0Ueu15trusYlIwJSLCycJnK4sKd424Ch7z08+18PmwE7A9PiPnMORCBYWhQyN5GFwrR7HV/Vn
Q38OzluOm/EoNxbu9/CMpUlB6u8X4Ncdb+XhHTPHhK7owcjFFD7rkEJ79dvfS/bGbDfsBxzWbNng
HqKhrxAQlgfpIy+jwvxIUDQXa91f4yDfL02/Dtp+qgKqO0s73glzRxpgJNe377+UVq4VyCXaVqNu
B+wWERP661DPfFfkYdCImBCtSEPFhvpTqChvmFOWVDX5U2VEI6kZQmpm0tkuKSa6XrRQQhMlRK7z
G1/uMaH1QMXZjptDVa81ntyDjud3f+F2aQtTr8BtXLVoB/lhjoatWenCRxQYB+hr/2QIQ8aE/wwo
L49sIby4IMl9gR9XdERhbuBpn+gHWF0c1Etl91wQKaTV61dMDC8iOt8OuvN+P33u7KyEUwkcZE2W
abCa+9O83UvsWykMkMy6NHE+RF50sNOWraUAlZP0Cbi87ocBVPy9IEZtLR4Bq1QgejtMUiVS8vtU
RDwXDXimti2mQmiHBsYv9TXIHlp7INKSy86pgQwLKUg95xoLdI4rUEgezPeQjtw/IPpdtw5QJSqg
ra6yyU3w6c7qc1vGY0PKmiTuKrQUQTd7EKSvXTyLFA+S2qx1+tmSwrqcdMyD7Fo2cACkpTDtFqK/
lmDNBQ3vAwgQL5i6aEKZaQLcG9Qo7SDg/CiRLt2uiMgXHFzgXjNUHxoOrFGHbTCVEXF9MdOhfxrg
ulSIcr1+E5DtlZ1huxcKTx59OKdUVzZTiA5pjjX1aZ7FD0xSMeUgNfB2CAwWrOxT6qM/K8xTwgqY
GkF3woOQt+tzqIApSX7OyjKrww8Qv4a02//peLRTS0zUfc8vko/KtmitrFDM9MQ75g9mKwkIadpW
LVuPQK1UBfnoV3flxwuDH1zmxA6iUpTTbcyK4TnEeIIYHZ13DlbVxGCwgsDTVYpxh7A6ZRBjfwmO
c7bXwqTD1YW8H9aK3XBznRuRf6PpOjiqGw0i+Yz3zqQnx0SFpNkk7WHL0ZnoxSMgE/Tcueskwv29
D8w6PjTo2I8NtsZVZ9PLYJ9JuFX1A+hDsz37N6piuW+V6+pBhpSswXMMXRumMmThsKRsZrNQ0nFt
zkLZqVC88uYacyC+6jHczCi7ULSUfN2pbAgF8u1+yX1NTFI7ar0Px1n3mprnfZeEjcTCjyxgH3+J
GVPpAHKsoURS7O5MVXhlFjuvHl5dTBK6m+xmkI3AzSOxDcHH8UANu86nC57/Di2QQE3XYDt9/L40
j1nBSoklRolsQqEaFbxZeQzANercZZ1LAWysmbXapDaQdx9XQ6oQPLvu5lBXButsceoYt/P3gZCh
gNWIbXg8V0HKcbgk4sczJHnYibEIfDN31HUHGbaPSr2WxOzCOkAA0XvaA36AtVFCuSnXEXjspkr+
TxTHrqtZeh8/M2/x83XHaK1htcKzztdbObFLQIICMqveUzH+W+TsLp/N0md+PSAk3rK6gwLoBrTS
YshTs4BozsK/PJ4Pkd9r4eAeyecqNjPDM5DoKfJyeSDLf1id9Qu/0tqyEN4s62gihBsmNEZULHoo
D1PvT6z8NcjOSExFCzkW45EHjMzwVcE0BakpG6AwiucOLwFXvCDiaaTNkCABFyGbdL/OnGiTTUhN
IZuXjkeWiB2i9R08SbFu8jlY5WQ4Bmr10ljlslHjs9N1dFJJIuzaHLNaS4O3tkGrntWcFi19Bq2r
tXgkf5mAbS9AAMCG+sMGMq5jl26JUSXIMMExJwNnYvo2kdNrul853or1XPX1R6bN3tG8ndy2/AeQ
Oz8n6sBrfk2XRDL/A0YnRcZUteSK7VQxVaXepVpCZTyQDpozxfPn9sfZgEq/OLmmpVRWdIMReubc
VDEy1jHcjAcGIKY6SJIg69/tN3IPMQ/9d3pR35m/z4IPHwA5qX/HuvhnjgLFvL9q07eQxiKtSpho
Z5M1Q16qcySlPpH7yLso7xyl0YP1S1ffTRxE86V8Pn+6DZmVXANuYz364GiGV/yUyfjcvOubumwu
SFc+EVDrOxH/1nE+Q4Y2Tuj/2W8eLuROlPiqBto3rzAGkmbxZwTHiqkPwqL6WhxLF35znuH8s2V2
fyKyrE5U/842nlmhVx0BDUbx3UxmJalAgZajWNoISta8KDfOfi0sZNhhzospFxpj0BIYV7z6jrna
DVnrIdS1ygCmCHk/JzzlVK4WY301d8C+a73fIKLuMac5YUd0iTTPxCvc7WubNhKgMJDsbqNSa5Sg
sUM5Np/ZwhKjFTrRbqhKD4uj1JRKyRUqIF2PBiI3HBqfQZILdiNKRVRGg/deSi1Cs0LrnaqoRM/o
MI+dEmZeB8ETRDlqWWUDG/zTtJ+hP0i5llxH+ZSZSxmh2lxMKRVGrQLWQPChFH27zlvjF0G9SjGS
DhNTQpFtvPJvku/jyFoIUZ0FBspCX5sB4aQT+AFT1tHvm09KlKI73F0z7QEX0gEOwToYYdaAbuBV
/IST9W7gQh8x1/zxCksVLONJ/5EuxjgwQDk19SP7nb0GbzVQZAHx2ez8U+LqcT+Mt6WH0wezeKSn
ppEm45Z91WTK4/STJJqfIHG5USyxLELmSpIB1AHa8XdOTy1vIWwkKtf9ixMaYEEcI83S+Wa//0pI
wNqrx/7KuRC5/iVlMgfwL3tJXXiX/UABdN149l1xAQSNa/X6hGS7UV0oR2lh35aSiWgqs49W1qdC
+q/EhcIT4ELZmyy9HMQVX8PtV7goRFlZK2JFrq56Lnr0IfOHDJGS9UEY9pjYMmGdq5YuvDaQ1SYF
HRaCFg7/oo2uFjF9zwLHuUgyXwkVPU0Nwg3or6p+ZGL8evU0vbBM4I7dq0SOMngg6rlNVBiW7vK7
yzIFU4psWcuokDyt3vc3JDqv6+ILnQ6zLBGxLT3R5Wu4fHTPMdpzzr3YDz/Zd1PXYsz+teJGDzyy
7OjVwQ40JZ0jKiv5KkvFwN19RHbxfOaJD26ghmPTwSiNtz9g7yLwjhuiETCcq1U2bhd4G1ExAqwZ
Oil93fUFqreHx9KhB2Wv84iWapLt3N75zzDIRY1/icJb8OGIeLatdiw+wzI4psy+xaIzWYZpDtdK
j36bhjY+1H7z8xs4wHLmhzN5aSaXxMpBlbwe39clj2I4bK4Ha6tKydj+I+xNgywvGF3oEpLBJvD0
7eGSklae1Ss3tv3ff2+6PLJ8XAYrbqQqCG0X6KoHbrH6DMBvHKUVE0DuTYxyjKUYMvJ0eLShQa45
SKJUaEHgN/1Vezngz2Tz8st5Qzi57A2eJUCcY7goiV7YEQM44gFJEKyyaoN7awGCo4TAwISgCaYf
+Iq/jKAfgOit0g4sPno/tV9g+15CkniW9jS0HqPe1ExfHcYNC+HTZfLRrslZItR1lnj5syFKcFbW
T9i5AN8+cGcHk4g2vquZjQNGt+1WwYOsJ8HAsfsv4jnh8YvGkIR2dTNopi2tL6zBxaNb5XV0e4WK
Aq+eRPjDDnnir0T926tazsD329149Wkt/7peLponXpF69+OR0By9IUpNRpM1Ab1yxjiFs5xDLSJg
p2HftXiMp6u5//gSeydm0Je1gq6+ZrR7GqNzV+1QX5z3KW0O1B184+t+1oKhh6n0X2F8JNoM2AIA
fdDEmkHryQJX2BuwvPv8Ra0YCYHQxCjHcLmEkCjRbmGyLCcWcFw7tP/V/iGwfpuz2Gr708HruAIB
rKTf/k06KPaMK5DNQxi8d0nnZq5fg2axCsmrTQZGX1UOXk4mEPnUujrCz7Y7tPuIRjqdghudJ2PR
oiHCpD0g0ncJmTMjKQBLY6W4siRx37fJdbJGVptMuLIY8pAShc0i1ONc7ECl1pXQ+RaG4BTAgCC5
sN1u17KLK0qTKhbLZE+FAGvA1RxFd1sYM7yxA16fCcyBQatt9L4Vzq2wx3Ey+NhGgFyB/ehC3Tvh
6cYnZwYmw0IUUubFHwY00cDuYide4dF0CR2Bhf2Y96dGgdEvk1pxJ5vNTqUDhV7KALgLmTgR9BYF
t8z7fKPLA71oSBQZwFCQPWr6E7fi5TlkgB53ubQLrUMy3IY+wy3PoI1GZMD7fPRtDRfvN4pZBHOU
w4OjTE3md3kbBz0XUnHzM1/m3OAR3XDXR+O/zXMl/CbLgXY20bGSZoIat3FLlVgYiGk+PGXMNQ/T
cZUSpKrINgYZwao3V6qDMy96jXGrN6Wtdc91yM0fPP3fb5a/dulJPdfzPtoSTA5fgh8rUHezLTLf
dNp6FuJcOZgj3JWn5cmrZKYz9dA06NuobYWxNaOIyE2chi/JCfXI8Ngw1+cJEuyTbUaT1j/kVphJ
MXQfPijZ/Ls9zod9ZHLTCz0K8A2F+ns/SxnC/6I4TcvqCy3Acaqkxy49LN/HHiJ2KwElAq+F2GVJ
lK32TeQrVO/z3LyC5HOp29VYLIvEOmE8WzScAGOMvAxo+zsPuULewxWaXAcwogfRDN8IC3PK0GbG
PZiA0Bga6mx58BnVj/fg4b1r3ZkA87RLCctkwBePRzCsgKoii9KiCpq2dy6Iu/+ixpfP9x+/6GHm
7lMxaRldQ46Mt6V0hbvvKaAM+OaMVWzrQ8J+Ar/FzaPKXo1Bo7hRKhnA4nijCZ5JYFv+tkgvK9DW
x9hEvrho+BML4Lazb9J5TGiCvvrlptjYcPJDOiqUBd31SNB6PgbE2Xz/ksUtK7gWRgsvCzvbedaE
auWI4y+qXja7r8h8b+NX6si92VK6YfzqXIkaWxqcf9/4oXj4BPj1MTwFMZVLrUhdJ+5iocIJyTjd
9SH6WTi7Rkc1MqrQqD20c3owhrBkX5SCRK/RjUmBe2/AhIkTw5nMEXLEploPfLuz6vp8e7of9EQG
0Ra0yMvqxMDcxp2lwlJTOU+wG+0Ae1dV8m4A0msk3p/L9xuCjL6bI1E+TmQ76DGP0Puo6wCApWyo
xP5CibvxfZkzAO/NnUzgOwklgzBm6rBIQuMsVvD3hrzOytMFz+EUczew1fdc08XyWfGyr97czVhx
q/bBJvPabDb2keB/qPuKKurGWvbakrW5C1iCwvwKED09j1CoHZXw4WQ9Ir5jPKbAfLjANLL7pnh4
scbNdBCpg1b9sDBTM01mSRH7bw2XBRN8HoYC+kMQE8RnPoerbGldLYIu7LmLPRaSxc1+L3aRZhs+
FqXQNcekJ/oQ00sRearbdg4WjoeRwozsmjeyDNgaMr+6d6RXvGhG8rTUyFswcYLxGwbNK86i8qMt
YYAZd1YOgp6MFHAjpa7Hl4WUptCPGUsXAZ4FZWL+u5/aYSFxHMuj/LXg1fC5lLJ7qAvXYTT8M5cN
vEmUjHM5+tE/WryBhGX5ny3J/7JfkArR9b4D0bGycl4hXHs+8ODaf4ZtlBozQKf2zXfuOr1iT/Q0
uiJtYR3Qxz4ZnvVqGd2LYotQMOkHjE27f65bwR5kevp9FfCg9Wa6UjLPnQPnPV6v3QZ59e1mweQJ
mUPb77Hh5y9o0mJ8QM8aU7yJ1XTqgYugfyBPzh8DUOQerMri7EjEvrb61qN930n3ee+CxR4NoVA3
i9RuWNFPTbPocZbujtuB+sxk+diedMYKVt46DnO6J6WBEbFwpGWH2HHLlRCcHLdsNJ+rwl4Jyyv7
rqZ7L0+gsDG3q0UAlLqZPpkXdSeusT/1LlF3tWZVQc1tivLYXDl8Hs4NZmifBigplNyIi3vT+ZAW
H04n6F19+IcQky9/BhXtqtlZcZ+3XVmUjgQ15cMdZn48EFloS615oe7xeKECg/diuBsYmtPn+xDb
7VEwBsuMe3iw8P641KjohSiLrCmuZQnRdoOZE5b3WNVj/hnk+wd6o64lXHsiFPcWoMeaA3TO3mtS
P9CXdyrbc5mpPZ6vEVp0BedEQde8US4Om4wQyPg6yQj907K46lh4CvPa5LSOI5iBj3lEmH0AxEfu
CxbODIOqnDC80tHiX+UtujAAy8iI+C+LnF6ebCrHk0S6Vhn3S4vlZX9fPnSPOHy+AdGnsnGJiaTJ
pOPBXiInqgfpf2nKMTH4SELva6TqfmDq3Oafyhih9+WCGN6mwb9oIqhSsYsDvILXeCkwy8wH4rGR
4Y3g1pZf5ec5lDuMRGCZmMNHPc/qOEdDTTMDrHLo0/SntEROOY04RqC82a8NCD5HPmm8ej0MnwjK
/Yfl/tMV4izb4Q45ngYnVrMzuY9A+ULfk1MFufIRAPygB5jCMy3JA5xUTGFQDJF5j7SIpbH/pGBl
Pkd6+/3H04VeF5ig4WE8jVxdJO4LgHsECln67XBTmp+el8UUK+lv7/3UWk7rHMGgk9tKeMiF+b/h
DAk2OZpw5/NINivm2WjPhLQVBZYBr/QPEQqlE8CB2L3Gass9cbVTjWSd2kEl2ts/+YI6kGNFvy4q
KpsWWhZjO5YafLrLs68QK6GscUv3gmZq1vlrF5UTl2KNv8XD5Zwee0RxPam8eEhwS8t5bveCnoww
NhMkdGETSXJXbSGhHnuxk2Gld7LmRdpiya9g+aGtbEFGDBEptbjBG4vcELA+Ji2QLWurMq9SCytu
YUy1CY7v4jW7MsvBnXEXUA2qlimh9H7RMTVzKEDdvIBt28sFvUzaF8WXPTrgU0p7opv4KrG44apa
7H2aKgt8T3FPHOGIz2lFrfObAnjfyRSbtOmgCAV8HHyienB6TCFQy+aMVcj1K4HS15t3/0MloT05
D/UO22255c+yY6Vu/I1JG/6DyLIkV+zt4D4T9fNx/5fdaXsg0xxbj0XsWG6uGldpKVqX/tbT7YhI
LxetwDHs6AjAMnWx03wxS+QlWS/5Jo4HjUSLR4KpstvjfasrbT8Blsz88J3JmbSqcqLUwxaxhRNz
7ILu7MfI+dGbGqM5qOheFAtp+0vJxEzXKZCBKVLlfjvrq5MWqGQvLrIfqgcGm8XTokzwyA8mGXsB
JbGv/hbaksVckhSWx2XvxdthnI+6L63sx62PNdUl/pf9D776lI8a7Nos+VZGXd0OHnkBjZ2UpT9v
eDbjFBfowe6IkoJUCf6vVVEKQshzeeIdlz0cLlA2yfFotUfzErS5javEGztMJgHvksx831zs2Ry+
FyCQahImYMgXpUAqZFTEslNC7QVbPy+yJWvEv36HImmXSiCCL1vUaqUeoJbOmf0XcLl/bMpK2IIQ
QdvfZru1hag9YgXmhSKcJMCac4/2P5WpWcnXIrzKp2MB2SXN59jEiXqORUBUXFypt3GX23bnu4fP
lejDNEAq7H9s5Cf5pUrcYrPEkN1fQ3yr3SMJlk8097QI4DLYQPLcWyZ5hL3ZHyGcopjawqzStQ3U
rYWlviycdzlNQQQ24A3qIeR6THC8LuAXlM1Q6ZsIj4tODryCbzeyAMAy/ybCgoXDzMEHNIznrUox
oD1KbRo+2+F9OAHRiGbQsRxGU8UEoDpwGYbpsd5kMKfeHkaqY3iBNEvkWVGwvkGs8MMR1FJhuIe9
qyTO7+V8TJg+G4p5bpgtxnMPrHsgkTm0uS9+W7Io/xrnqOMBoW2yxrkayGXjuTBo8iQiwI0kpLP1
XiFpPmrdXje+CJ/Uzkoal6jTRv87Ql7+poiiVu3Mpe54e5dLJag1q2nefKwuVtyKcf58zUZ5JRXp
H8WIYsm8tgiBmnrEeooN68zeQ+Ahsts5F08yCPgNKLcPMnCeURG1P6j2i3YvfRFg0BXxPRkW7/tO
2+jXdPzeQbofBrmz/ARUC8GqCeXjZ/qIo7q0nvGl/U8Uk41e5DwdZHRwSX5nay/4fpHuEdC4dqls
ljonyXWgX1ZV6LDCgiei8u7dshj2BUlWrfkA9TQYabyCEuf2UN9Ajz0HooZNdPuIev0AEjfsSczW
irWNkJwnb1hv8YEzlGEik7s5iAND5fU9Pj+92L8AlquA/NVMUJrOf0YWoveQI4fVFJ8uE29TpTeS
D50HDyD+u8wYsgbUbqjT3Z6P9z0FwvxWY/kvCbt9a/CkagHEdx9UJDpUkb+HXqmgkS6X3Y1c6/nb
xZQ31sCRx9OEzFiYh236h/a5VNZQdLFGCjs7Jfu+LCtfm+nE0VaWx/lRRlM9dmHeI6+EazHw8z3X
SReM/mFkv7fAwrjTfefaejIiYFPp0jvlp8TuIfqj+ifjxJdfQQROZgXzfBL6Re+Hl/Yb++pjB6Qr
tGR9OVLnASOpSZHJcw71FIMjKG2l7ipU+vAQOUf83hbtnrT4R7OKx9yM2MyRmyMtRo69pwgC8+YT
xpUQqnNy6dafkiy5NZrv4qVknHwamo6owJXD7GxQryz2ZUNmPUJ6LUUO95yBXqRSVCJIYoXCO/jc
zS8Ly6VXq2Z+X/zKhYVtleXH9yPjgBHfGTLw25g8cI04LZUYqhDdLgtRJCoFpVhxLdNxQ0dxmnWw
kWSUceW/UbcK5Vb1jfl74axm0n+gUHZBu/LlysifI1DkvfVVdiFqKxgxzv2CP5uxaOXPA/E4KiJd
6l/rN3GoZyw70JyYCye7GYglby05LydlhJ49ybN6UAN5R0Q2oyj2D8zR5fhV5GWazvsTxEqh0Zx5
aoWEGkSbMFsB3TpwTPgmoS3xYfUiKSnh3lB+iF2qzDJ7D1j2lwPlUsyUYIPkrcOyiFkfF1A7O1Af
X73aatsDP17s97PU9SUqdbao9FvZXlJJn+znkKP6B9ncM/tEJEAVg3y8Rk2nQqIb83yXdYOBIR9m
hnKqNBMyphNZJ7h2zyILcy0D/BnlJ47bP80zl8619YSLjP0t2i/QMX3xEBRyEqalkH29G4hVmQPf
S6uMZ8/wcZxMPqOV5I0GhJdyJkJylRfnjkOXu7d2cq4Hr8zzSS+n/GK+JXeprbo52PyS5LJ0IXeL
ES+ySNc202O+vu2fTfNDejpCski0Wlgvww/z8lEgV6KiJxegeUD5ZNEWdg8QSHwDdBxYmh/Mk8Mm
GBpcKpBvcqnieLgvA8p6vr8UnO+iq44/GeqrW+bBoT6lFiLLt/VIGZxeqgd30Fk3qXMkFGzygWCA
ds20rSIr2Zbh/yvjKn29U8PXLabjnJuNKrlhT5RLDbHRu4rqaJ0F9/CUVqiuZAt/B0Vqb3jXHr9+
o8p7ip9clU2Qfo/Dhc4Ndi18mG9bj9Bndbhh7abDbvWmmrx8wNy1QOSh8KvKDDfg/KJ/vUeUZmDD
M6brWWtUK0XVvsVZEzO8xCwQt8Fda/UT7uxl2caA9cWLcQney25DrjceosVoGDH8DTCyrtjuxJP4
0eMfIi+qRmWqSxHUoolgk60tiQMHls203DMnmhwlbcEvmgodhv4lFtDAQwFWiE8qHm46mRrmsGb8
Sl1GOC1089RmIBbchMxpJOsyPG6eJSpMftZGhd5In7ijfNbNduJ3hHy+Ilsg2xxQUwLtC+BKf7IA
Ey6F6uErPxBh6W/sYzjLyz8nGanQdak0mjGGvTP0AKIzb9yynf4OtcTrPB20VMzULlVzmcB6I01x
Y0Si/rKu6zQ8M9pTh+MnG4EEugRk5VTPKJqBf8WUCvfurdzvk9wYwd6bl2VpzOKL5/LArUWjmAHq
xseykB7/G2eEehpFuWCoHtn9d/Ood8JA367G2f3+P0XHM7xorn9uRnxbA7f1WkpFWVN3GK8UxOoB
55L4315cGfBn98TkpGGKlpmQGCRQK1FRpDfTy5bE4cYUxLrnCFLHj0v9FMAH+HMcVCOKt9e5MpbH
Pu34jYO7SI+p6+wnFEnWojWSg5QzOZr/3/yUTZgYFsd6VHT3kjbr9I6l2e4Mpe55wAj5+30NXUV6
qF2fzlKCs30Di0spYHQbkBb2RoRBo9HTm9CIu+wcGFpATUC1vedrINVGaImJsDdRnfWBtScRIiK3
cuTwIWZHdyM9Ejt3WbPebViGvSH16uot7oPJy4hbaIxLRrOxp9Uv7Jx/yT+CULBYOXAg8rs7n81b
mxFuzr91HN0MQDSe/q1f6HFuCl21h/up5A9Io1kZeOiJlIo9MW/UKUW2Lrhqgoja7ppNrPsZqgbi
rFf8lI/rB4Dcq3y+xfrnnwkL1VYYZG1ZHxLHN2jDMAt15zrCLAwLwtE3pePd8Pq9i7aNik8vmPn3
LBLEMLOBMJq6vtC5VK7SrJgd+1s6MMAX4PZvaa+0Tru8zLv3tiT2LnEPXt6AtevZg+Jkjhhd01oA
E7e579hSIFsVKVjJkzcB9MEKQYOCWI5A5bPMJ0c3jnUzk+lu0JQFXiUj6UpWEOxsH/3H9tMKaY7b
0YLRbM4yKStng9jDWF8I9BSL6RpXMVz7nltG34A28xM4Zob6UTQ8bnD2Eqpr0u78mZTMQNR/bxCq
7/gj3WWRPPTagene7T6dSCyUsgBkiqC++RXMbnJvFea0XPZ/Mis9CM6GTdRaF4DB/DUH5eJ+zNfZ
zJyqqoYwcjwQWqcEk2hTukyyMSH83fphkiz+aVpmv9b5h+3SzoJ17oMUiq3EXKYq0S1JwpOW8pyD
uijnhpG16ev2t+sYQMEXUCd2qZDdMhq9mdeehuWguZSPP/Ohpn8BqmuaeX8KTwGtrLz3ARKSgwdT
fv7JnaRy4ipNXe8SmWBbNI1+FmMIslJdk2XIiPoqM53SBIZn3FlahNXa0kSnrYMQT8fWU+ZNx+Jn
DBKDyKKfWoYzZfXSj1YWuYvJP9CoSDcfm2NAvis4VtDOqqJiB8rRcVEea7HscsCgrsxydsWB8GSQ
S6NAhzhZzC7mB4mVEVlxlSmA/yxpnsFFpqrh+FwJf9anm7HLEA4T+eYHc5nfqp+a0U5ChAQs37wZ
/LY0pb1vzOVUcFtsnOQm2/RoTHPkZ/C/U1vL/lVd9VwCQjMt21qulw1XoOVbHuo8A/XPIB7IfJ1j
SGMuxDObmvauozPchfCIQFiZMYt5awJ5CXcrXwaae5jGnjN6rKW4kw3vemT7+s7AyOP07QZYuzvT
CY+nCU5xJ0PxrMjU909Fjp2a5xfAuVVVPjD9pFCcGpe75K5JmvvsHk++V02fNUg2jd18GYcvqUXi
9kQ3WzgwxUYJxrp2WLl1rjlieBJGHD+uhvBC65Sl4e0jRCwTwdQh0CylhMeafbqpfj6w8js+HJGX
nvKWLDVSLkSjNWrGFH9d8jEIyGezSp6ta5HfHsPJNZjJUciQKOjHFuYCXhjw6AEQVz2fZVvpcIGN
H24WbhUyohr9gELiUkrzzrpAkJM8oBDVSXTZ6g6Lao/FI5IMHJek7AwYRkT1/oeXoarD2/bJArCP
tiCggry8m9oW+RT3gclNuvC5mpGmV1+f6HQAvYSanFGzA96fmtra0t2lZXyX96EBkU+QTH4SvEAT
NgJXExlcm4O2MUjFSO0+au4kE/kqmvjvON5hKsN/MKjBr9vNqrOdrUxBfP2ZxuQJi7EhB9brqvyE
l2i+A3hGbWWrlkcOQ7vLzxBPl3PXEv0uCECMxy3S6053wWH5VJ4pmmfhUDAsh4ZJC5NYwWwN8Xo9
a8CTE1R630kWiF7KVF2cVSNcPe6ULAQ6RYX9Wpaz/15or5PQ9qbcy8KGG5DEyhQE1tv0xSDsU6K/
vUkNK3Pd/sSqoYTOE1Lpq1+LHssNCC57UDLOVREKLe5sRRhJguw3Gyss8yeq8i1ISypB5md/60b6
aLsPK42wJzKDG7Nb8fJlszNXy84olOs0nNkajhpaC0fUhGBTANZLGpD6CkIeqYkZ48gcQJaQ+p4N
rXaKVH1Zj/Boak++B2OIJCsBUY6WNlXOIzv080w4EKHdQEAHUqExJY6xXCY4g9yGYMtU/wyeVj5K
a3vTvm5VJLXyKCg3cukY3rnxjRfLEQda6VqBDELDGwH7T/rW82OZFtWhU5gaQ1tnzllzLtJ2Gby6
djg+MramlZu/rVlRtLzLof/HPkSyLrPVWuHdXB+VAyKRniQ+jqepmbXYQ+b29hENopBeqPElVoV1
WpNwSflSehwc03R3Cl6/dNy5uhpAk5V2ijE/CC1dvP7Xjg+6bZqQcSAzWNLYOY4j48c9DK6/hFSc
1oCl2Nf7fqPlnc6Q7j6pGrvtvughBjvSJrd7/fEIEPvrcbIlSLZP54vTnjz2GMsHkdYNgbBgeE9y
wlHx6egYT8ER3sTQ6/2JqjbM0lseYfyBJUG0Ztz4hZPY2dxVVrcSyh+3wAVHdE5bAmbjSpd2YInO
Fw5MdV4GT+PV+5ICONPlgs1rlf583V2us6pzvdSnXHNv6B2SujtotgbxWFt1/uFkoVdsrI2qY3G2
F4aYu+44v/Nmdj5+/Xw9Ss37yKR/5Jbow8zAXt4qZ5q8G7e1X8frGdv58+MfvjqFA+gVv+HGRasP
6ODq6nKSHMgb2ij8HALuAiGSM7JO7HqqTOcQGLVDREpYDRb3DeHvQB2r25WSKE8v9tz9xuG2a330
Zto2Ti+6xmnfXkLT38S/RVTsJB9tua4VGLQkEbqTJAzpBSQSV7JPc48aY051s3Kmp1v2LOH5AJmW
ubn4BfoAWMlyZYQw621BFyOZX+0CdSAz3VSJVGwJF1TvZ0U90GWF28g7zjZa0K7HNVPVuXGoSihW
M9W66aeHI3mJYmqVvY2HVTG2JDbs6ycdJIVIKwK3UqFehUsIEbb1c3GdwtnOodXBIwy82rp14jXV
/3X65Ikf6lSU5u8mvOMfbR4WdzFz4vbzI7M03t/YehDLCyTvvO28ShbyB7X7oypM94c0i0DChuIK
oaAk1+NLQ1bEgas2HHGMPnWVu0jMWy0/KwvJJ2ra+m17i/k8GL+Dc3RIiR1fDHpG+tZVIAd9Wvr4
wjMzfsw8dvHRmvvfIdkif9xHBQWmQZarvZ1r7Pk1bgUbDvyKLXuROekqDtVTzxwbCjmXFD7ASWvR
il+EURX2Jl1ZPwa9IO3uWEweWR3F2GwEVbI5K9Q8Vgb51JeAH3LUxovH9JGFzC46UfMyyt3LuUL8
vtoYEycXotErVk39tzUml1rnKFlKqNdt+PLsJ8HiOmRFLhx51mtifW7xq3UddlSvv5S95lmNAnxN
8LfjAzl9UyUDzroGFoakRB+l2AtoMz/Q7rGsfiwoffQXC3qb0WhBs30ruKbEWLzwNMA7r6vk+vhS
hOKDonhKx9iO/uNheWB3LMRkgfdB7pi+kJzdMN6ganHMWROVVtHS2ga5jtllfRTQeJnrqIWKWcnr
IiXnuXzIf0LzVHVpUBF0HkZu5bnsWxykXcNb3AEvq/k3WhUaWD7Y2TNVdEIvrLTTlUh0SXRIR7vS
GChQn5IpxHqLJSX/asvs6+RF3AWWlnsIusrpDC6HPuAuzBDlSpfPo3aH8RkhTYyCL/y9v4PUxATq
NL0oQ6mOrfeAm3oa5XFezkLmIRSG6VSthanLfQ/b/psBEYi0Pr/v+K4Vu/2S0J6wGl3CwvddAtCZ
MPrdynym2BlYfJXVlxcmmb8Jewph9iRCVbd6yTRr8NYpPAqXqSlKamP81p46D9DOgxpvflW2UbWp
0VHhbighU5Dndeh9gugTJLNL/VR6vfGwd+bExRU/5IQyYSRmlK7h9keUPTbosQYbLNV2nSSbaZmy
FrUNjJEdQR+LNbFFB7QxG39vlObH1fUhPcDggFcH/CplS6PIVhnv9R4BnOM5pjZq/JdClckWvDGO
H5SXuqCnrkts3f56IEBayZBT/iSZmYwqmCEmDtvP75p5AIRz4X1CsorjQf8viM0k9pF0ee+Hip+O
leOLUHW7BHqA6ov/onlp3aBjmG3ELeQsS+UT/pvHa61OXGXIylcwDoLM6oi03WcQ56WeYyjGDu9F
UNM7VYusQfALjvVspFGmmp2sEt39n2kKep/L+qgBzmZ7AM6rKT1JhE8bD08kJnnfjk0Fdht36uGw
xo9GTaxC+UrkqA+IY8CQhUfbdT6c2oGIavYxvjw6SZEB+aalFtxds9cqiULVoBbJf2Qxh86MwHB6
W/1E7w1o65bLmqehVJrGoR+eMjCssk+2dyZKvoc+aa6SWoh1J/di+pVzwJMaTY5bfDY+2NoLm5ON
QkRpTjNUiU2TKz+VGowy78+skDuAVv1vU+BzO2Fk1nwQzCj3tx9ZI/TEEQtOTIcGN+v0GVQrKQEH
bAU9sZVTS59ESlfKazC690jsrNLvSK3kiuAF6Qk1MGW5YSE1AcJxt8tYPKP/BR/fO3Sxm76UiUcd
Cl7KH3C1ebepokjjelFK6heijftsq4H9KXeLhKvutkjOjgpsoHztWYd7dldUT9tV6QJiJhsw/eWY
Sr9rkODLIs6JL+dl8Dd3+nq6T3Etqs2okvHJTM0PPCc+hstl4Kx6yNfN1rYrvIDDDbQtBX5BQ8mc
9p3NDCM3R4/RRmhlB4SUDm1sDg60xD2jfVNnPMA4Cwj9cRs22blZC5NoYDjNifdRG3iVAsc4wWKB
g96RPc1xJQm2yQJ40TXgoiIM6kh3/JZb8hodME0SGKGyhZphgfhuRRDgP9onoa6uzJZPCLAP7bol
5Q/DrJ8P9d1OpXzziYLdDtUwEOEAoLkojqdA6qwo4KlYbhnCVqMmKPTXmSRZP3eqdlx7DA4Tfauo
vFxDOBoBbqJUGwlzu/bToGlkYLfM+/KmHZJumzc64j9FloACWwG2GyMDbJm3nAiFy8o81u65G9VT
NPL0UhGYHrOUnJOR0Dn4NhoPJRMAKX8ZCIE5zU8hEsrEyuQf4qopNhI3EyaHZbFjE33BbaeIOpAu
WqFfP9gBvywJZL5+1C4KMqA0puIWc8QKnIZ93EznU7g55ja+Hp4Lgu+wmRMlgvDwXtAUWwhkRJzY
1TodDdBoUXM2XReNo+1oiMHfFTxoLtQ4jqRJpECCFKq7He1Nj0PipxtQU2BJDBpgK1p3bXckchgx
63Fmp2n0kCYYDnLtOIl1qrTHBE15v+1jV2vtHX9tYqpIBXVb1i+QnxqsXg/B/pyyL6Lr4ixxZNeq
LZMTJDLiqo3b1NASJMu4MXkP1sqbaxsYwsvji0WbwtOe4TT58iGEuDpUSHTGSpRtpliFKjgiIf1d
YVsdUv2FvEI6WVUaJ4BzTy0TcstO0o97trBVr3VUNT4FHsJzNFYV4nDxGPQpdFdD8DovlI4C0MXh
p4D/7w8GwvlaeyZFfcR7Qhr/pbl4orr8odM163NiJ4tBhKSNo59eX3NKEZlTCExDeAJ7FYhoxZpT
22JFph5mdP9falPb642RPU5lq30iZhecoCYrULx4iz8u4dsCFfqKGnrGEQ/o4fIqaMlDhXV2kwAj
fjdW3h/wi1kxo0bAzxHSjhg49RQh6GtEkm9yx5iTLQgmsxWC0CVQYjePZ+wZv/WvAuq1R44gmXuh
FF6uV59ZgmTXxlWVGZS4CPM5ZRNGddrlASk5yTjMJ/iPsrg8XYeUNlf8d0IsDwR397WEiAuwSyxb
ptb15BwTkiLH1LN1AElKVoFe0CM0jY1erW80L0lM6bWLpaFouNvOvjIbnCmupYv1jiblp5SDa7py
kIKwwfvvU4iLEdIeYATohG27Lm9LFYhfuDbXfEhgvwfWponVCneqH1ZY/qbZA9YwYrDNLU5Gr1sq
QxbGOmMQCuj3+MAJ9hwB5oZaoEl2cEI/Ol15NTM/fMa+sQ6xUoASxuEWSulhMckkuaBceWMIqcgX
bA4mGLPMQQD7bzdrXQKYvUrWPef+vBR34TEfYCtSTgiiTmxYeLBImaJZVIBGby4+y1fzq+TqE7EY
aikJXuOl59byCCnPlvzoDokWRVRBI1KWtg3MTa2ZLKYyQh1Qsy7PgQciuytwR3Qy84KTn89BHC9b
CfSHiZpYSPQ0Ni5k9eFp3cPRJrWQSvukOzgsl2aZTLNxSPRvLXzczHaAlwaLJGIyQ8fFl4L+zg0x
Bef2r1XUGt4pQJ/HmIPHCHz8Y+oxgCFCNFn2tSw95nZPrr727E7xYhxUqRlA5LPdezzEeBxoH9PL
qJuoaXwuSfYkd28FRrhERMLvT6aUVNCtGw/1VB2eyOYNzs9YtQucDAu6jAS2BOHcF78NWvOGuD9b
mhSEnccoXLhC1hVSFIZGvzm6T/mqub6f3VeEA4ugN0drVgk49Caz3pg/u2ElXpORXhvHzpTOJua9
SNWTPwc4lokHe06JSngrOxbfO39xahJVv5cFnm4LVgWI8HL8OqCQY76JVgA8H6GgAn1kftGgCqQc
xDiLiibmBMHcQ0E0HytGodn1NdoI0AQnzhXfdK2ZrhV2leCt/0lTYuta1fIT/gD9kGzWg67nBvJW
g5riw2XuFPJJGiueRGu2vu57T+aQiIYonfuce6Pucb1HjK/eD9nBdt/xv9U/Q/YMdLqnCQwQ3rkd
1d7sl/9Kw8Mv/fHN1n0mEBjBiTppXPMhA66vaRORGIVLo7XT4c2XcCQJCsENFOtgGFZFrctYpuL9
Pd0KzdTHm8MKlqPifoaD5aiGvzxyWAAJ7E/3nQItPexmGYG4DqDTrJcQDVeRbSk2NVnrhSQI/RPN
sb4iMdbAqLLFtxeX/y+8MumfZjh3CXLPVPVNqP6fHuE+91hRpu84mWApmy56JqPMK1/pAwxz9B5r
x6HyLO9ZEM9ma1SHXPuj0ZiP3dYJ2OTumbIEr/NjbuB004y3SHIpS3ecg3YqBI2FSHEmZ9mMiRbl
iHNO2mg0r7OCROTm2SQp9O9yke7B0kXYK+agL/IL+n2ocBC3hIdoPsYfIbUzl0Rm7rU17xp7R7pV
oUvHfbUe2/0aY5gEZSnbIbnCBy24teiwjdCui1lWSAH7kIaB8bDgvE5kGXauQ1iemAjqHgzLwep4
CH8mMjl8BSESSJ/F3OlD5Lkng7yC5dNzf1IJIeNZaHchgnM9pJWYGkzKuNWAJ9Pr2McHw3Ueo/wu
M77Oa0tXFLXubEtMhppx0lcR2/ZDc1pbaX04y1FOJtQ4eqGt+0j4UI2mW83iWaQktirh+9okpP2t
x2ETofymjJeUtl+22ROI+68AuiFPLlNpLuBWjViFPo+e3x6L8m929a26ccyDGImQL8LFARTD9lcC
VVNvmnA3H3rlYVq38hXX3wUK7tjdub0dsfO5YupzUjJ4G0OBqSlm/wKL7ZcpyECiIDW/mrcuG6F6
NQ1ZUCbURbOX9hq+TVZDh13lK8adAIhfCiBRNod3h2Tq0vZdcQcIZVQHFtps70fGDdrZWEOYYu6q
zgBrlSB1Zkts5lEvcTghltxqAeccvfQusjDiwupMtps4s5geBTauaXCv83aFfRmoaA5o7jra71Cg
AfKEWhV14SWWyE+aP8NH/wxDSub3woywnyxM8XZZedC6/E8/fzXZBLo7hqyZk98asjPSI1o+37vv
HLGf1HqIgvKCw5PB2N+kTR9kiFj4oylUD5Dhl8U3zwiIr8ctfOWr6w7GjXS18qtUpFFpClNi+OIZ
r6iFnGCGg+lvB9SzFIn8qp1ZnQJwYpAKTkHzwK77SKxRKbELbZMnaILFT6javvlrP5I/QVZJs5zN
gPtJNbYoe2H8xgmhY/TrkNg5TmtHrL3hrhsvf6cmuEMzZaOvy5dyxIfaTxBgOKpmpFcHuWnbBZFn
47h44QY0Ywd4y9F+gJD4ARz17Z+IPUyuz8ZlGXYEJXpWGrftQXoGgtVgLllA9HQPb+/5wysui1D+
WoYqeNo5eOztlMFwhdbOvzmwSsgbMPGOpBO4kvcf4KAWxhsk7repLOCmM7Gm2anJzvic8aoyepaW
XDFzfPqpNP67hdX/hVWoTs4EAVQRwnR9kPhPHMSsjGxkZSyiFP5QyF13045VduabjtzzgFWnVC9S
rGVHg1mq34D4sWJBfsI2U4mfv3YMlwRlYcEySjT3lugH00nDZRw6mOonI/jKr/CPlA9TMrit8fZA
RqS8apx3iRTWvcJR7pslY3aScBW63nAiyy7n+L3c0ns6HjSj2btHqA5utEDUgwE7q8Pf3CazRJmL
JnQx/KGyWciYt34DYOuB+COmyAZ8Y8RNgBPB4XD4q1AoS8CgLIb8xDvoY8c52HjpBs5UXzZxge5U
7m79zSzlFBUCQFWL+O9YZkREoBSDRvc3i5tsqwT+5SRghL+slH/AooK3Q0tedusf021eYMVoUSjX
SEl2RoUeh7gcqG1iNBE4boWJqEO/8dO7cwdZdQYmnKOrLAaIeud/nd60rQvzDfB3/naHQsXQ4/RE
MTRTL8VAp+R9ftX8TbkqzZUvEXeij5MBhnNlrwaW8lTmQX8sVxaG1tWygmvlq1ij/qGymtspFTYj
+B/Wj6GV44r10EpUN3nyAqigd00Zjo9oxnM9d9jceFEav+OwvrcnX0mknuahj1qfghOedZCm0wqp
kLGsoJDTrwcxbaZfJx986FAWyIdIIzQZhNenz6/fqRFRhmO9N1nN8sV2R3TkjLDd0s4F1qgLl0jZ
dKkEQs3JtYES/uqGrN26WhHOu4HhaR76bpAHUG1V1xFm6kLDv7KefqjuSQMbLT4FVMUGBFZnM+8B
E4ttM1aRu8YYCBcyWKN7QlNKjO9m7+EGJ8vv6hrfrxK21cRq3sJuSvgf2WL8tU+d1fQH43FYpsCS
n4ZFtjc1glY5lSBA3XqpbJq+TZ7UKLJ6tAuGucfA/hosr5Hc6iEraQ7DN2VCQse31JsTCDxWirjX
YTTO/pxrW9h0+MArf1P757ILeTMp8tNyz7SfdWzWdQGa/j04OTizJcUJ4nOKVnCBaGMd6uzQz4yn
ffdHowvbvioKCcWjKiz0fQbFjfuY1J2Dk1MbCtUDAUGfmAXTSMImR2/VSYS5XTdwcURk8p2XKp+/
EPHGgATiI2wLx6mWCqqjYUE3Ybs/qExbQQwLnU+pu9QrfkF7bsI3ohsEOdwcP9w8NwbTzR8VG6k5
bUUDKoC2pKj2ENUEQLA8oQRa48AUDlCLNqkLmWAwKmw3XlwVLXb3TIPtc2KTFpGXV9ZNs8kKU6Ts
aslSaNtjlMz8zte3RbIUTdHkzfy8NMoT/oe5bnJuMnsF0RORXpsNTuA/3zyO7HW9By1MDDRAOQTx
VEviDmQowNzebQa6oaaNz1zlhuCUw+LN7yEAERLvavWVOlQxf5/LFeKU6huuHdHdcuDwM1OTOxzl
T8jeY2pJmjpCWTBPJgnalITZQSyK6fdvA3Yz/BIUjzTqmHpJMCWyPVjiRkiOR0Wh4jOHsOyadSZ9
NpIaIYx9sCti1/5AXi0HlsjWw1Ksov4bedwV6SxPSZtYLvHcML+pBvRak/XxKANRqCS8uG/+qV9g
FZWGa3T6xQvY6yjQz0JIUHUZFqYBGKlnMdJBGkxSxXLkUSna9RERcyXNr9CgpHNOqsZYywBbV4X/
L9zH5NgH9Yp2owB+pJn1Zmfjf179bcUYOVmNjSuvft3CAmfbxpVqnMNQy89WkaznI5dvLSkdBZnr
FSRZ84WzrGeTOl4Y+/1Ncg+HPJJ7ycOSDGXBQGdljYK45kp7SUK/1xI8ZkFuPjn+YwkglVnDM842
x58+GVO1hXVgPBbO9oN9lO+LXOytoyWCHWSDMbn0xDdMJ5hQPOyE6EXmtzB5kTBYJBupC7vkn3Ic
mB2zUD8QwdHUsxESx/f5feXu+CtxctOq6daGgAP/+B+PnBC+SngoMr6g2VYQFio0+ZYOa4fqWAhw
iVv/UnEW6IHsgj+UbFPn092a4mleMnxNguRNjhmqo97EB7G8KTsJRFkrWOvlegxtK/WQLcCkxASw
huPxpjJqJM898eEpfzc4wrXTWVTlI/XB/Ni5TqzQXFWBqPQyO4gG5PbhvZ/+vfHBrNsWPsEweNgh
eGDoiWpJX46rXMIWlNougKzthmiZv+TWrQew9rkgkGjdxKZfz9zFqMqbDBTM2KL7xAIQTY956FvM
gfk+8EF0ndQw/5KiZexGUmW1f/AXqa0qcn1NCoviuE7nQrmIUHl8HkC4GF9+jsJ38c6TEmp2bZ5b
0harp/38tQmZ6/5BxoCsK89MaWkNG8KrzuSs94P/cNAiZ7e2/CJybqekhejptcsFYRk3FTF/k2tH
PcjST3EQyeCsksv7OUQ3ZLb7v8JFNC0h8rzMa9XJNOJzgxuzzTotJls4ynne9OXvQw4oCOA1lxAX
Tp1dV3OM0jHyNJPzeOKRGiv66QVZnGzbWyyF8TwYdeLhS1UxeW6IFA7737Rz4GF8RNBuv6HxyvQ8
0oVu+83K1xY7lwdtNDsrr7VBPvEZ0ICuFKBzzvy/nTwndmOyLA6wJzrW/DU7szCDjB/39Ey+i+fZ
shwTjudbCSynE0W7b1ssJYNxU2vgIWwjktv7yxiXjXHo8HG9/aN/O4gwkkschp2VYtFoLoQR8Gt2
CtD6d5KiPMMo+nzlFoUlYD9P29+NIOTZkDalLPs4u3kSstH+zehemeW8SPwWPuN88aSJS+3C0KqP
JYLaXe/G7i3vhTQ1iRfLvK2E2jJ9dtNF/g7EghulAQ4pz/U5VI8bgf27zglQuLvvRhn3ad1xBB4Z
TDz2p+WDiB7azS0vv7fUN+YOo5DnrYaupY1euD9nj+QQLEiXe1cO3uFiNPhNObOPTpZ38BOI3KQ9
6i1tyWMje4HtVZ4xIGq6r9M+FC+sQVRhNMFCnju9dG4kGLmrCzAElJzSxWQfsV3ZQJ7baRrSOc6l
hux3SGrjOFEXtfk4FCc28iDhXrnDGC8AJlxeeYUKZlZWzHPP7XeYXTt5PtUGQtKA6sieeAAAJxJ5
8GoK/fj+T4jy80yNDeyV7/u/tkO6ZP4EIZOQZHDHIswH63CqbQjGVdqnvB9+uqFtRyMAyeO5pqvt
ZF4OtSEwnnXApqa5Hxq98TOWle5qJpYVSpUSDJ5i34ZPTpGDYYUC5Lhdv9IxupkJPgE9e0dXOoUm
P+ZpHlCdu1HgnTeXhDKYUAQr0Lq9v7QbkoReTNb4eeL8eFf6ZhwRPO6KFoW3SuYeOnNMX9Q/Rvxj
FCF4sUJVxQ2rmzNA9hxrKVnY4PpszUdCniHwu09bOf/ZBeoZcSrjWM39cz9SsvoXaZKzRcVj32bX
EbhsAkvuPN+T3VZcSs21vDVLYC876TQLmtHKudPXGFf8O6ZPAeenwUC6aKTLmUdiB9kQLL7eTe5z
BIz1Uo5FgVrfAZ5ULsH466G4B/qd7ph61krBxNh2zBJYLUPOMQ3IargcbERkV+eCt7gZeeu6x0Gx
4HMeJ7mnVJkafBFHD7KV6AS59sGEJNTsM41Z3Ixq31IPegPTBD0yJB/nBpc6XMv3nxT1dsoxF011
DnKTPmZzqq1kwMEItT5eSbQk9qbevrbhvP9/VUTf08yBgj+IUVQP8LFmWir2S5ngxAumX2iLdNNj
fjoZ6IkFj8r64PP80y2dICNovIBCczNCzifK3L946F4A5gXfODG7V9ovszbjJA21YD0aX5+38g8U
Vll/1ZuKkCbORLdVrlPlP0wAWvNkZGv4nvyD6Nyb7y3yfoWC2FaUyXKn+lFNBbfHixAqfjvOG56f
TklUI61sXV9fEHNrPXXl60n40SEqoObxPWxbz3+ViGVs4ZVA2KSjk+dnF21KH8JX2+a+N/HBSzUG
n8WH05A8j0Tt6719e8JndWUuqCf0+M/EsjCUanmRfd+rDhugjNAZsZsPS6ohCngM/+TUMISmbkuW
lTkVVGQQLiuKcjWnlv8lK+u/9A/OJfc/qp+BKm7dbpZKDok9+ALTLkxSthX7GK+K8GvUK9sL1QDV
12LJPvobnH/kaXfSMgq6fd/8G5awS27dywq2FV0V9um1BazqTy2Uy84Vhzs/Xs6QOolCc8bUk1x4
YFbMbrAq7CDHsmFtc9jY0T44Sy32/FXyn3qRTH+d1GgsYkj5dsvp4tkZX1fGfdYY8SL/SsBDMZvp
h5tVrBqUs5SbMkaIIpRRqtLkU1xms31oO622QBHdUlKty3HV49q9O0XSJHHY1hpty4JB/U7qj69R
S/Nq+TTAJyZMSDNGybYUFiiL23iFDXmYZ7WcGYYhZoc+mHt8tXj5WJdAnRwY4Pj6RW8o3UDttdiK
j6eO82OKkfGg718JqwvixEmAhcoHmygFPD1g01F+0KiPRVj6+fTIibVeR+GT7/txJQ+5vswJDpWr
30qU72MQWCppNZ2lnc+sGuQY+JPwRwydXA4XZOtVEgowQAzmQkckdrdPKUNNAmL9iOev7AXzUYyo
hhySxlCiJHbq+p/NVnz+cn3qQSZPnPlPWBy1UxHap6UhvGc6AhXl6Ml8lwVD5sHbsRfgOrwidx9V
PT+q10yEFRjM1ea8ALHMUsiPvcwfI8hw8Q54pL7AGCxxwoEaMe9VZt+T9mEXdRbECCl8nSnmDHvx
JZYMs1De3Z9Antx2tOp1YPu2pPaOyQaQsnwrSetmybfI6/3GzSDxhZN+2iJC4SBgGP9fw1sVzdbs
g846NU9A7+k8dOHNqX8jgP3+yRKOjsJc/kXRNI+l2Z2CDFJ6Kg07cyjdMmHIdwaqE1THOBpqm55V
g+Cen3e0PnHGH1ZT/rAMH6dyv3NhmdGMTgdleR4RxpGY5ktWO1B9WA/OZPP+8HeUQE7NaLudmlI5
6l5r7TD17BYyXPNt6i+BZlWX9Wdp0m2pdcaf2dw4N7pAS7dw2iynctitWCqRUVQGfKolB65u0pLH
d5bGQHZl6zpu6dM88aVjxabNuNvqW3Xb2APbCCRhNcKNrS/ly9F4Qj6N88NTJV4QLMu1gorX7/DU
R9VSoJ+xMRt/0I1TVC/jhtLx93jNFKfJndrA5y6Y9XoABfMspmHEIsLOQHK6arRYpZ7zg+DD7OOw
JB+ITmPVoW2GV1pAUy1ILckSNFqU5+Tc9teymz+7K5qEcBC8qPRLuFg2aXGONafcI9ZkmqqyOh5m
Bw8imXGfWJ7QPvd6ED8jQ10mnaOl9oPkjjSti3ReUSELscXZAvNCidt5VwYoUXKK+7qQBelAVKUj
eptaJDsVURRW8GKLK1A3o7L7vLu6OOlwuNSCFj21K/YrH+dMH6yCuKx27NoRFrwxonUmgycSjQ+k
tCLA3OBPZenB5HJhiScTcioJHu4DX7+OwZAZPS8K6IBQkB/5uvcEDYjRDxmyZBsEl/XNCzehRYKt
wfgPP6Y0YSeU866RdJuWbsUvXqBV92suNyQ8W5d8O3rxcnGPdgDSF5mOIfDzPnKtL2oqGuMOUgGJ
5yqr8ZyFz7081MxHxowfgXkIcqCt0JJvUbCdyr0COMepQTT7BDIBWZdeGlMM31pHOg7RBb7cDfVp
VOkLdu86/Br062rk7ZyalcmJ0kYBEyAFmoeP6xE9yR2+r3cItthp4oSoOzwri/eEzmFRrrc7nV7p
7JJ7JWNDLNiUwJzyjw638eVnal9jve2L3MOD59Xj1OFzqXKL106CuAsUoPyvdvMShIzLvUl+YSQW
FrLNwNVgWHV7eEO0ci1zGRcu1Qil0UhictpBsP9Zh+8/Ui1+avuRVEiS+YGfE35JoRwlKCEWo2FH
zfELnnVOTF96n3mqxC3x4BUmOCBTKwywZ9e+Fu6B868pFzJMdTEVAzoGtc5CFhEeds6dlefZQwas
E8E2n9zOB0TH0FgOujNlFUeKAHMs0t6mSgmOiYQQsK/ID8omIQ1OjAcsPLKE2ca2JRiMONJCRpYg
VREupbER7uW1tT2DWSEH8+RN7BWedGgOByBmOKQFHGHgao47jwEDviA0/KvDecI+/A8qH9mCG/Wx
jj0RCBNCnKyg3T4MPMztdQ3i5o7JNhthgkn5b/RDk4hKebudgxWW74d7zjYMOc13LDJ4oO2vyw4h
PvWn6TWvIT0g+3wQTlxOcnm0qMc8cnaKSkI5pWfgWs7jSC52uZR+2Z5MDiIH7M70ibsOkCmu1mTW
eurC0lDrJqsRGuZBevcCwdH1ZYk/FSbkHpIWeTLxCUeQRx9Vw27dPvUKMN9jFGv3uQZSiBmhU5Pf
D4LGqNMx3rq6Z9sUDVsBHlajxIfgSvjkO9h5vaTx1C7bKzZG7di7WXndQafObgGTb+Uuzrbba92i
GKFz+BgTveKSlApDTSRFj3EGJDtXVN3iXZ28p46ZHT2VJicKu2DmsbQw2MDRdyNZzS5Ovd5lGej9
+vN0mNZdVGn4/LjUIa3SQaRVRHpj1VqNB4TZxJMihJveYqGX/ge1RpgjYbNDvYKIerzNZeSQkrk4
BV7KmwsKPqEJfL5KdSXF5tpLQojtPWgUs3TfPZDxPITHv5dx7StiFPsOAljXJwrONoxMcuOiZd79
cNLKnfJI8EdQ6o1imfE9N0BriHerym2rUVXAVI3+Tbp4Cg9a6cN2c1jTIVfVqtHbQWtXo0seQtKU
8UFQebyyIem0tmEVxYZt5Las8H78y/RSVwdS+UUUNpyAMrViJfYHjeGPrxmqINdSBZGrbnI8vwp0
s/IAZcrlBt5yziyKv++ks993Oa2iRZhXwCw34f0SM+FBxoKnzGuL9irpqxPT0VZ3oeLe2oHjlSRY
J0cpY6YkA33UVi9vRBpEFqmKr46aw2ZBDQXBiHmdZpH3J0cM2xBV6juCns0gUpzuCy3352evvAL2
vYo8L3oH4QRoZnvd3Z2PrE66Dpp5+494nAOIrStIppHSmi+YO5zrlDlDmS/PwcjSD3FwWwWYRYXX
Q995ciClMADGuVRN0Sf++XL1C2WjELk0OXmdrOG6BiwSo2BlU5rr0gonVnwW2vt1Y9o1kL5MRlrd
zAV/YOk//B8OQcScXXZ0wfVOSMkT8UzMOsa2HZ1SbkIYXFW7r4OPd1PuCYC69sZW8vxyDKCNs1a8
WB0kswyo2nDrHx/uUoc/daqwpIjMw8h18CFyT1tqf2iQF6QvoQ/9LDqZOEkQkXjUrEvq5PBIJsAW
i6DoO169s36XHJ44UGh4zouMtNbnd9pI6tM208FgCCZApzX/Ar03lhPHQFdnuWqd6m1C9WTQnL5A
Wd5Z4Lpmx4G+XDiZ8m04UYiJpoAQ/xkavKcgwKI5WzfbrTkCwXbTRuAg+x3pOVXhdqhKVZalwn5s
JA5EZh8YLoRZfozwMFAl1bt/dFSTyIiEjQ3e3lisG+7HS+/3Bjpt3VeP6GxZ96siNQxMdNM680w1
X6jSGuY+0Rv92Z8ZfHK77NFMY+ZSyQsya6gCuQVPuGeoAn+5gixg1GVMerSNMJkw6mfEL32FAXDj
aBmLKCabxcl8NhPNclguFQZV2Gv7ttkC7Nye29mX7ce4a38pGzaPi7upsspJa2zYQLkNgtZGf5bo
jltkdC00bmvAguFN7jqpeuWWZMfCZeGxFRl6yC8YaotAbYNIapoYgXTXichmNB4ArT+HI5PMUxoF
jVQApZ3YUMC8aR92sSnBmoYSjLHXiNP9WfGK7BUUL7MDSHbm72NaRs0AuJx16tXtfsc5oqHDo9aS
/O1o9Iw0kZTN6jMf2yGeS8+Byyj1Zk3RkE9sq00LQVl2Ji9bGP8YRNvKB/4cRr/6F2RYKLKBJoPV
Oi3fkmNbX6sex4ubJ0zPWdZCJwZNB02xqFWW1Fib81YpNVvit6/msC9puaEqJwLnv2iT05SLHqDY
1ah5sk/5b/dJWE8zU1N+sdrwjj7K5xAtYLvff5AdyGKq+hpLonRi3sQXeyoWcMNoPS6LW/fi9swD
w58acShD3yCH9jlErnkl8wP+34QRfJcCHlNCmPr+6b/TzYn33SOlXu/wJ3FTID3RlFmbZ4ATnuV4
87THGGCcKomzrXXade7pKU6QqfqBP/1g0rkOR5VmM6Eobbahe0KSqAHg0j9Joc0hVnavXJeN8Ggq
awDi4FgW57h7tvvQ4+Q0h+Fzx4ke+FiKZm2cZ23STjDrm3utMLurhPPXW0Bl+jPJElFPKuTzUUqR
d4JW7xTMDXhWpk8RNQRs8K0wSFbXYwzfkOIfpFa/BvySPz7+qcEGgCwIzvus6R7GxLbnK+3/36Iz
JZn7NvnBUDCqheP2MD686i85cfB0cng5BxYwsRRy9mCwkuATPYtPoP0mHW0WPnmfpU4FfyCVTi+c
05uelElp5s4vwSzzNlKe27sKmg3sP0hu0NkswUH4O2ZXLJwVA+POJXFgzgQ+zboJr/P0Rncdav3h
kTK32snJ7jvHxMWQtanNB/cP6oGRFWxLsHsEVvrRdDdisq9JemqucZpB80wdxmHAJXOSgkI+TU8l
ugydFWHh5G0Ib/CzNSTCj+lAMyMBzyOmb8h+ilNAdu9yqxY0EDANdtLJIHrsalP7SPA5aPMWRv3e
bgMBsOxhXG9Kkws18tAF81VTZnVljU++7htwDXrBZfAVf+97E6lL0bSn+Rg35OOXjK51ILCA3Vpr
rF9faniB/omf85Ya3bfLc79wLAB/clpyu5piJtyMZco6F/BN2mlWtOREeU3JATkpxG9tfvzNH29s
O2GhUE7gGkw9EEY7g+u0hgiccwIXsSTsaIl8gSidu5CniYfpW4qo7UqgMsGTzH3M124eYgqqZLwV
YiBmpOr4YD8vubHq2EByEVFrNfddmcNDGF7VklnRuYUtykAj5CSr8JeT8Z0DVoP/RrMTJuaJ5pi0
17QEkslXCk3WjHDB8+w/VllDxbnYFHA4iuJWk5aoagFhDp2vZZBkjDvR74SINYL+0RUVxmF67qyQ
hJZIYN7/kEFMd5GqrSuujr18ohC9lM3kp26xFmKTrMWjElpN9/QJcssBG5vWHNXOl0WKYbGv6wUh
zoer9TXwLCVGtU2CBNCjB4vkv10CrZ2jrD2IQjza73ZzDwnXNKGC18mscnzWdwTdx5TWcJjbcM5f
wRl7fsE3Ky8JSFnz7ao3BayxV42ndb2IgG6WKNV4rMpasSN25MaOlM85Myb4oW1fDwmPzUbsxMMO
I6ay8Zy6bC2QTlUEgo273zbC2rYPRAYc+jXldZzwIE3NeWEXQTW8S6cKPMyI+u3mv6qwtnYdCEc0
DBENeX3dqvhIdN9MwFMzs2f0Yk4N9ZiNV6PE3v9lgiD5mfeeKkSw5RYNNIj59UjTpTdZ5hr+d7qt
I9KQkh29PsauWI+FGbp0PGPxmXBMaSgxEpDgBcfy7faSbdATrLTGfy0EndKHVUV6RT8YvgjSXYi5
SPqkG2iXgd9pqPPra/3BGrlXf/7ta3+auauYUlp+bJWqEE6LlfQMX817GX6CZb/tmgdOQyoYZYNF
ujC6dpiQBY2V4te0Uax3n6E1CMUKwVfEKsyKpvGlaacbFVqI0F6m6tRXcVNioSojc2d4tO9Uf4vu
2bRyJflGaI2zyWO/bEyAOo6FuMN9U0z8gz+XTtoLxAkzdHwLkJceAHT/MlSD5Hlg6JTIg+dxCw6k
DPr6n2KXvN5iB49IiA/M7yp3r9cpvdUYp5aaxhRZalmZsOmUf54duvUZVjXTg2zAK9FnlGIYlYB8
jGF4PyAnU9EOzQpqllOkyhB6ujH6kfAXGBsq1HUOoGLp8w7jFKFmanMmc4ZTw/evKA4NEMXTMVxC
heT/gH7JVOHtFfWMxhEpJbjdIHiXjb8rZ6NkCUVY0/dEcvu8lWyTeGmVdR6uDsyRwkbm4WhqFdRG
wEv3xJLB3QvcIsbPauV6T4as9yagoTLTR591XxPO4wJaY/Xz9cwAVoEMekKtwm6zCg6E3oTxSp8/
RrK0g5ZssDh+D6L+vJOAE9sh6yEns7/IAoKLlUMWRAHy3knppMHqKE8Ub9Pm9uPCl8MFuMFMrI/q
qXmUDaALC0D1bYiGNppIwr7H0EVshmVLH44vaEGPjHVJ7r82hQW0tkR7G+fG7xEQTFn6l4smjA8M
4hJp5fa4x3Q4XBa2xJf+82HWaaC6nRttF6awUSmTmD2nkl+5yFw1zry6O9z8vr5KtwWtZMLvf4Y0
iRe3uLpgEQECNvFc77SM37LkVrf8+Ya9hehg+ceBDAOMoAqN6LULu3dRugjZcngmZnYOx1bXznJK
3UdsveZRGPyraetPssJKXEvEjvOyu2NB+ul5jVa0rGXS8LD7eCh/X9HIsqDm7dwoUFIx9JjI8GEc
NHv0eyJrgrNR4vY8VEv8xVuGhjc4jH6yfXywv+/agxoFOoM6oZeh3et6kjTIx9+1lqRi42aSCMeL
099CJb4Glzr5BR0ox6BNG9Fad9UinOa2PyM2HZXacvDeT/wO7EsRDWEGxyQMA6fO8qp4ZUTa4O8i
3TfYsaNSnY0VhPPzZ2hcZi49jXwICuJ8+eCJ0TYH41fhKy3FRxorpDqze4qvBnjW43FRYatPRDjT
ftrxgr34O2j3XO3yATjP8N2uqPXX5noicJMsgB7n/XrEcwa2NI7GbCmnkAgazWsNWqtA0xExzl8p
b4siFh66nJ8wdaMHea//GkqBu9ZnRaVsZ3JhgAnffYC1GWgDQgavCS0/K/saF0M3rp2KpYW/xV12
gYXZ9aQKIWTJRbH8ZbUMSqg9z3YLQAlyv9peZJfkpxURpN4Aajn5qkLI1uTUSNVTV/j8xskl3heB
b+amTkS3wJcjg14yGqIRJpKGQQTcPkaPVRCrK3Sx9kTdJ1+93/aLn1e5DK3dOadHT0biM/UWDU23
+JiZdJqmcr+j9+MCh/Khlr1/rkvEcdkF/Y6Nw/qfNgIN1r5UrlxGp6lsyeNVaQkLK2MsAFW18t5U
pGH3eINKEP/J8wLDJ3GEryxhJ85BfFCdHF2fTRB6MDkFuK0f2x6VN9lAkJw6tFgrhvbc2dvZWQwO
GV7+Hqc6RWR8tqFpcEbZ+vOmKjaPQn8uNzn7ziuQFQvGxFwOLTPXyWM/B2KYCMZXZWAE1RwFBc4c
OZYVsdcZJAsZCO4XiwBph+M9fUFmWum2V8Iz1bYtNWHBvtnNIFyDbBatsZeswpojLAaHjHHdWgEM
KBAJKvIB97ycBsGqJNQ0oTHHLzYi2S8H0xrE+GVvQwPFl9ej9JvYYu4DBFGeqJk8o6vkyjscHv5b
PnZY4CabKgh/1NxSr+WI0bmwkWQkC/rT/ZT3SzTCFpRpOJbfCQMaKnIQNyFoFVX1q3PDVXKusMws
dNAjBYtRvo4GRJWAtOOQa99jpN8M2y94LZuo5cGJr4FHt24Yi8AcDh+PbfKU7EARzGw0OUqHkUKp
JBRL20hAxIVGXlRoY1iFk0oOo2fGY+j4LP5mfbTTtc7KXrhVanPPZ/s/3uBoOPsmlnVwZLpgKSU4
p79JpYHza5yHUuKZcIGoxB6yhHFN1II3mBCxWwZro8sLtTvUDuYQgYgJ/8Qbcnv0nFCG8vG6ZUpz
HpLmIK3OS4CjLD0K4LCK49yya1TEo2+D4gT/HeC8pztume7EQVZ6RA13/PrFnW9PMwAKolDoMjC1
n3oFbUvHB35f4g/AkSEPMnd2SbOsQ2jkEUxVVi3B8anyItAFMpzGiyx23zCHqnB2FsRXH9FwtMZ+
Lt4sN6+v1/65dcbTDw0bbYEL1dWa+lyt7jehHKvgmEwBm2w6hs0WiNAmg+oBye7GBYV3hN4U1KDP
rqId/4jTB4u+7RZvv9c4pDGh7+DDlT+SRi90Vxs8ZDWHngPGH4+9Bnb+aqkC4yTC3RNzJWIvyOjq
hCYyQWGuOJ9maBp3DvfJknLpbdaw3keQ4e0eyK3S8Te1WulKQVodiFY4hzj4h9vk1UCWzzafzCXx
pnkqvUvKdJn0BQzX80xxmo2l87dBNsN7Up9QX8LOICxusMOibEDYMKn545SlL4OOeYW9tgE314+y
gNaPCyCaKyRSfwkWJk4RmMtHGMpDVJ5TdJ4XCNgSKTOPHbaeBd6komVoiD/7zcZlkEGwSzC00Z1S
FhXGmsrM28xMYSukSncf2LjZ3OEf/daBhILtXCmvEwQJRKBhjz8HbWa+AN3GAUt7mFKm7VOD0YtH
jYTyzPuSqnn9b7ndYG+kb9507RXpdt4mBti/iLaqAw/AdAVRUW1ug02s+/iGWDfUU8pILGMtqcmJ
tJdjwjDXAKTXFZ0ed8XI9O/x9w18BKBhidiAsMN7bIgHv0ataPyEg6PEQrfQcYu6BVRknM1jwQrI
PMKqC8FkE5u05ky22G96lFvMrpY1LtYfAg1uI8reS/D72di4nyZ0+IlSlZ0CIXR6xYGX3Qu8OTjo
zOYO1DOSvOOmy9bYnSrFDh+Bopqn2RhGNkt4+OWL7Msq4OZxJf15Z2dpxIOqaw6H1O1ei2OzFhwz
bc+ReUNmqsq+8mCrNI8LtvHtxkDGDo5EO59OrkfORETZWe34NT7vqCjpc5JcjX0OPpMEQbm++U/c
4dFtAkKrEyqWv7Ihg8P0TmTFRGHInhO3VMv6ANPGHEOCFaE2BOo6mZcOm/eOftMgNJwdkxzWP2uV
oW7Hu0K/6VW0vz8UeXvqPIVqigD/azAt5jQhElaivwwTmgaQl1wf7RYa7TXyGkaTKPQgV1UJRX6a
wbRP5lrhqY6BV58b8YAPjwZV/LKaO/sudL6OeWb0zzDCAy77Nmrk+w1U4YRHMd2a+eztws/5F9gc
nY/aGf6GHxahFukh0p0Gh/y9pjrdv83Hl2FBO2aWv4pyTuMYoXxk239SfOcqeLI7GLsewwd26h/7
4aIbIqQt/38aIsQtPejd2goYrbWxyp00VO7jSvWd8S+nJClzE8DEk/8ZY2UwgXo4tlDL8znSD1ud
1lS0erze/0jSZzvn6P6pH/mTS0UFllYHSnNmp6sHKK6HWurFefwMBBgXU+GVZIt+TbkYiJz6FsB4
ODfonpRt+K5m9SKCbiY3dQjFkKp++GJPH6gpFlx6m53JsW1XeBSIquUoOLgVv1a0TV/adH7QscAH
EfnakJcwtxr5RgBk3yYf+C2qknCjgwsyFnvPvcdcKpzAc2Nf5ZjA/cnzwv3cxQLWYdEOz5Wzbmww
0xpFWO6gRcMX2og/flP0wN2LZzc8XTFRNWaBpVSNg5g1vrjGmo9S/JrLLgPtjLqw0JhEFXLcdBsA
3668tKPY9QwXzMa/TY7xqbbhr3qhiBrT2SnLzkLpVVRaS8EHnpnZY20KHMeK+PY9HSwxCq+1yz1m
e56vFKpS7CoJbAo/vu6EkcCodJVzQxnosH4lX4SVgAmf5BUJCPdK+ngfqfLqa+edbaKGV6OjmGGA
D38ZPPagJipGQ8KaVuJOOhX812sr0brJ3ON1jy4Qfl6CMlQ3CUw/mpSclHgFT4n/Q8ta9EpiDWaa
SFqw25hSG/imNuqdW+XW32OTfi1lsgXFWQDkSNvziKFKD0xnnh9rQrao+JX3jmjFcpgwiGS5tvYb
fBxqiq2vJrvs+HNam6ddg7O3ZkpJdj7fu+ZXwZ5KbXCHBbUTItCsfv6ZJlZF8Vce54CDhb2prGfE
0uCyXpFUe86oEq+3RwV3nJA5jpOZIOAR2XkgQ37pgBFFgWMlpQfxYOROyuqOUhNN10BHbJF3asLG
oV9pwRcQ0SQspzBnz1W172rG6WNM3niGX9mXDTARbhaIsmOKVVqTJIp55sLxkC4lc/7QJaCDSSfA
AvF58IWjw/9TYrOtNbvZ8KW933duYVBmRlEz3lO2hG4HlahooHMIE1iha+dlqBwpA3CDRjjA10ku
qFUXixnQfdOH6Edd68FccXG45rNYhy9c9t0hM30bYeOzt4fmAe4F0kJvhog1R2NCEscixL+ZsVpU
ritSDU0zx8AL0fLUIwh9ceBqfib7ltAfrv8XuwQkL8Ca7xqdCAs9+tlZ6g8F35rT/lNy21WV3+9B
6bra9+IHz7tUuHGEcDdthC7fltzmWSzc49rQ8z5uvFB5KLndKPf3Kmu4h/wdVK+uOR5R/CnuUH9Q
E+UER+X0cO03dG5mR0HC5LM3zBd8ocLYaFuBA23Us+fkHx/gYtCxMok+mPdy6jcrJ7smSI54Y69+
Oyi+1WTu52s1hWBgf5H49C+kHx3jnIomyn3fTnOaycIGTRFGHr9jnPykNRGLqvkFL/Q0Tn1PlCsN
e9A50vsCDHfHgYnfid6auiWCxa9SiXV78fbNJePbEfK/cfX6BRAV8tXn+ULhy4wtTFrQYcTM2ig1
CfBjPM7BOaBvXPNSzOnzFBxSmqsNzbeuSXrSFDCCdFGeWp/3/xijTbw4Qa5KXNiqdZolayvqNi9l
KCQEi8ZL3f2JcrGto1mpTizJS/Vy+NHn6C4wUNI39Z/2UVypXo4a19HVMUugCPm/+djX65jv1tX+
R4dptjrXvW+31GuK/XmAymTo0EYFFzg5CCoR3maN262gF3ktAE63EwC57Wses7z6aH29n8n0vFAc
CCgrQF0YbcbO5H+xHX+Awc7IM++nHssOr1M+gSxC7keauIcP0BUR8XyNYaDoCFcriACNKBMZpwBC
mt6SJSDhM0jSi8pY7fPiylv38ALh3df1EYXdWk2WvCqCyounEt6sjojdKAN3QwyUfUUy5qJPv2vD
XftMHNuev9TCZ8JvAh0L1lIldDZlwYq4Nf4oY8MJQx8IzQdgwid66E1SBsUpeTHGpO1NpJ8V3LbW
FOU27PRmMg20lHhu0jSGrSSK8PGH8LqeNDNmeQFtbA1Mb1651v6SVg3PDe94S/wyXgbPnT4TnDOK
AYum163e8b3/gwRNnp2kFvIUVHevwj2eir46AHZSLV5KYeIQLCEmPqyzINjF621RjdV0D+115CrX
bDD/TdbqQSq5BX8N2NpM47oVWgTe/Ahk5D5DIXGoQoj1h7Iq+VBNGbp50r1pzC8Vd2ZAs74jh3WM
KQyssvYmnstbos1bwUSnz9wivRQ3IugHQxYQ2TcVv1wWVO/SfrnVr87xY+pZLs/rv1c8rxPsmuT+
nNASzf777Nrri+D7h/BGLeWioU9jMIsiBkzI00PYndPCwCs1EzTV64ayimtOIGR7nV3sQXNG9HZp
NPc0Kp4Ul2lZWF4ps35LeoWWtcvZSlXC3L4eY10MAvNFlh0QDtDJOmtARaLxh1e5kDeGU9SdZ2ht
4u+BPyYFxmL8SD3MSGogLEhpwgK22Ojh9MZ+j0CrFigo17yuhqVYWrghI4ksY3/gUPHhheNrHEab
rmTWA9e39qVK4iIySzt7VG47XrxlHZTim49s7435UGcJF9D3e7ZcLlWygSMfG1T1WQkokT+8Kk07
RTbULwouibwUQxcvP8YpCv+wzvUsifuWSRMXSiT5dLsAt0vLtX3vFQIBUw5h/C8k4t+8hQ1Cn86E
CfnvCBO6+Pshk6aapmZMDB4uiMLwZcU2N/EmTbCAXit8Vl1jiZq1e7bYxFC5OssHLuQx09X3exUd
eL0GCbTbKG6Nle3XTGv30ShhwChNbccWLP83ZJUMoASRloLeZ+VsXGQTJj2+TC96Pab5aIbYKJwI
FO0M96CG5LMapia72tDUrERjNkNmK6cuQumxlk/dcxnvu/Rbb+4vpQo3TA5HoWI0+2O+TdLuY/RY
TMUM9vdweCq6S9OgD/TMyD1OEaETj+zNgpZ1Y2OwSCj1+pbkQ4KjNkCVGoqXjMyFh669WJhNwdjh
FT6s6/wC9jqxO2qYKJw/vhN8t6hl/L/oucbUqeBZ6eAl9BrsEH8HAPkLNQGT1+AVKN9ORm3tqvKz
w+RZZOVlIW/Sx3b5F6F9tRhA0oLC77RzBBajG74485rffGA/WB06L0vWO87yXdnNEuP98GEfj/RO
itn+Q+btqiD43VlfKmpnsoQLk6qKOyY83hxqn3F7/FQOgKQu0UZRWa+FWzCW7xd/42P6hL+ECqW+
D5k4+85MWPnxpbc4OkGUHjHLAbhOzQmdtgYe9LhEJICh93Cr0Z/Av/neHmXaI9SqeztzNVPcRJEM
OcShkDbErcGLxoJ0NndeFo6K02yBXfcsX7RdTzOvpNxBBr6tjzYNg2Bv5ufnOAqTsUUx4tacFeIh
feqf+fK7BDjXvy/OPLPmJ40qesuTF+szVa0OBojpGoqIWoQzG6XP84k5Y/u6UA7Bl3Se756UVyCh
rimY5fdmL32LEH9ldLsFqGj2XsPts0alz3lBz7YOrLFrUH8CVM/1ug5+MJdaqd28t1TMOYRs4xcR
Hc7qFXOnP76vMYiFACyJa/gO3wAkljUXIYK9e9s282ahW3IngJony3P7h2ATEmD0xuhy/goedHTS
9axhMapCWPA+SyFwQkFdKBO6FeG0y4X5lB5s4LA/EMYLGpSpeCdl0fvb5tjNOkHXzHn3rPoQtRwl
noB7VFFuTEQmVSPiTq/rl3Qe00QsgpE3HFhFhjcaosNPWolVQJ1cbCLMaZbyGqSmX6EwKY3HrAMn
HHavNkAXiUokVTGuoeze0kg5z9dYDGyD8TEy1AP+5/cY4+94tOgTcV+67eE8jUVmrb23LKBdwOkM
MO2lE5VOfwAgboVoJaMhKplKr3QvhpN7vdwAAbfwgvy20hETgBWYnmckjofogU14fN7XBT0Al0zA
qly0RLBW0+aamGrAE0/Cv9wZhuc8Dl3s14vfJYsTGV3yAcbn1heTGcZyF2T3KeegNmshJk6aH7LD
GOsytZ6TmtEoD0Uxf2vgPGuUzwJz6VdTkq+4zJfry56OJbaHhfTeR1kNcktk1V7MVAIWaozSEGny
NSFTeYxG8+Pvo2GXkeNdpvAJBVOUsrrhbfKsrlRNRn3BzlgrxZoLYTURGcdqvwGYn2ZsQInYAykX
kXCRHnc0J4ErzpEwGi8aXEt5HgUWw3mX0dfyCOYPUp15UdPJpZC+0VCcQDi5PbfBZ3r566BCLLTK
EtXrdf9ouDX9HKXeU1oZUDEpDqOk40Zm3KaT1XjaTP/15hgjgGmqmcaNYcA/3n08XIE+LbjTRkGk
rmOnExsA6xU3NpzkC7n3WU6KpKvOc9enjtD8CRzedt/8LvNKBRAIKCfh2OKn1f8I4BdoL6k1P74R
+R655sCLJyvR85p4BkF3GuqM5/fmBJWp1Yhc1roELnAquZjFRnEPrNXvLjRVOjiCvg0r5u+IQVff
Q3TfRDIlHteWR1HE2xLra7L3kY2vDJmzczHC4mM7HcZaH1GXE9dbpcFF+1n1UStOuCtVCV0QdYEd
Vi1VCzCu6SYS1jJAJ0ASXQT+4G+bVXF3GG44+hf9yrMyF6TGz0d6kQqFi2HVfbWWSj2ZTeiq1ir3
9YJ399tecOk4ff2G0gnsgagz9KqTYyqT8opvi6zUcQvj+6lNI0BDl1x5Xax9BICvV9PRH/cAWtPK
Rh9OxYdKq1D8duKLrO5AfwYwuBIMsPaf7UMRXzLEcp8sVW5pm3m8ZZ0vFEnHLSkVfWGm5sDrp6hc
9RUWF3ta2gOiZv6GPZVTVOor6mQcIFbf9Kv5ST/mV9t2b/jgza2i8iaiez+wJxc1PhsR8/GlH8mV
lih+VpTWJB6PBPj4CLJaAhf1/Io6ByRQAi1FzXOqBDqNJPkKP7DOCkB3acwjZCbQlLFcSBgClE51
KpCavQ9XT2a/7GemicQs0sGTN2wbf1JZNlxOYRMrym/s9fbST0xcbd77otOG611Ril0aWaAvMUO6
QuSH65JcRLmqztVG5vmT4y8GxVFOrzF4YmzW5m07Qm8V+Kn5EkHD2qzYZBFhMLdeK2UDetqVuiqq
qkp9FZPtszrVU+KagfJ20QqapmVF98RjYQcyyc0qRvnWkyufTYSNk5meIjdkLqm5swv9AddmQBaf
npb6c2gv8N3WIesoDtsGvliUSt2bdOFuiYS0qsUZ4pWqqdfYvFJmuTg8vU/XvfauwP3EiXuUT0kY
BxYDc3WB1c2HqL4P0it7lAWBsUc6YYfuCeYeZ52AMHShGk7SxblLqetDkbc2o2YVeSngpOaWtZwx
V2ccODc1iajPyKECo7gr3Leeos3RFi7e5z4GGtOLyzIQBeEC22gM6qS870gIPLD2iogee11d3ARZ
fSqUfTBjrvmG+/70mcQ74tl14pPoEYnM0sS3ga8v/Wkv+Qp+zbgE6xPKsOK+C2ltGLkA9GY9VkCS
REPihRTV90czKSorD1dQ8N3I5y7J1qFN0f9/+p2cusK/K7YaqTIdVhWpSyiNhJ6yYOi4k7Z0r8GV
vtQeZSRFiWaFpdFOixdxUUZjV1BRT5hGeB/8QUrPRB8DdeS2AxQY5z/RgFo+hullPNu4fuTnQzzo
pzZDofAjt19bHVIpz1gS6nMKtZrvKp1mC8IGSHM2uWgGIT4dD3pEEeZEFRVxBgKISffNRo3YAJm9
yR+2Mzdd1xfSZ6CoJSB+RTvo9CqbN0rKeThTGvnXC+BS8jd7rfAGKVS48tNP1RisLuGJB+uUDWQx
V/94yRbm6TpTR531i3claSE/7EgoezgZxuNRh0TkgP3Y9u3ptvH9ZQSoOJ58m4vGcyUp7WlxIwMj
elBgR33wqhb1S4OOYtP0UIIrqGYxXYbg5OeFG1ZPWionFNP4Oubodec9/a4RLhcWg+SlHA21XXb4
OMENuAVGFH0tzu7oAuVn9f0Z0mrWAlauKvQFz/VyCPaVtO0BCEhBcxcMypPoGb8BiKIifysT4wW3
xXOte231Jamhh+hUJnzOitnt1RC1UFx1rTmomzyRgiqPI41w2Ff+ci/1NmD/Nsi0+LMHdX8/Fnig
fNni3/c5A4ukdbT64E55CXKiA3hW6e1yBUuEQKWxzT474H6/MSzrpMClH6yt8Ju/nNrG2cI/N1pw
Y4ume8Qm8eN2aglAXz1awmmoUstqSVBZ6pugi6yTHP1F9hS+N0VbN6MBOPU6ZZoIBIwrwXoxNCcX
PkjyppwBhr06YYh7wVBeGPRTGk+mSIsfCFTS43uDymCApF3PuoeR+K/uV0wPS640Oniu3p8HAN12
rdRg27JuEE2x5HL/57IeRlYrAYpL3gq0Aqc1kmLHq9vD4o5244YuFVkr33XKPadbMfE0T3ihLRBR
FndWyQfdbY+4iNCGrFZkdmaOjKH5Iag7Ew6RtyADTODR7oCUo1mXf+RUuoD76i2ITgmoslFstuok
KPQJfmJUAGNlHSzocfQVD11R3VYMn66XUyQ6j6eIkNURgLwrwUomedY1JgUoTZR3HfN8LYYqa1xw
XGghsJAPK4DfoNRdqk4cNClRxYWZntD2z/WW9KiakWMKbUrQxG/VspYhR/YswGYCltSzQTuVV7t0
kII1eejgfF2brTCkYr2sPvRIaEW5MEFz9XR3s4tMN/01aQdACuB0Cp2vE4kwbRBIZgFMTHd9h21C
sCLV5AA6M+WyUroTNyxDieeaNVsf91QrpnpV0l9MAbf2+zmewp0p6vEhRGPYj/14VRme0oNPaA05
zI1k8EgFHNCrO4qzRtnyR9SgZQHAP2ih98ar59pN3+Yyz7+kaV2JHB67b44p4uTUUSY0HYnOjVcH
c6Dj4Xtrej4bWCY/VzPz90tIlKrwcpDQSHB9n0o4/WRvEUk/oYitM+tTEIa3XMb77hkKjlM6Y3Yy
Tf7cjSByY3BYEYGUhEgPirmXMfaoRfz5kWaSzqT5Y8raOeNLOSQYon5CPJ55aJFjYzQttKwdFJjp
7kRsQgIIxRH8DCMXCfqSZp2GBhFWvDf2SeUITBn8cjDdzE0zkRoFSvCuUohBAkMi+Z7ICRoeIuM0
PviURaw+WTDL3y/u5/F+jCRFF7x+dqGkZcbPRbEByvglqgdYwWIsdimb9e+z7zV1uOznj+QjoCUR
hD+W+iQw272cbcwPk8w2FUfsVuVxkNy10J5TBxoJBXT9u5dYBV0AEoHVUXAPv3B5XFWskepYhlXj
+sR/8YSGq2LYpE3TzDZN7M29NdfJ4ZnTtyke65wiKUpNG0/KY5lYcnBcgllG6nK8qWI6onW4yMX7
8yLUDHV0p7EKfpcMCddGT5xGy74GM9w++4JGOXBmxKCgqDmJ1eWqKEKQqN7gXooAv/vDBlfYfj7S
Vt8feMKxS9Ln27T3y8xq38ozryLgFVzgx/7339eb3tkZRRZaDBND79eBhV/HoD1glgENU3zx5euY
7uteGWg8rydEJnvtbtbBJAlYK78f4EpH1iTskNMkfbZR0wUPM3htDyfZiLynB1JPJLxKhAq0/F1T
6kNoxyhkiduUZANrs6mUqTZ7WFvnOr6ZFqy/I3NCcstk2btDhbhsnHtrIUIT1nBd+gvYTDOzW54w
kqX9ZBEY4LaPAGDXyLuFGeF06aXsQJkSBCkyJXzUKfy1HjQmDchh3KpbWmbPwD0QAFRbZ7lR/kAG
J7H802USJg+wLWZpq6q6JLTrqXzcIMMmeeMki8w+HxucvtAx9vUJUC1qnBvfovKIAgLH+NPl9tcx
AqY0cHs1IgNpMug7/ia1R+yv1SX1LXX2XrorESLx2He4+Kw+MCNqKAQ5rtmyXztyVhKflo0OnV3A
17hYUC/ZFo9zS7PJbWdl2yeDrc/t+6tQjqDVgAHASTNiLwcz+p0lrySZl8JOxZOnK7pzUeces99d
aChk8rV9W6ZExF6t4w9W9gBNnRHyGAKkXhIaCPYQmS06qtKeyy5+0Eoacv8nvJCbMOFvt7Zw2CvX
FBq3lInWLG1qxYshApUk8WoineOmEL+mnDtew24ie0ijKQC0nIHrGIB1VnnK/u9RyFaTSj91ETwZ
EvhJzTSAlt73gCBJzKA2n7E9FcB0cSGS3gurFLEcHI8tBYtGlufvvjhqs+P3saFKjjOKe7WIQ1XZ
BUO+MEi1ST8I9VH5SrXuTiABxaOBzWC8r27/W9mhR6r2jErRyO6/DZmbklU4PSpsEa1PoOfHwdjX
F/JjGVtKMBLPO58b55kYTwa6qYl5a706VVJ4U0cSxaEyxOUPfVr4a8YwglW477yQELETjgASom2s
ATYU07J9LPWU4SpR2KpSLzHJjrxPI4UI/YrNhC9Kyfwm9eUiXpCe/s/jCQNGQDgti1QdUNbr4FFy
MXXt7R7hMznP8xRc2L/Uz07JatCDXGaxI0yKo6USdnyDcq3M5vM38NF08Ya2A91SE4M3vpN7KkBf
lirq52LfuoISWziEb0etXO4XI+7e24zpj0Z/3otJ9F09Qc1ClJm1UVbDEPROdhPmaYXJBLNabmYz
dhgEtgLG06tTYdQVPIg+oCDZB/mgK9ufjZ2mFGyKAlUkezlxDrfmvIHkGsxeVDG0rnrZ2wNVYg1f
kMdvUUqttIUhrFo+etBT5403E8GnBKmgKK3uTnutLCLsSbAXeMbF6qlWckpTJFO0OKpKc5/1eRdB
TOAwXhscVqCZ2njE/XjHFzo4klmcZd8FPg1GC6Cb3E9tvJzLBqKBWxDuvwD8VShHlgqGjWrQx2Bh
TPAL4m3GmabVjh/DstEH4e7YFNidNoHdIRPNKHjINQhhY/210/WCibah/BwDu7FqyfJQT2E5oAZx
zKGCEP97ITteSAwxV8Tv8srYnvuC9UyhGjOeB+h+RIL2G1azmN0BkiVZ91GxwKoE5sDThcgHjgoe
hEo/e2wNCKxYUuALOu1RzOPR6VR21gcGfMhTPNzbbiTEW8xyfniWspxbp7kvKP2fFdndxQA2VGFZ
84wK+1R+aExMy7ydrRs+cIcJc6NIa4I4lho9KQA0QVSC7aK7iXZ3DyFdHzOI8bJ0LNwvQCoAvAs/
WGBaBK31u35X6huokWfcB9ZeJtpCOs6YC457BWqChmLZq87nZScKJdlcXVkuHkB+DziN8oqmLubd
rARtVK2SvCI51TQmTd3FKOAk2xxHSgOwSUqol7uU0KZdyk4Xwl7nFEVT0Mho/W+7YznAhPjxijgg
3UHqq8XSS60+HBuKFP4046i0s4IpwXWZ9UBvYLoVAPdOxEQs68QoOVRdkuLYSEqmidfa3t2BC/oz
Ms3NJe1yZM1nOygmT9zSJCXAxNX3xslY5iFTunyo+baaFedKwTeLT3RX42TCmT7m4ofiSxlzvHkq
0id6032VmGH2+4dMh/H0EQRgbghCaT7EzR2LYaDtSCWoQ60DlDk6B9hHXGpgEnUZspw1navVhXXm
zFMUyyT2AhE1BkGKwpPVxayOnwTOfOHoc+howUESKapY32amIBkAf0Dg6SeTDQNdHsPPIzJ/R2Gw
o66H2BofLosjWDu4aPKbkBZRvhalLPox9hMc9WKsj3KdZFYW7NpVy2Wcy5rvhaKIYih+JVHRjN08
0OA5RZHbTw12sz30Myp0M+VyOHlJHoWl9IlRD6LrYfVx+I4+5ERHRDc7TIJPL8XgICcjyyL6fnld
yUdfj5iJIlnGt6rHgXwJShutPaH9567qy39LZWhFirsDutZ292rUdJdNU7zWqRJIuzYcZ2i5FagW
3AaqzK+P+2n4rCaIxLz2IpBnQ4XEs0gVeiSBYXXtJ9CYWP8s2eBqpgdjvWfeFj48pbLd6Q66vz8Z
iXk64bEfg8gKpC49hwxF/jIkCOyclm4FLafuZVcpnQNgfCh0Fb+Yct5jonyFGDFu97J3y5t2SMYN
v2DbgMgjtb9blPskN7iGT5b5DaWqcUDcy1q/Wl8VPe9bi5+pH1ZUvRmTeWbZir+nCH5I6XnY8Vr4
LxhU9+lY94aUCc8xY/gpd7TB3Yn87nNYTnl2WdmVGdP3kD13LBKbV4FXIs+c2ERBW252Tlyz3CRD
KUcutlX1Le+bgDnDxvoHpK/ybKs9WCAPQ9srJKfl89E3S3dewjTuVvYmga0axbRmqiXzJSmPzLo2
stTX/89AJVXDRJskJzAWkUR2V+pkhBrHPvEICsf5OZncBoQbvgUPFHlwYbtVQ7MO+FLYxvjG6+Qg
m3vt6ba3VCaNO14xMVNoce9GlR0M9EK6m0zItf5UfwMPQgnco/deEu17WUgjwWc4tlp2CHdGxK5C
IuL+gombs3rnmEodhJDILE0cLc+1kc/8W1STOUQOvNQ1BYaXumvCDs3oQx3GDhRmuBc96Abcq9hA
GCvTKMcjosF0n5ejSxKDmCr35hzZbQ4V6A+7mdIttTjpISxos0U4NmbwK9J11Jdr75DmIrZluzoh
8wNEpa4UuDwDKQDvE2WEehtxTjvJrcaP+QtWfB3FRNq47SDIWvdu3yq3tdxv6ahgeMrvrZDGOikA
CUdogR2TmH9uSWgRjEXXHma/FewtyxQIOrAPNwo7kfpgs8Lt8xrJKTt4f0SdF3/IS3Qf2JLFGE+J
liCG9gps5lwLEnlrtRJBLmwz05KsfBHj+oJkhdTQbHT9PCliLb4Ied46bdZVSPgUjWXjxRT5R+5I
s7C6KC1+5RNwxb67p+Mlup8pU/ts0t6cIq21edDM56D+be9jaM4KIM4lj+LlRfMfIvPJh801wDhh
IwdslxvLzO3Lps/Fp/7sH42sfMC6pIDEENJeGKmNNm1Tzlh9v8D/GiZTig7PEhA29BDJlByBKwWf
j9v99WxopNZrwVe+H4jWjjv+zv9S9LgnVLymHcY6aqU+XfWbd77lPIRNgTJbGLw8yN8YMIeat5aM
eQiQHpt5UKWfukKz6zRrg6hxWdTb4a0uYWPmIlpyq1x5SrEh/ymJv9Ij8MJtg/yj2y544gMMPQuk
v4f18T5ZhQeBe6nMI/uRidlLPtqiM5QouWBT9jIP3K6bnLoYS7Fh1UGw9q9usf1vveIa7XtCvQcf
eDbAm+RMGfKwX7hbSiZk47kCp00Q/RLMvgRfxyjBwpcuHL8tKybqCjAq41z1IoHZ994DrH0xd1S6
+nLq2XDoJBePuCxPEqwBzFhDGuNEaNk7Mb4tePWCpJQGuS32XY35wgOaJPVDpc4rXgNHYsDC3TH2
pZ4OTwWL2lutqTOPffak9pprRy6fwYoP13lBObIH942K/MwpsA8B7Ynoro+bwJkn3o0GYKpluk8a
DqB5cYlGJ4rcIN2IhM7eAdh0miyxwb7D738N6RJJSYx4NrCMr+V0ntc5noj2TNoIpM3jPvxk7zxq
TxOzGNfSOKxbsYBjCbD1Y2KxSE6sN94hO6xwpGDf2W3pfREGBINkkt8ZAglgQfJyiTlj0gBqGcWf
s35WmpLAcMUT8437tuUcZIcEQSiMUnDZQxQgkNrbAUKQ+NDKUs+xStKhVGyUoOVBZfLJ2s+9EPUC
5fU0e1N+JdFwGUcJQuJO8NR5MhaoWh8lF/BeH7yV5+xpjKigiEV0Ug/XPQ4hhycuBVRzus9d7D7P
pe6XXZCKZAW9UwPiuOKVl9Rq+n2mWDgxLyWPmAM50gYz1JA7Umcqc9GaPiB3E2fGANCDCHmFqTEQ
Q+7wNJkm1wPba4ClOA/ZkbX12pI7EE1Dk9Ou8jHCn6ngEommFXG/tBdonmfJ4d4CFT/+sp8pqVvN
FhAj54ZboQfmkxFIvM+hC3Z3tzBkeq2xGykxrym0nsmKyyH+VuPFcIIiVDM1jD+bcF6R1Zqa6ou6
f4HQHdkWS4ns+UI9kjpehVKaSP9o5LZCFg3zFyPnRFu9B5itLGQQWND+29SRyudUUsK5rUPnnSlg
5BQNhWRXiSo+gDmaH36ifA2pFBdwweAhWbCkU5ljyDiB4BS5xD1lhIHgP0iyFd96O1xcoye5NFDb
r2X6w/6zwPEIjwSzdt1zKr6yDOVAcS6D1xs4jXySC+xtfxs8XrvJEOiP9WWr1WJhlASiHXQTQUau
NSeEnsFwS0xOBdQsoW02VLAfd9JNCm2PFNu2rO5nXnXq6G2470YPlv9vLqKGL2r7Pvogcza8XanT
I9xsRfXIb28ukmumWFIOgjI9E4esYBxSCMOHZ1fpmv35LK6G9c3Za0MayoHrHubiV8jV/lsF4w+J
0aoNMfbNxbQuKAXRWjcqIg9p6yTNY/VDqbsFpvJXQUaBYDlrviHCMYy6Yi18tZ8Ce1QhxPPMEKPB
ldM19VzfoBfklTS0znOA1ChqUsO2kOGxzf9vbzrVfa9B3Txfb6dS5JWC44US8+tfpDJbFFbuXJvh
K0kSQhfdG8eUi3yiyzxr2Fa+2D123KbFsA6MwLcCnuMBSCPgROQKqf5Vmj874gE9ScVy8qsAkVI5
42U64ZM3k4h7P9c7vYYxz+PTJYX+Z80fxF4zecP82cQYkuXFEpkL4yaN+8ws8TZrlxImjlXdVTHw
WEB1NGm0AMB5LTlKqEQ5xa5s7DiqiwjfABqUtNnPTTmVsj/5xnamhItfy6JOxqefd4sDNzIjief5
CghAajpgD2/hi69HXumJ+KJFwh6kWVWZNPvLqCLESpPA01lIcOeCI86lFIngxR9ZJrGXJg/PyM5Z
n3FuCKe+8mKDBnpXHjQZDvgKOUmG/SpgP8xklgZJp77q69hkeYA/eEyHtqA/MTYP/3Pc3j5QMthp
GpulEFzADpYh+l0Uvm3lxxgZSMkwTCQxXLCUaduHu1elThn56zc0vfo+YsgtJlX2n/dpwVhQLGci
FfCPW5iVrB6NnuA+LvbCLr62w9neYyYDfE2GClxfvqOWZH9HhEAKzGijTsL0ipzo54VdtehVLvUH
XIeccWj/NlFoukeGtFT4GxFwQGvlLcwI045uDzPUNlvH6RG4DY3qlgiGdCGs7Jjo1PYLpfNyR3zO
u6Gj5KwdYvfudjNbCV+uid53uY0poErjfB2RDwU+8jAUy+N3ud0d+Cdla2urFOU7a+O/o29AXdlM
kwQ7Yy615E6qLXuHRXVy/ZLAo1ibIx9BjA9bo5cGdyek406ml8Q+TW6ZKvG8qfzNd3aSXfJew0Dt
/FV1zOjDqyZRVzzG36thiEdM67t+P5sRxfbbj4l7f9h0i+y5Qxi2g0W3g4gxZZ1eDnCocc6y+fSZ
rKVN3lrvsnQkQtnvkX3bJzw7yXxSXEVnecaYKb03dAOrTR1hTzI4sw4KB9riA9i6b6OpLHOgxc0M
9lBeNakegE+M0YsIR9MEs8s/ctXLsirHa/gsB4z1sosY+2iXYwV+eJCRFW9c15nQ99po28yA+4T7
3FqXJdvM8xlIU3LYMZ9y337c1pk0NdetzWBQVg1OOrB7R8/hUhUwt7zmpr2SCqtnIN++37lmozm0
nq131itpUed9Yufb0k0pk+FUPl/x1QoJtvl3K14rlCEQ4OS0Ds55uuSX/i9mPzFO09iw05GX+9+G
2gf3Noqa8rw1Hu7heeDH5IptqVlRCaIaepFwfBY48Gu6aOWVffctvLbf6uoe3oxj6fe+2vK6kasw
oOogvVgoeWt2f/mUHVPDfdr4GH/v3tsd9Ggpspwby9u6iSmz2wDOOYerwIRjiDZXHt+N6kRGt0Bn
VYku5yX1v73pc+IvN6cJWUz0w2a3fIGbS6VY7vx+pAloapyMP3AAF9KfpV6MHbWq0cJzVdw0dJZt
bOwrOK/TUD7VuQzU7WdhUkUUtm5SaqYBEUZ8q1SFn6uAX5kRLOmdOd7WDlqmnITmhoOx1DSiUhK6
ZTURWnNWYf1SkqFrPKvMj79hW/OVte4wSBuUDYqV6PbYLoNDUPpeBVM+c4/ZukIU29jGedJhjKES
URX36BTMypcNiZSOapue42Xms776/7KzqM/kCmcT04hEiBBSnVMKlLF2VilyZmQENTj4uPdWewau
NsNUE630Lnu2MPKViR8Wpl5Holnu+ErH8/yuWdh9U7K/95kYGYTyMTULk7O+xiBWzHXg+5MgckS9
LPUqeNtd8CHBYlAR8/PQx6ZRIFefssgdRBe/EKR0mcJAfP00nYNOqT47hg/1qJ7B/1pgJINTJpbn
vACab209uc8ekC8t3wRN+hEeZ7TkaRXdUIEXups7cV6MPWXzW/r6BUjJ+cs949Rk3LP1EixMAy2+
UovTdg1bpbSPvSlCFLlKKOmcMisPFTMsNwlB+nDqhf5JgJFUlMf9cyFIh6iOHQqyoA4ea1yBdGbe
4QshkfzgsqsIrom8u3xqGuo64TpcFilg0tgVqvDYZe6aWtgYGMwudXnZwQxmWZ96awVaSsDsuzQR
De7Dc6hMjqmP9gYLCL+UuMaNdApselTKueXOAKK/AdbySIYpshTQQb27DnzylzB1smt64Vu3VTld
A0b7LhG4hzf1vUaSvty0PCa6oPmb5uvsJD3JLEOatZp3WasSW/ydSW+vkYkZJTb2mS3LoFpYnziz
2ZFYeC6A9KDuT5qirPayaxTzWYuxoNhybyy+a+ZODjJDfhs6E7RP6DQDLhRam2L+NuwaoVfyDDoS
Rs3ocEK2Tl2Wq/RGUQ8SFV3OezJReFS8mbAVXcwv2nStINY1/GaTL4ArmHGv8Y5BLpAXN7JcTH8V
Ce4z+gf1YCz6Qi9GDf8o+I7GKGB2nQWv63l+I1b+HS/nWU5Mj7vS2HmxCuKET7qyb1wMrYgRmKDJ
yQESR52wH4LLCjjs55HpTOUl7itE+RF+r8oTH3BndHeGuyPa1sALLUzlXT+SQGNs2hHI6TO513sU
+uzaHJljmY6FilXxPd6UOUTr8IhWshohxmXunhHhS8s3qxEIRSy5pu9dIuATUogk0+9frf+Nj5X9
DFlq1X8QUdEetSMNXeG+lDQcVilU2wu3IPbWK7VMKgiasM4Vw+EwR1yyxAe+pu6AILI51NuCRc2q
c9Le6ilczBfzDlxyYytrJjjC0/LwIQSmLZl0v27M1eGRc4yFDHHDrPouR/hlukAGSdwRS8Dif528
IlLscNhuv2bwdp+VOWI6x3cP0GZcMtdlHAh0Luj9AtMhYAdMhWuiVL8zXeDX+dmedqEiGAXP0yXb
PKt+WnGpO4fEG+UBlCb6fwmbkyDVH+yh/Nlh3YcerCERa91bYeZK5v9Ibs1D3OjN6kKTVWMuo0GO
1ZYw7QDYCGWiKJ6Pj1Ht3IS/yW6PT3r6XJ5zv6O7SBjpVM0TCbfYQ3YWno98ZT6QGO383Wzx/c1C
OxE8NCw8Si4cF/0kci/YZef7xAgVQlBMIvfanrmfYsRgCIKpj+MlyNTnOXmoyMStX0DaM0tu4NdH
0U+hwCw0LltrnXlUjUT7huVtcYtRhwnjwh29UquPfQNzAkbrlTI+QVGSXG15MOdHcNPlXw1LnSkY
Dh5d7labzUtvZAQIra2QdQPCmFkiikS1YKXVwdDju4dUf971b4JJgtpmuIJNIuS5y1ujf8DLpI/J
IP5bDYAG2DwtsjR3NkJQ9ERtpiWpO/doUVbdHo0XEbOFF83MXqZP9M2jSYkoZYBPmSD3h14XZyQo
6iZLK0Z2y3PUoo4E2ED+2rvIW8oDCJSAoPqzZ7WLzkHXYf+GB1bpCb78HXjY7JCc3SoHIodlj+bc
VRsgvWHQ7x5p1EMzzQNd53cW/tWjLBFhd4dW5Zy1Mwmmc00IUJE1SNbn0qKycAOMarGcQKpofgXQ
UcEQRo0AWxsBCR+pNP3anS1hH2iSHZs37NeAa3gQf94egxW9tiGGo/ktponOzWlBz5SFKg8cxRZM
h1AArxaot9TUiGbggplIoQ+b/YklWj2nXfGfOg9IaS9pSVgpUEIy566OTMcXdbnht36/Og97aRDq
40+qwGk/z0B49P7MH0BI7kCgYxOgi6/bLXsCUP+iKgKi4Afg80Xxb3JS+zfsGoSaGx+ixtSMUbgE
UQ8mfnsOx+s2odBK4PIQupFgNjsUcePD8WJUSZNxyvurh7gC2Uz2dl1kkGVYVz56mu0Z6OK8Im7C
YBPbf0ir9o0jBOM/mcxjr3L1hbqxKgfIRh0pLd4QuCQ8o0dgW6IFFLK8+75aTQnDN/3th/dWTfE7
L7uNvXF1ObzLDqwlFQNu8bBbUx2fpu4wDX1s1BPzhPS23WAeM1+BC8PUmWCOmLNLHgjABwaXgWJb
HZXFxTUITXBKusQNS9gPP5CI9lnfMDNtv1MYE/xw01Y+BG3V4jaLfcADzmyCDI+N1IgQE7L7Rgix
cr557e0JsMPdJ/CKQHFJR0cTqiAjaXsuXjT0laeJ0uLdfv/xtHohOiKNnBCYUZzpr0Ih7hgH0BiY
/N4oTapmliyh38WZb6RQIMphqaYL8x+T0oH6jmFXt9jLNFTpHh85zoXcK3WJDUD4EXNhxtKQTMF1
qAxkWouwmiQx0P9pGANITlFCee0RH30aJRAjH4gB2n9F2/iRZFxJrXYW3DxvWi88bBSXzI8c1BiI
DkOjmm5AC+PNekiQ36I+jEtGFHfmy6XD5pqdpiyUMeaFgzoAupVMvyWn8gL/zU+pdicZe/WROMG3
F2GKYabnzWldshDAqBOd2ix+v25vs7mwVXt5XdpuERCVwt2j3BO8K7LmyPyJPsSV3xPv9s3TmLzE
qzviUs+rnIC3SJB01DXrU1jR4iId14jRfvbx3nDRQ1kA0pWUsC0tsa1HBf48RFDe+U7LlQ7kZ7e6
aW3SMp12hVsx3DqHv8PtS7e48WEqfzNSkoD7Tg50i11LqQETxLyemexHRslQEo2oXItQkH5DRcyX
YieAjZazrQ+GsCIWfYWot7rbrWh9ajb4X5WxgxtUwik4xxLhh6pMF7MskkVvmuJvjP55ddfRDYFP
85aH4zL+eV6gsJ3u6yxtyNMe8R+EnEioEFz1Ci8VCulCZVLZj5j4dlf4qszEpNylY2FXGCFVfM7B
rrjgEChA3z8uV83baZAYRspxnzfu3RZf2/ktbh9tGrdzz923V9IzvQ8idMlUYowCfcGeyLH1LbYE
LfUwb7e2IsbHXh/Nd1BmzlqD+3mPLfL6hCAn3x2v9GGL+EX25Fh6IlRflR/dbehLBRVUTmVgLGcb
5UKSNQxp9kPEh0GR0FFm4R++hISOV5ULPjP86nNFZMeGd87El+AUc1MwQ3tSWUv5ttpFk+1pegc9
U3ELeVNWzCccnDg8Sjsl0I/eoSnV9ZuJ2esE1BrPC9LytHj4joZXw2jfmKInHJNM9BG1yPPuwY3E
voU70oo5jw2JsGDuiDUbOfh8sjGCEqGa/RuUybQOZvriAU0sHk9OZ6R1lPcx8xm5VjRKDbodRD23
50Z3obcVldhjeUwz3bY5i7K5iiKZIfI7ULGPVgxU//3gmDigkFvVUc5JoCyrKziS5FH93BT3gFyP
YXXw7ILqi3g2C4tqFrrXbuAF6QDqtCCoPbAlHDfwqYn7sQWA0zYW8k1EEoBUKCsdc0fg0uHqO6J0
lvMY6pTGW/sdpPsfQWYFupqvrVMvrEqHthDR1CwYgN8zPd1KC/i4NKzUPsSO9uCyiZWmHG/4PVnW
vBpmd9TLKrnFa7ZrWRdsG0i9SrSaRfzSW3gunpF/FkEnqRbdexyGdRBX/qD8IJTHluQDwuT32/eL
bXqEjz7pSByya+mh2BoRwam+o6CYAc8PrxROxHdaRrNOhuFkRe5w7lD5VDu9Vtom1eD6ZMpL2lfy
aqb0syjW/5C/J67CMuJzu8jPhJ1YVPELnxvB/l6iaC4etrBYAWe1utoFr3+oXsM2CRurmJO1g9gp
Sf8jC/gHvWRWOUyBwnXSEt2pb/VRfTkvqsLtx90ReXBOSuwXinmVS0ACj2FrTJl4+7xfvwCOl4Sx
Ejmxi3Nd2LuuvQlJVJO6A/fV+40r+5HYjflkOaZlS85CAl2eTd3kuWtKOLHJdMTe8GuxOJexJm3R
uy8/H0x2/qqcWnIlGIJ/WabRvN7Z8ayKPpHir1Zw6c+g7duDsO/dJJTqFrj+K1SPsaFttrhdjhrA
gSsq9o2dwpocRu3tbgjXAGl+7J2xdFNlXpxd5JV8MGJkHZzXXm68uclD+uA8dTjbo8QwCBVFOzeC
0w0Le/HHvUBbpQE0V14gjlM0LKCqxxgmsDzXCqJpkODtsHudQ1390GrNj//Shki6uLDx7m4h+Iyk
2svdJHiaW2vCmc1l3kvQ7M7f/6bBHKkgETVSCmO7CBWdndvPG0CkxNG74jOIw8H/9SwB2MavXTVs
oopoCmWe/CA1fp3LIp/dJZoTbJqiEi4f84/0tmWSuXr3dtwl/tissUFESk8EEuPdg/g0jSY8sZEQ
zY2uiw+gYyXYC2n1nGtoWwjDVgtBEwfMnRDwXjSJ+RkOL7rCjDVMGPmTrMSELEOeLEUy8I8eXs3G
L4RmdAzJjJnu2omdudCAd7YkF6unr+Zew5FSG3GRd89DlYxW0k4plnJNUWRPHmAndJbDuOr75BJI
ZQSln33F6nKBB5gMLFzaEekzY9mzLizIfaqb97WpNlcewg73KVUqKHHsWRuDpBViIMADgRlTajST
1LXfOr1NLexiz2ZLmsspDa4m7Utfk2zpVfF2ZOyt0v0ua9MVVlIInpHa+3elgAEWh4lf0A7upXKh
wEvzsdf8MYHZjDl9MqFXceS3xblTvx3KFVvolk4AXblyNIFne5hg6JXztyjAxF8ok0ReyF8qvNrD
UQ1KfCtZTRznH8Kr/FiHbe5AgEd+oD+zxpF9yuYm59LlWAE4dKluHfoyJF7ZXqvs4wecPBaGoSO7
KSArPLTlgt5A3Lm+2L798sP9M4rGETsHQb+xdNYf11JPfwCBGA1ZP0Zj4cIeGVyV4S0iwEkeGsZr
CwqnQeCu/f2eJWELZ41zFMqJr5o38m9wad3QYDbHS0xaHoF01abV4G2FCLaPv/3GnP7h+pBc3065
OB9UpPxSldEHA0JKwUXzqmt0BhSur+uS7kMPTezef62/H+/yhRatRlnM2VnUWwoXMKR/6WYOP98B
HBZyTHuBGsVSecBh3BRDj90RazoRv6GWRvGtbGKMPZNfcAK3hlyo+Kdp14vWVJ5hi0Y9W+91wpy9
v/VLHBGNwSyIcpqvKf0qdYgMLV9Xv0uXBOEVp2bHC9voYPv7L0Agl9Sd5nZbQTJUU5u560ceKu5C
v3aLPdF8+KupTLF0S3cz7hs56OIX4AXm71mc3dub5hciDRjMIYp6G6ozoN1xGDiN1iBVqqGus04S
YWi67n8E7B4S8MLwf056YyhzkrmDO8q/YWB+8orOjc+YRSu8p9yYfbZppSRT7D87vUpCkHfVGdQk
QfgtLPCYSBO7yGN6qy7uzBZd5Vb/vv48eVEugVxHpXYxN8hsaYG86k3Si/fOxrL6VzVq/9qSfIgW
H00DeiABtenx3YYkl63LUTJhqvLdKgR7yfVx9ti3hqAfua+Yxg91jLaNdHfWgYu5UEtnUoAxaWoC
1rjhIUnjcQZBn7WtQzYu/Q4p43LLRu1FVPEDXTJJoGN8jqgh6Pjm8/HmNJ0VS6Dd8K/jSEdbQlii
AzyM0u0PIheQFD7nUvgYNw8oauZiCQ5shnbtlnlqVViyXXcOG0lIW70u76ZiPiq5vc3rlpWqikcM
ZpuQsbK249KH0SCFxrri/n1ZXADNCYgBDUUcIN/G/99ebIeCCDa/YLXMLiJGKaYrwe/gdeeZRDHb
yUhVTjHkrN8Y2BYxBnZ5roLdxcR8RB4LhoRojhPj3FonbwQvdcYxDvctTpXoRS43BSeYW66c6kat
SO4VHGj0vmL5C27Dgz5syBgPJd+PEcOoglKkWUMNx1zhXD9lbhC/B4HNi2IVU7dSHYH5f/zrESKG
WzvB4ewmEVxbe1tcWYbdiqHeQaeJGP8whIW4Ld/y2Gndy5O/C7Bagnj0d1Vbqwohhb4LUWfNndDh
p7/b3l2IFR5PNsddflPUXwdx9/+836RGmBfBtTmApXE4gw3EsMeLXouVCtqh2P9DiSFwV92IYb7P
umFkJiOtDRerWCJ+cVfz1LsB2ZE9oCf6bMhKUkoN9uCnEkXei9mhHQZrWT18WzcgATosV8TlUj1G
RazZ4gXlBLMfOL+9z5KJ+hqqU34OEjW2TANYwMEDmb8rkHcH2PmvRJpJ/gWDspil3IhcaiKvZii2
6paG16t6dXyLkUPjGbXlERIlUFMR3PMSgHCZ/vR9KLRcovl8iMlHaboG/RrirXn7r6+V6sKoNtmJ
S04WlUR630zXPeoZy7rqnI3QIih8/oxcgBEKFG3SMaL+wGJHmRvSn+q4b8idPsqV7oh49/G+Zo8H
cm5G4uZcAZqPI+vtEEkftz1ZThZKsz1WqcnOeBqcP95gLbhBPAVyXxJ8LY16FCGti/2OnYgq/udw
JajrO1SEw0jLT5ScwtxvL9CBwssY7YeXW4nBwfw5LEcGEzkFk36BRNkr6Wk6x0ysinJAinIixN1k
7U/akeOFukk6ngBdn6rPwc3iHHXtlX9CYkBDynQquYe807Q7vaGjcSKTpuj/sexYoWNY3R0XHk0X
caOsZ8fCHwIYOs+RSnKaay6xy11lC1d4cMQSjfonMXkW71JlFKAUZtCybC9U+FMS0aiO4uHbrQJn
VDGP2TnS/q8FDIlV/CainbunZu+c4YWOGgba1PUgY5QSlef8XulH1bAUbP27CTjJn38MwPoUXQ+D
E9tqOB1UVe9oi7BkX04+7e2ReaPXbfMAz22IbPqp2rydhQIGLE2FB8iOd4dOej3PjbuUNyIfMTpZ
PfLtRoPjhmmQGn+sAaDuLhQ3eEJx5UcT1fPn0mw8Ox3TXBrNCrvdw7KSnCj5zXvxuHdywxu/POWZ
0ARC54fpAzxb6ubytMUsTtceqWTVy18e/Ez1BmX6BLVY/79QyRGbfJpazJ4J0DjurEcA9fpAjVyF
bbdD97yLfLZpbflqZrHLDtxV/R3/u6VHXgW26vUh90eu+PVNpOzGrq0vMMJsBsJ08bdFwFbgpt+I
t7OUGnIuxQZ/Mu4EXyDaybV2r54UChBPHQttRkXj3PyP2+6GnaLbPGHwHH+5zdHg2TuPTukhPV5c
2nSW64vGj+wMImXjdI4IWbn0O40Md8iophTO8X4XBSOSIuT+si1ywoHO3vypl85XFQC3LTDClDsA
HTikQD5sYG+dYLMF4NJ2Z7PpG0aPWKRyYssNP1RkNOtW/LbdoLLPpF4f+YPCBiiMhXT5BF0FILC9
uul8RvHnbO2xnetTJh5W8BXnY0uj3RTyykSHs5T7adbc4r968eUTzS4DIWJ9mA9McDO6e7yz3Ypv
Gs490x75tAUeCOD4rrHgOQNQO9/WmPMc8cysNcyRN2eXkUoC4Tuf564FJvAovjSQ3ROgZCahFu1z
oVfnNRpr3lOtJoZ0qX1EZvdMdywzNtBYsTPVSg/7jfzo6Bvkj8+rS7hlwVYU887UtyFQuXERHBeU
oefIdzq8PxHQvzXT5jQOsIK3Y60V9XpDER4EO7inkrwdPn7sLPaVJ8YTYy0ZerSAY+12wIe342JC
9vj1+VDnGnVj1LL3oJ2fk8dFCG3WSNBNVREA4JLkD/PjRFvQAQ0/wjdnxmtPCCscaf6++yQwCRwO
eibWL2k4drAfghiExDyK3v/PlR8s+17GVanNWZO+a2H60pnMWGQaMP5yVCcqYoOdNd+vPp7TU3pE
YIu4OxLCwWY5yhtslaz5j/Cc+sZAAhs5AWFajK2t60nju6L+diE3yLl1UgjbAFhGPMT8OLKKfGBT
dUBqWgepQ8Wu1D0aSRmuFTUqWbmdJOYSSPppjdbJe4Va48x010oqA2aK4e/PPwI6sVuCcv05OwXH
Q81Wa6hnOwS4Px/yZgvUUzDsitlJsqTXmmXi2gshhPpN8rrAQi9UvUcuFViIUCPBjpCyqzNVy7vl
+5LfiSHF2omtxGSmYDPRRDuUQ2cObtPKdy8maaRTi701xAk8R+tT0vk6sBD5D+FxBxaQWSSiTAgt
X20D/eZmgvQc1wYM+WgNHsoUnJw0BxJL3nqi/sIR7QOIj2zQ9GLdeP4D2VoGFFMe45vbcNA67k7F
rxZvo9eemleNuSu/WrPbVnWlWn2i6O59Y0QW2eiq7oGsbQCWd0t3cSwsuuBYNnV38sf8OISqW/ye
HUdgm17kUwRibA3Ea5qtrrloPsyfPtVBSXZ2aiLr9PkQMvPkTE1rDksb8GuSIe5yLY0HOtGp9SZV
1W63U1ui6orWaS0BnCn6Eu/XtTwELuEoiIRPszDLRiW3nP3x4n693CUjbHyQthWKhwvT1mdsH3WB
5I3gfUoklCZPUWjHT69eEJMZDMm+C5ULlHe2sNbQ8tp2RZ2zuOQJeR1N2mqp+8a++KRx0OjkpHh1
D5/11k3IqcKRk5pif/LCmGbOg/P6wNZeXSnXNMG3/P7zyLcrOKLDDHyGBXsbFNAZ99n86zr3XjIb
u3AuQxewRatjnFyIm/qUcQQ29Q9jTzzuLL7lPVHTbJ1bhmcaAn3JOCy0NeihHOUFVlGAtU+PbeXb
xh4pLtUddyv7BwzG0MY/XCc1+XUTFMFabuyWAQ1M52Zlhhdf11YfCaqGIgzmJ3SnjbcUqtlsQ+rM
p7RlAJpt85jJMT4KptBxOdittRZ3s/zfmIvdPwhIhm1Owd5gsQg0CpotrEBnaLN4ybcqp9M4lkKi
kcwbF+pM3sRMoEhKKr75FGIbz3lvjRYF8gYYniBKE325uyw58vrKj91G7lJGxzVTHFXL3u+N7AlF
0IxjFfSEKKJHpKqvPnZKI5kpA0qSqy+AWbKn49YhXAOseAROxQxS18xwRKbQfdYA0QH7tenG29Q1
hGnmjB8R/hD49ogiSPrqZhIvvffGP/vz7/G+GXKYIIG2/DSByXFQiAp3OB0WPMlVnQjUcDaK2K7O
FRxw5+75Fg4SEwB38TpfCDi1JxYG4c7al7naEtV4RZ008GR9JaLCzvuPmlpemoVh3gYb6jrgaprL
TbaDpf23RAryq+r7PPYRVnw8IeTsTam30PwkQwbphAJsUMjiT54GU1mSG/Q0MltdJUj6w5Dfh+VE
ctXFuGhX0kwLDmHoSznf0F1QPN2i4WZkFVw4zOOvP78AtaSMwb8Qn0bdu8kHxf3Tw6VJSjnB4XIK
dluDLXtjxlVOp5aqTncG2F0/1VcmqCkD7r2VmXB5gzhL2ATbyXjYpsSN6SXeiqnsWoMa3lUn1sj6
4FzCPhYc4iMT2tk5DaEhI/ihGl5pcqHotSkkzh87dx5jy3FX750iW0TjjTMOk/efFBpMlnKucQY7
HSVQ75rIZHvlvyITS79OhxGYyvmYO5lAmkfzx0aEatI0CB8W/+f9Jmyn76tL16XI65yGDZCXP7mO
rffKvgD+XhEggRVmhceIAswkUEn0dmKsDkUrOGtKa9Stw81IUqT1dQooOH2oCMN0jQmsaN/lmj4M
9zO6Q/w8MAsm3UWMbPcgvOJqi21mCtRDNaU7D/R2kYPs0OMItTSvpCe9WZV31qSE9m2UyTmskUc8
cLf8X3EfuMQGgLyePg+8wPehqIzXzkhToSquKOBJACugZSsVx69wNn/5F5cnry0lX0E/BB1qbRKg
3PPTll+7ce9VMhedvqq8APJTKiyxaB1Ji+V+HrTYbHWIMVlBupJMYMkVE41Ug6s7noZV9xcx1a9t
G222zGKwex47uqlU6yB3OeHvFNi3jzA1QFUGDmdPybmxO/s85JVUOFafcBoSPQq82dDJFQJnCHIm
BfYkLheNYEuhS4sprB1Wb4Bi/KtVJ6qiHWeGx43tdNYlsQIh0ndhsli8qmrXnL7yHtLLqKbHgPsp
E4MF+KjYh8kFyOydpoztY0d9ovb/RFJimhOsGAnPEZMESWTLDGsTA8U03AZhoa4rrZ7oh7E5WEwb
bKL9qTiCDkrqaoBZnyctfN98l2u2PUw1e13AS7w0E30BtyC5ZVuFZesSfKtgDYSDq6mns4t5FljV
z81AIULOYeCSq32nANV561LEGG3jHIc/ayke0swUz9cuTlt0zu3Bi19CFX/OD3cPEngXlSwOa2V3
UoKpn9VYw5grygEGjDIUelMndv5N0y462YecEqAROo/Ngq0a4vQyweuktxVwcXiXbDUxdTPyn/aA
7vvFF2MDPJwGuFA4ALR45nKp8ig/e4cwfjJeYKaB7n43AZ9xQCnhSg5D0ch7CwVu+C4ESVyv1cGy
v9b7RRe3ZTl3xOC3fhIwlFqapmlA4lPr5UlZxQx4k9nc3w0LIgS/gQNus/VyAauzjjpYpCJxV8NT
4zd0m4rGdzJlBTtYqLi1ErK4fAmJThntvLjZPPLCJSqyXiIp8eTxqMf3nbU0ulMiESCVc4sIpowS
DJRstmJ87BcT2Gi/QknIJIt3OC0lASyxhSxR7VJnl9cb2jJnTyaiIGcG77PN5OQ9OjgZ1TLg1zTg
1JPHZ0pMHzbA+GVX6k3ui49ugDewmhSODIq2+d+jdaCoP861nZEa2rEHmL/16U4Hm2UtLgaUOiZy
oipkQPSTWuH9EVCGCSbNvgb0ul8D1+5+SwPdfGcrSG9G8kI+mDyZoRxcRaaoy7QRAj/VhVM1n1yA
61DIPifFvCauZCEB9fav/AiQ58EUCOXi8Bi1t7BdDGGq1uVyVT5VNGRjL3aCFAK6g9s2hm7h/QXE
U3p3qMc0IcHSYUx10qPPDf9FY1MDuj2eM8GddDEjX0JthQiJ1XgE1yaFPjbVyYC/3U7TkVKXREjJ
1skVZF3WFHJIOaYM+hc5EL05lDZoHggD/jGhm0vMVRYMI72PdDibqEaPH+A1TYqKL27U2H5B2Tdc
I8YvMrTV1s+xrxgXyqevnsZIlF4a/rdB6h/IbWLYnRPrOYEticSUMTu0dutNhfoDNlTQImmp+bZZ
Mx53y2acoJcYs/MzP2bzxhzQhtswhxUMha2barpQV+Y+9ig8NZxSN252yy8/I6N2DtDGhQmYnt8Z
XMD8jiERa3M9z2L2rVSxV1ghxsJvWfSj812EVhaat0uv66d2VRtsTKiWCIDkwhB/fB59FyJO24SQ
jNU9h4jERyoig9CcfkD7gW1rxzCDbmUwcxJucvfORKL7jg9CXhmYaVfBkiE6HaoQaOgOtaku5bQ+
1zyBmZnzTczb+Lz65eJSGAh/etw3HbKWfAdtVjuqtlILbgaMyK7qQNJYlCS3bmBjZ5X21YYV1fM7
sovqammzxAwPGXsWOA0qWc5irrB/FVLj5F7Yb2vZubsGv7+Bi2nnmuXPhdr+Z21VOiMxe/kwJ9K0
2ghrSgaBjwo5qFufNLNZ592jdWKlWPpXrLSNN3zLRtVsNuTEiKaI/nyTfTs08FLv4aF/9bMeym3h
qceO4CLWg6/FTBHKmtev6YnpVvwqzl0OtQdiycJ72WFBflWobFCv88cqyLQ5z2EkfmtQIHP1yvuG
SbnD5IZMB15YMCZgho1FaM4POcSsAEDmGPjy30XPZK5NnZo7Wl9iEJzquz+SUmaHr6lqSbA+AMXI
rdB5PBrdEoLtQppJa4eHCnNIXt1uQE2Ia0QtQDQQUDGlbji2sz8p7yeLdBnV4lNce7hYhxB+cZmp
hel5nwxQyjV793PTKGZZQzt28QDAbQSE0x3NMZjatIu7+gmH0u+XV9IFDGHQXn1pMMqoMovg68Af
g1oZtqgZIC3punM3TfnSPFxZgTYzdtFPayYmKIVCoKyNe1QaYr0jnx9h/SlA5KgCGc6c4BW0wj2s
H36Egc1/c3cZwMrYhZxY2JD93azSF1tWwYRovM+sY8nYlqoOev2UOpRFb3UHy/yaH6/dRIlIrgqk
o9oUbx05VuY2o1FwyraIp/+Q54T/dhsXOS/UxvHKHnjQfktGhgwiHZOFqEY0huz1IckHqODXXcqA
vWs5h/LOWvXE2yYekaKu52Sf0W/V80HMek/57+2B9RlwufWQlEGEGfe38jIRZeg64XkvzTFR7jyH
bN7bZPRLrWFP6FjGju3pvRmgkIu91vpA5ghsoSEmecZ6I7u2hswJNSm/7Y5QBy3dfgDG/FTfas0x
8mwL/xEIrACG4nhiPfgKvk71KOCitS2bOTI1KUXUvK19tJY0l/ggOEP3uOOtPqZidzGVnq2fYSj9
rXkFgptMRz5Tq991bekFgGJJIGhFMUcD9FCKRNEToYfNKvMqgPbpLqY+yMP3nlMyfBhNwyZXIkqZ
cdmH5V8d9eY0B1AYEuyLzf+QlbUh4KzL89+AVcWh/mgbjP6XfXAz6QyI2Gh5lMCd4gRwpiyQH5dB
aokg3TC/3fdsNpTshvP2mRfJw4rmnjWVYO9cHWBnKi11oMfPhUtL/0HVwefCRPscuZyixPjJz2og
qNi6Ijp4Lp5mc3OAumfJfowwaJ5oYhokZvAYKeEDqWmaCTBEh0R8DXSpCn4iwuewCLeFISjxjquF
0yP0LM676xcwYRJmwUqSgGhVGyVk9UDeJBK9MGXWNca1pLOL3l8PWrvBM4L8plMO+INkcKbTSxEn
EL96KxMtBgV+61pOvaYWnrf2l7xf7/s991qv71LeKtPPOobPTdPJmVWbtdY/jJz33A1GVSBpF8Fx
TIlyez5Q8SvEG7joRyzCBewWDybV7cYR/o6luy4Na7H1ZlpBHGMjjgEKC1nsiaTt96AGad60faxH
2ng1uA5rXa/5BD1zN6NPRSdkDGyVc947jKVFHL6pfYL5cienDeCABrtw2tn3Zo35TNb9gPxG6cDf
jb0TM8r0L9notHrYOTzbQ96VULoofzBGL9dFHnGTLHBWF7ztJ3NUNmzjD5GlgAwFU6vVy/iHRhOz
l5XNiyQL+EwYoTcNXWRHJIMYfbsZkAssgNKvRr9EqqdxtlUPmltB9vyWA7xhQHWqnXaUzw+jHs6q
ijM9ZzjNgUHexCXlhv9IBtNMZU8fNthQMxOTvMcAMMvpSYVzm8Lvsb1f6XS+TkjW/uWnVRMPqZ8Y
mBs5gcLaroteov8vPnzg4WzIpenoHrmfq37Qjpv3Q02e6h8E5kbwzMDoKLecYOPl2oaxJvR2uCvV
SMmeKvcaCFSyRZ3GyBPFKZQ0RGHfVc0XPF/AjotBmMg9UlmfNNfarVMfWlwaCa6EOTuUqaSqQCRP
ftvgyVEM8aNBLYP5pcS4hUb3jL+a6J6fNzUtSuGqKzfIpQcwqgJum+A3pTYZEycRpH5HV696rO9y
Pd1VLt0eO4TrKEoKoRPEHpXi3LT/hQYQ38PjJ7464c02lrS6l2iyGucSbAyXM5lzsP+EFcYHynlM
qg868j3BnJRF9BRoxxOcU2vqWTlXJ41La1fZvyoxOiDnu8KlUtMmtJ9XA2tbNwhJoOHO17SjOzhH
4tL0TkB/KwvAyJ/dHHQW+3Ns0Pf9S2fzmAO7NZggFE9LnMA63JftQx8ViD6iv7xZs6oCmpHuUwCv
Su9kAx46yRj6PvVGu9mzwKofdyEMXweWJLLVcuKy7oZPwpFQtOGEDqTMyT+qiaMaZHLtyoA7dZuP
AoQYtgc2WHjOIuL8gRguy9bWX7gmuXvnwer+vKndSU+Qv+1kHDfvvCALjBpnomCv0OfVEEXlAe8i
c9ZUd0aAJ0KFn78BN6Dds2WpfBs0HDpbNaHjAouwaYsHtb7P2Obbby6jkPga+gJPBRTbTl7/9FY7
5CJkdHXiO4rxhtmFmlWEvL7t67gy2Lar3DmHMpip1/7ALiTz9BIxY2vOUBKNack8MY1FSS3WMihM
xB/Nn0hHtyUm0h9TFngqnW8q4Mqsaz5ebhlcFUS9ZMZu9zqBoXN7mAmXN5b+HH2TYlxNccIDwpxw
OCP3f7pvHpt7Qm4JGgy0KMSUnXUsr5Z9whNm+QhQOrciIDubIOK94iUdQ2H5Oz3D4yD8JPeJ/UHX
DTWIL6po8vpl5hpgkHAIt8qOyi5cjy+7A8EIUhz0sHDyyZHpD7AEe/vhFeB1QU5pSGWEYHk1Q1Zd
m4fYztj72sxXdlfRfy+sFaxNSkkJqUXeHocIaFbfomH7AMkvuAV214ZHg5E6bPzY8aSAyFtAH1bk
+JFY/ZcNAdE+3PPRTG71zufi8pifFBgSL8Ibht6tDLCLK4LKiIUZQjE3uiDfjI4HCa2ejvzKSZ5j
+Y8ThHkFOVY057/hkrhhGjfRaEOlYvBvX71+x0F6FWvAchw7PASzsSgCReal3EVqxSYI6ssxVABh
+dEtBvAYNWY5R+Up5JDQEdV6106pSHhxWSpA5U/B70dT0FW5QmrXY7XH9VWu3JxYoHkGNm1kPpHz
0yiXvEmcMaft5Ma2niIlg5PLZ4J0D7F0AWW32ipRQ2+/HIMAYsUBmdW/XxVplIeyoIRIe7owiXjy
XtjHW6Z7KRE6xPjfIChh+1vuo1TCCAP9r1bBZ8Wdq4uYzufjzTIN/mMAhQbeoSfwEzq7WGZSxPoo
w/udsSBVloMjZJwyxkbedktTITcPLxynEC5nyCQ14Lz7eFsQVsmS5MvMaIqaIIRuA754ggScIA5C
0/vAYtY9fuy9ZJfA2c/YmFndjyGEXtyyNToAwB+DXgPyl8+Y+kd/hV/4mzAtyX9rHldLsz5eQQXf
6lgIuK1B9cMIMsz78RcnYJuYhQvEFq68Nwom7lO9amiYNUwf0siANg5YWOTXqK+INdLqT6BP/VBm
6G7Eb/1eBsllLOcANz8JHkhe6U8Z+L8D6THaoyFB8twKzBkma8c21acUA9kKU2fVB35SFuZPXhzV
cnyOhkgWfd7QGbiqEOjmj1rSz6GU426UrL2uthZUCy8wn9r3XBBKM4iuc+ulyonglNpXkuDxpx2m
XtCcHtkmMwvdQd1dYKPlTIyI7sD2gyl0/NjI+vgLAou/2Vtj4g+iRpte8YsVsp2m5l8IfPbiOx6t
FQ3J9uGMEtlV8Zhwe/VAq0PDuH3tc6/1+m8MWwRVH339/KRDdzZEe8OQTHaRZX721gJJUO8S/BHo
IK7gRuZyKJs0bJIbGa+ob0zc/PnUbget+KJ/yllwUWJF+0yt8MK0N+9lP3WFlTnOa2lUA12u05yI
k8oM8dnFQOYJ0dNF7BqETiwNaX7XnwWSf6MKpZ3FR8I9FwfNBMOo+z+sFZVd3vAADelJpekqN1Dk
HUaycoFBMkksdrLCE8AttVSQwYBbcWijg/mPLua6HjXE/OGE5b6XB4C3wSlH1+0LZ/Om/juPw641
MV7Nhr57zvH3HHMUfVI8c4/urnb5R4YW65HYD5DFYzBmBSO12Yz/7QrnL4eK1zP9mEAfooIpd1DV
bGz/EoL6IBgwg6/OkjYbxjmWh3EBYq4NEbdhL9q0FLHRX3PKUp2WiagUn2T44xGtkEovPbdgE6s3
NAK9oPKcN9jIpLP3kZkvbBpBLYZdSi4mn1PTZjppTjHpQsGhgHMAzCZATbILedDuztgDKIXvyv+F
l5Z9MR7YihzhmSrxK9B1b4EmFp+c4tAmXRBtwaZm261jBPCfbbI+nryFh1AkiV/tND5ZG/gs0F5L
rTMXt3yjdx5lTF29Qkz060BBsrLebZQ7IvGbAzA+dqJT84+rckKxE/b7au9jmjeeh+Ctsx2UPqrq
C04JzWVU6NjlS1Eeka38PZd89hD3oIKVOZOcxAhNWBqnH218MrmlJhyfL61TCrbnfZ09KgReUTV/
uf08IDvUP2+2BiHz4Iy6kL5CC8+L1PBqdJf957gZZsdR75sMW84U5y/VFChR87JujcYe07Vpqf+N
plfzzNVVJJwFJ6XxkNApbmA3rA0pw+FRdPIzD/YPpNlZqJDI6cAFFaTvC55MW4RFUKIjE/stKAIT
W12PTS2V8W8Z5JOR901mmDVoH/w4IAr26QbcupMT4f+MeoZUKxKYA2100eGucergeI37mX3fWQAa
FooKgnnc4BpO8pFbcpu/8yEhIWQIRepS89TtEj09hes2PXwlIJq8yzYV2eO0ULHBrtXDLZQhIQJl
3k8npUwai7TIgsx0qVo2WEtD1hUltkZoBf+pnui8b6km3t+A3WfPe/Bk9Q2U8yu5fk/hUoXBsRgD
MeHnYEv2fpuR56NUrbMsFP7PzcrX1qEvEyV5Cyfjod9hW/qgdaI1dfoPmPImnyRQDOUZgTO/x28k
V5wgFkVq7+jw8d29Y9qX2HhWeeswG2JfXe3QIfDrl/cmasUvsWIWbUUomWjYJN5SvFjYV9OJbbyB
U6sCu/+iJzsHcXriqoGadda8gPsj1LAma5+bWr/iGXWZQ7Oy9Fu/tfLlGscoc7H/Su+mTNMq/Gt6
a8chY2jSB5WsJDTndzIr4FVODisF7k6yCwT5ska0Qw6qdW8abOKuna8+q9iMNHfb8QjWeSpiPhHw
QGYmWOpoiGP4ic9VXsoSQtskP07LWIdiZWO9P7jQztGMMlRLfj6RZJsLK3rHVxcLchqVOb9XtLos
BkRWLA+/OqILG63pGyZEHVjxlNL3UbeO4gWIu5qsveyj8xsz3K7wz1VUNtH3PM5mz8CgrPn4gYTc
f0GdPyfZuPkX8N+1UlJ8JtczQ8osdRwEWz+6qwFRSiHK1eeFnWWBeuA7tDQCZ4PsrqgqvPAa19Y6
Mu/foLox4b5nhaNRm/PNX7v5xLl5K/kp8uumuc+wTT+nJmSwohFJOMVU5maQwVyKq2kz+zE3Xiqj
h0jihDfmqnK/cJ4SgRvq0+mtdIUpSnPK7MB96Hsnzs/2BbbBJFliDJAkezVsQ3oaEhhOIf6VWQr9
a1JbUyf/8TgYICtYYDWgLKaMl5lZl58cYXiF8h3P+Nzq2SPpnA2SU9iUt7oPydDUHDX9EnHYb/Bc
3GyfTr38Bzp5d2Icy8EcLo7l0Tl4bpzUyH6FFMgk/mTMyouHs2cyML12JeZjoEMpAOcLB3I61CqJ
GMHccwq4ekmdqM2Im66tG7joQ59FfxYMEAaVjw67Xcd2N6BIwodkma6rOQof3wUeNuiVBSH8yuov
foo0vxlM/GiE8PoBB4bEJaSLfPfukM1LTGfWUJOuyCSXEyqNjsKnz+mdVkjuk0BJNGXq9aS8pLaJ
4GWvupG1bxTHI7y9e51GNeuMmd9ILfZb0uEaNQL2Bk8dG1/Wb1aBSvHUnT83Vzn959LNIygFp2DO
qySpxhw1L+0AOoQ7qmPstiUIdP+mBxGC+R8g8oceoc+ZbOvpVzlvLApdR7RJvd3WtjRdVWZMCr7x
6bTuV24pozMbzaQ7rsoE0oJTuEj+p31BWfGJfqhbG+73hfsftbeZCjF5jSMK+49Wju2i6N7YZ/96
cMhJOlUJWwCL9Zrf2S2olCFlr3t57cO0xtF/S+W2p0m+7VZQKLhCBIcNJPKRUYQgmrFTf5F/BLLy
J/Gu/stCvXqKErYfbUE+CezDXzmRPc+KfCQg7cQ14q17b6N+mVtC4U450WPwtDBLf+90usEkEKcZ
vEdsbBGu9xXFD+R/ep92+Ges3wI92S5Ss8PXgYQ8j1zkkWJLdmefeMX1TGpfwD/ZbfcPaRr3ejhq
JsqDE4fxYNmDPoN/w/5akHuj4O705VSOASM6o2OqcJfsmfcfU9vZ+pEOJQsYpTwWQEQEcEeqDQUW
+3Msfyv50fJZAdPNtxS4FOO2v0Uj2yeSPY79/CSC8aoOs5887W7krWfEI3vm5eMhRPkXN2kdh17M
EhT5hUm71O2fCxpTAyPvhI4CuX3l9n4KPwVtsLl1zi1GwOUWWpvFMlfroB2GsmZ3gg2aO+zYXoJm
bMzfywjgznQcbSxbc6mYIMjxzbiBXUrOejcdSWQI9zhUknoTlzN+F/VI0J2DUfNN0jPvnbHNGw4x
ALbMoN/AZUVK2kvpBm78MphaYY0bkp44iAeyfk7Q6sorCuNHVd6pZbQRL4rq1OYYmE00b0NWu1yq
bUUks5L9+FQ9H85IvlHP1KtUwTHogk7jZr921yvueNNg7VGyL0Q8wgZq/u5jV1y5i6BdEuTXo0xs
noY2VWwPUzvmchK8j5XYTiqDgG+ynNFmll98oB6qZzRGAX2+8iRmdvrQgZQVIWKgN0iQHvERZt/b
fJ2yKy5ww41L8TkFpFjAL7TkgYILGD/RLythBIxVKbOutE3r+qDHw4Xb6OqBtnHlwc+1L/jMw1h8
UbHSvjLB1OYvgn41eZUQELAldfPO9AuXKvnsawkk8OKRR2OJD9XM3rdPtFZ46w/OzShGg5FQtQlZ
RyvFaZxRueOAqS/d1sf0VUBu7b27VnfmTQsLnwpZOVwPK7pfa9QuzaBCcdZXo4bkt4uhFpvlg/O2
4WyLLsGzpI6cG4JCulLn8eo4vn+VIIWEKt6F6DN9VHzeXOTwwcPeo/szykqY2Nk0X6xocQBY9dgS
uW6dRgMW6p4u1xrstBejv8W1nzAc6GT+S/8qit25bgdGC6NPd+aN2nNZw7ckTO/sl3huVrxh16W2
ZirWNrdTihaNuh/KKdHOphGK0F9K7o31TrZHwMiHUyXuV7nAcIEcPotDpI3Gfxcqegx1YNVORu0M
YrRD9kPvvwm48qWUwzavsvQlKoZA74VaUSuDYweBsXuqzhGM7UG0T9LqhGiHzjqT7khQS1YK+WW5
595HgETgnL5eoy3IMdlY/KNdRuO9+w0IUihfxQmo7hLYhzs5f3iJG3aaSTeAVqZ8Hl3tA3qQrpMW
t0lpKkAcmAfuGVuyZXTygh+hMnY7Xs85WAnnE7RO5kOVHEOHZ3WR2SaaCvqGJ6jYsmGZP0vR97l3
b+Ad2kwaTfcLSU6ks9cAMFAhJBUVl/zRrtuD2F2cq52lz6gbc4ShJ4Zb3/R67n4REFzgtYLCaBD/
tg5zkijmlmfgrXhfhZrRAlCxSChQoV33W1cN41jEG6Xy3sI0B6cRDlUEyEIrm5fqlW2kRDemxbx8
bAUasJqp6yPcfP6D54HrhZJg//+C+Hy3DMJBzYsgpEFLuyU86bPP/Z9ojwcTg+cpybwewLKVTdJQ
LKf0+diWSTC8zwYgn7RtPcf0ocq6wcTXIRpi+mIDuc36E4KjUttmNdToMzza8aHA443VTNGlgjDr
D1Hrd5mnacKliTguF2MgBzJppBE5rdEJJoaU8fDdyIOAOl14KcVYqcKSpAtMqo2q/yWTnCxiWDiM
locbwfT5F7MonG5DRnoaqipO1XjnWgP6AkcWSRQeizMaFTE4S8khAvBJkwXRpmpk6N6x2Dbe6VoW
8gfp7YzXyVoVS4yFe64tYYGxvB2Lcd06phsA+1fdpzzD2uD7ZZkXXaEQnYhvUzEgjFPLNoYqFlmu
V9ePkqoBHrzYdo4Zy97X4yqK6ggAA9FpEb9+Ouo7wCMxnXCCjhGPdxGSwGf4ipy7jLepmzdeV4SV
3nsmoRz/F+S3uaeKx/KvUo6d90LCvWmD5m1iGMI3NQs/XjIY/8pu3hc8+JvA6Krxwt5fchsaFv/C
1AO86ojPCR5prt26e3IoXnhGPnG2yFkCwqvWuJGy3zk2i4+85pcTHMZbzC2C/+28oZATg9Qqj2fA
t2pbuuoExz88Fjlh9pSihBdv/vXi6n1nrprNm+0Fpd9tC5w/RL68fojyrBpC3L6vdYzMBPxV6QEs
xFLB5hto2RGE4rfnDXwZuBu/LqOt22daCa8NGV/7+AkwUdkjlmanv9dCgHBZkA+yVUTUukp9M/NS
A150Zfl42iV1A1AvErzsxyxva6/6mk+dETbpNf5RfnhPI+B+fz4qVqQg6vhWwgq7PvwZSDe5IwB2
7HaxkboQpLhY0rswvyDo4Tn9q71CC/bdyKvs9hF60u850CiYLDZMLDUFS1YXLPzAStEib0737xUZ
WP2TLqgQES/m+QWcwoOQETAIEUXLp/HSZDv4r016MgCJXnLR1Usb1Gz84xuvqPlBoebkeaXsVhYV
mpLiBB36TywoNHS9io3REotdhrEHCp5Z6TczFXZ/buK9pIyWQBY5yruNYoVJcZbEhstgwFQpIoTq
52XVpNXh8SncNZ/DLvUrufcqbeW/L1TLyHxwO4wni7MEArr4Pxs6Ca89QcP/iQJPL1CbaowWyTUO
ijZX+P5pUXV3PzjI9uUXZzpWXFuECmXxn70YAgR3suP0uT8FuQ+sdViXJfU46JEWlieUKU1MCSWf
X9jMv9vEUTk/vjwHUG5ifpy7sMl2S/Qv46WPl9uRBZaJovxJraBoebkdxAqbrbZ1W2QBPLwDWSjy
FH8KrO7R/U4f94Hug+gCNOXIV3U67iodE9k8kXRIv0IZ6/0UAGaD0+kG7bo++4zMtn8oumTljr3a
lodmwrrkYFRf57uB/WQuCzae0wOOTqgqGDPZhDL1Y+1bQ8cQYRi0G+OrluTCn932OAo/UlBjlXu0
03IyPGz2OzzakVOVkQmnBXV4qDimlUGLpLMV2x7vyNzeh/D6cAkbJoeGTTy2HwvvLuL9YmPTISRU
HZA6cVS/0nkygJuyh1iDpoijS6HX4ujU/gxTzeYbcyIBptGHXvMkM0neMIyfPUWJefONjqcONeJJ
iFm5PCuilycu8UF7+PzzY1Xj6jtnzjRLu0eEV2EUEpm9v10I0swA7t4Tk6u6wSUWEH9eJO9zVWNR
ejMjwEixhREJMZ3G0jV5sEANB1NB69inD9t1mHg1sDFMFuwwQuyPO3YtVnicu5GHYxcfbM244UtX
O5oEO/ZlnoL01PG21Mqy1vYQdgb0RLO7k1dP9dLfoPMG3xiF6WcEvkQgxIX4M9/AGlLvY9mkT8/0
LpHWJAhrsb8hxhUUxACn1k3WVfPES2xDmAm0qJon10iq+6vaGZGuwRMXrVXM1Q/5FMRmtdedwlSM
RuQLlUA8SIMqmtriGkdwUh1xENfXLOu7sM+Ay+WtVa3TxHDJOK3jPfiW9li184VXYGiPwwZreNMq
kgrdrSFlcSELNJpkd0MhRO3lH90wJYDVZhywmBvdH0+5IiOvpmobtMIaEQ3xDgt8olCQ3yBr0cQm
M2NkG3vDJrk0DnVmktoKE8ROzVGOY0hNp3HhoQAZ9Z2Td0JyDXCC0bUwBXOFBIx5QLyV9sYbMMGy
Y2d42RVzUvnLnaSLv13/9x8JzOJ5RitKy7Dc+YZixSXlcVUGs/lKNNtuBqZEB9VDj/fLMTwAUl19
8LzVQ71+T4Rw0awZhaKPvLDbvxhDwhCQuO9G+aNC2H2WD1O+UyHyzGfNsV6gRkZQcM72mAGTAslq
6DiX+0FqgRSlaZggSNJCzgMlV4delpwZBgXy08UQuSBFusO7syRiZaAC2H4gmap8iO10YkpjkIt2
X19hsC3mB761/i4846JDWot5KlRt7bVXRlBEhMr/ZvIYThmWFdsH00kpBc/7zoCq724CDQON8XmG
dsJ1OlI2lrgRyCCQaeztbLCxtPMSH8XTHmuKIVnVg48bfF1LXuXl5WPl9P1MU3nRTcol86d7jIMN
nvnrPw3Z9s22xSNfp/YScq6CsnQDVipwKOiQRPyUk+v0mE1xLvG+0pRC8UZDnxCfgZuj6q2dVEni
xONdqpGnKGJF6rIedNU8eC2t8LBNaBC0gBJaFVKWDa5Q5ISxU9K7Y4kByYuE7TC6wNlKgy893Prv
bW3pezfOoui2sJ96/bjSM8nxCz3iICZY0Tedv/IEvA4fiPV3TFfl7xiH8vQoHO3b7DgKtf04BbOH
dFOmMV0ag4Y8meyUzjAsIdA48OFak4Qp6cbbtaJYv3rZ8H6JJoEbBxYLbvIFLURsXWeFILvD1PDL
92OvZyEFJTU9rc32Ru1M58x2N/LZLwkhUa9/kc2gKJc78pYiv+rxOVz06NCR47yYvv5Mn2O8Kic5
/WYtCpSqbZZoT6r1nro7eUcHtlP+TLcActx8sQABkn77HU2gMTDjWg1r5CZvPKWHMeCmLxyQ6/IH
jeDkRtQ8aR3DHd6xvFJyXHRI8Osl0rJdzSpqC8xGTAcRXzi3C604G4rK/B/TzFUhAJUcMDWuz0j5
oUMKBjq+BXHoBm7fEIkhqPTNZXQPQp2laR3gIfvs0OJj2/OlH771zDhrX85WpJhO2gAU1AxxTbVn
/MfRTp3JM9B0uyfQSifpb0DZXQrPwcVYZngv0MNgYEaMbtPoni3wf30ZKR0q4RgT6zXB6T/TCI+n
nllGD8xwafQpSx3rnJP8y7K403uD6fNBPmTBINqT4sR9ojgxIbXe55YRnjHznrVwPbedi+EEZGVD
EUEOcHSd3HXhB/ufhC64K5qo7t7gmNe77vHOe428w4DS7MDzRYcOLN6kWfD1Qk0BxRaLAIY7MKeC
PkXYr31h/R+GZvRlFpoJSao0EkPu8JL0nUDhNk8Q3nP6RSOUDaaTHYjp1q4oqrv3BMgEAf2GCVeB
IkMFlktDnIJjy+ESBL7zttWfpKyR+fIZMhlY1w2Oo8rZszeis2HZvH0upUArhgdUefEm1n3pmvbi
mVL58HPPVMGyEVH8JehRpNsMCvaibRwQSAvOh7n7X/XUq0QwonSXrMTaUR3YM0NR/aUw1gkC0CVv
dFv4GJTPtiUjXquoCbre+Irlm9qnV2eOYKwm9+iQnsks+1vJnqdQKSey95ubx11SQS+abb+34zYy
s2mdfdbciPBUOP5ErCCCPJROwb8BpAQ4VLoJNFRHvmzaTxG+ntYvQwY9Gs/bUdLHZdHbxNb54Ok9
glSlpqSFsNd5hnTuxBjgNLkH7JHumIoI91UZu3B3jShAuPbGVZIvPArmXTdJxZEi3hrbUSk8P2X7
zt2uIApdvCI91zGb60c4UHAhgVipFUH2rxEXs/iVZWaMsdba/EOz+ENQ1pR29JBq6765vYz0Ec6+
K3dpVDsi39vFVlD3Qs/1OzG6VslvkjwvXJQqrQv/pNTuBb3LLULbD4VObhD1PPTnzOARDK6BsYqU
8bFpn92tFsnjZ9MNxr2NubzL8hwjy26/t37gs3trZ/UwugTjTPPvqV7sour6wLfWc4XilzcB9RxX
1f2dcqMq1SFO11uFMM6SWpwEap09k+mjNRQgl2v4F3cuhNnAKuvF+ALLkh48wyN6VFdBLHpDdgHz
TY1IhJLdFTcYWPrrVYVKoT4qUjRRBTQQM03jpCZqWAmSe+mod6hRJfSzwbqZGy1NFp+z5NDzWpRY
z6DpaAqSW29Uco10bYAWZQ1X1t2leURnTRtJsximIyu86IxvJUvsxhbsGHAiXsnzpHc9h7xks8An
Aut2popxomYqM0dPemhMk647r1HOlOGwflFb776q6uK7q1mhf3h6WRDyrZOqDwHmzuzmyJLNbyaA
3IJsvkb0AB1/MtwiaAy/outokNjssRb/sbtGgEzhC8nQ3rZA3j1+0mpMWyro+uOO6EzIo9CjZQAM
chUMZ4DyFzeOm8dnJYxWOFNL+bH+qqkL94dsS8HMmFI2Fg+I6Ceus7WO6C21CVK5DJSONLFY76lI
biBhiU9906b5mHXdRr0p1HLP2EqrG9ENy5JjYPPEoGkdOn33vtW4Q8+KGlLhiZy2Cros+aVxv1o7
GY3W9KZRPD78JBr4GC3aS7fmNYWfVDopxeer818c2JN+17wQ6kTACMZ8TH+DHgszYk6cBg1M+Urh
FThueccxm0eqcM8g0yPjw+mprE01KVCgXQqc6M3UMzPW3konW1irsfOrH8HgK69SSJFCYmTb/i7o
NPLqoUClbHCj/5fMeaWRSJz6jVJSXkwgGIuNaRqnG+edEkRlPPbENrq3Gnj5ZrB9di3xLCK6YW7K
Sns9X5jWycNGW55VcW/BtAr5KJGFL861cKpY7i33+IEIsTl10+ZrhLfT/vy64cV50qKdbwHBdGks
qVM3jIVObOdG5cDY5P164VxanKe26vIS6TQDwFVc2X/Kr6pMaEveL6YboJBYn//Pk+uYMHp/WhHr
TNJC4VXBpdzCHlE91B+Az/nVjlgazGFTP5NZOzGsfwNIFORNGqjpKv6MapH2UNHgjVgAVv1MvxiK
XXR3QRyfQCkihwRX1s5EMr0AZbozQSbLITWp4/gc/6DZMGhNqRdRdGNxq5kXgqLW+nEPI2ou4Z7f
G/VyWt3faiVkoV5CvxvQ+h/Kh9yzdG1GkCwapVv3ibKzzDCTLwCGiWYsbsgwv9AhaalYJ38xA+F0
jgS2sT6IhVBX9OHFC+pgFAzdb2wWspA3+rjybByV2r+R1YszQIPfmfAtYd4sbsyj0j/gF1bngnng
k5LT43mlzeflOTVhEs0lH5vaQ2lKTU9PhxMCwmRQWkM6Nw9qbGmF4OLAKwRDCDycfwdbKC67SVYk
lwmBsJI7+/uz1c+mv5ysyLvehqZ6oHPqHwJMk+OfPIugMKRjj1bLR28jH48dvMeNIWm/2+gIq/OU
3oK6drkbRAOS86BBla0xz+OKbFOagSAs6AYjLa9nwpjFL8SQil18+VygTgPshHS3gatN4PkbYvN1
Jrppczj295LMNZTMvqoQg5b9+jSzRs6SUECc8bTtt5qXyJf2AjE3Zjdwfrth7InCjPTFiv6118/0
Z+gcAEuSIokiqC8DgPUwtTn4mKvCP6je5+AfMtuzjMOmZ9t8SJNzkZNzWuk8XjTO090zPoCJ/Vjj
7/zdhYw4oz97kxYB86hJzGtOUwWa5FfU16c8XGBJBhl/9+W2l4lpJaZOtR7M4/HD779zh7lcIas1
CxOtOJmP8Xz5HnQbk1D/m+S2vGWrCSLbbi4KUomFehm495xM8ifB7kfh40qekqj0d4xUio8GITPi
OKGXR/YTjYaE9O+FEo8pe4Vve96GWLrXTYCawx4RVHxfX6mpCw3Of414F0cSV73hhxOZXBME/a4Z
5LWQO0VRKO9lu73t7r16EFwjboOJDtB4BmpEVUho4eUQ5loN7Tzqi3423SDVbuw3s+QSBbyYxeyH
Enog1HbqZsd7KT0mcBfuUdhTqeeYvCgC5+SaGYPwJelsDsz65Pg8TFad73LJRBdCg5aEe9Bh5gV4
g3iiZR1pHk+ZUhStF7Vwmg3BizMeGN0BLv/JEJe3NaafC7uSjRNT0zO4Wk20fwDtRT/dQOAdyQE3
J3tA4mQvsskSrxyDeR7oP1dYOBM4ukGNl+a+GvXjaohBEy4O1qc/+KA0j3YNeCijRDu/siIBOD+A
+F+VdBAypD39V8KtmLKtOqU4BeH80DHqSEd0ee7Di++tATr6ay3ovRGNn/5W3eLfHXFW8t08bZrU
EuJrnzZxXMU9QxLP58DSbnmQsVvbEflgo74vwAinDWV33WV6Q7216q1Nia6lvBHZufd1lZu+BUbU
ORdPubzy0QBosy2qb1Cxfn0JGNozUKLQw5IJrDsDGo1kAYXyX402wnMTO2gq8L1idqk4F7tD374z
D9a9EXWkMdBkg+EseJp8SQZM1ZH/KSML5QJRVpXYuvH+ZH3Gl/BbOUETk8kPkFM1s76WRuiA0X8t
B/O7wh9/o3Ls4PqEM9HyTDRW2LNz9BxO/7lsrZzwF8rIzM7R8RWsBO4PO+7Ha4j+LymCfc02ZTJ9
Qp5AL7wPstXQ4EKPcTrxNaL30wjiG+LzT513yOtBDfZUXg5llXwYYLsd+a0rZqYUdebBgnnWZFW+
wh9hNU5hlYQaq5QaBKvJKzJjUkN65EuD8uFtLdqRVBXdJe+aAUjEnza4LWJ08EwKjNGq8KKTHTmP
kpRvK4bdatnHJ9iAl30kFJMY++76LYZ/EXowDPb8a33KxISEOKT9u2hEDhj6rFciNFkZ013ZELAN
USBT9V6+ixHSP4fsP+LIRawzueV8Cfj/E9gXjBC5zWG3EFiQ0/cJBfFpTg/52tpSuIFK6c5j3tLu
OxV726d/ObPKhuM6al8Yx/xDSjIGG8bgqD66KhAFOAd6k+QSYmStgekr6Zwj11m3676nAjJAgnWi
vO+Qdi3nrNBEMjB23CSzcRK6mZNTLXAul4j6hpXRdGdflNUnYy256Hky9HKMjhGH2R7rryZcjKrl
+uZTdhQ7uu1MPHRdU+zrV6qpjcwPWeuVfFiAoko4x1zX6TYQ/JBS3AEFIdfgHfJcgxy8HYlzgNLe
bFhYXB2N0e4g9H85yPTKXIoy/gzg2Z290YR18ZoPF6+cO2+X84z9Pvl878EQWhJNVLqGRIw8kcoL
x8EtJlPtyDKeB3AEsWRWZHvffdKIDsmlYGU37tXdBvCDbx7JxndKunXb9o3BHUcEiyxszW7+HKG1
ps7qFwGFY/lk+egn1Tr3WfpCoSpKbe3+yyKXh34LPBom5IZAiS8VS/3O5mJvrTiikFydTSPTIY/x
J+qiZC2Pm9zDXmM731qj8g0jfMfvwnnGSfcyaUbkm3Qzq5SVKUejHbR8nL1FA07tM7dz8aeJLeRS
au5xF9ag171mPkXzW+wR8CLwT3AMMztyYW1ZdsF+Kevz02HMrgR0g67k291HDS9TZDwjv7JPrU7J
mJeMYp7qNIR3+af+18Qv1zxsKiscVx/rEIb7ZlymkAsTNG6QTrGNQBZW7nqU5KtotfFL1QGE6KH5
b5rCoqrb5Nw/C5hDBzJt/lxspEgOMzv+T+zegIlW/MoqoFsi+pzltrH38q4EDFLpMFkppqSedrTw
MFRQw6HXOP/MOc3bBsrLjsCnNskMCgM8gZ6Wh63CNV8pSy+5AY5vopneJSeyZFdCivITzsbPN4UK
Od2wUCuGiN4X+U9dkbcwlY1FW/NglIS+TuD14DxTbDrfMHitfKB/0Np4FAoVPyFjrrrE93hBYfOx
RT24IR3R/szB8Ycp+riJVTuKV33b1KnI/StkQxxWnT5wUyUWoFB2Gqps9E40iJG0txUb1Pyi9JMa
9H+2JhI1eoSdABoTkMuqs5R7/1BACwFfHSEImPGpPNRnCcLM2zYYAVSTAGSDbbSV/goxpQNxt9pw
rCzDmAlLU0Xik9pJp1ZcK3dXIFh7qnkOfqHBHGXVkKY3Qa2HO9LCcp1x1USL6Y123a/5F2sPOUTY
7zTbpH2YZCmmK2rCBOAYm7pqu20GW703i0vrM5BCKl5Trq2WU58m0+WfbRis9XxS3SWSI8mqGcRX
mr7PASj96aHCk6jEK1Eaci0tjL85MbyzvyXYwKN7jSCFJ6g6cunrGb50t+2SIQ7DWsrF9cpIS8fL
GzP3+1LEflMjo+HNj6scfM9JCLy/QeGVD3Nkf3iq8G7NswwgTh7KA/sBz2eReUtiaANDqEsJlggM
8sjF7/4caXVRjoNx7ZHh85ajdUMhveBVCzo2z23nK6wGqwIuK9adYjHk4LaSfSJkM3VUD9p95PYk
9jhr7GpKbIrNibrs1cETVQve5FkRZ7UvqEBFxjYA2Sv8Am+OoqwsWq/SNuh8JY6C737Fcj4C4v4I
ve0OdmWdBW9jrOv4wBmPf7/H/cxQBGl+Eua+6xc1s8QN1bIR/ooZB/XJbR+mXrnRJygfaZad96ka
QUgPXnJcMrbPPhMQeD6IXLXclARpbfrhLf5Yk9S/dMVlaCX9yVjZ6lkCaymvy+bZqDMNrCnPUp5O
ncyYNG4AFIXMhtui4mV5uII4vPKFc8QkUOy6Kld7v1dEl1rTRuDPYZQkNWwTrvttvcS74h6pyHpn
gei6YpylAsxGdbZcu0ZuUv4kCjiO0vqa0Wcv1tOs0TPoLSrsjl6++IcfoIls8YpRcgS6Ddu1SXUS
leXFXxSDSOoB5mdvEsAvNg8rgAiL9HwwwmFidC0qc9EYGv3iZOXkkvfW7I43Aro1EVZE9M0k1C6r
nMk7GE3yT0uOINohjqp/+hcOczr7NrWA7JeRvQoB8BEUKXK6lPMZLhRkCZC10ytndzoFngD2P4Pj
Hal58JFSTy+fX20CRF93F6f3a1p+N14dI77O+R5dfblplq5BFt5uly26ZNswyA+eWS8GYs9hEcRi
YxIqhDveBcS7pnctApX7Q+AVryrLOQKv3IcBK7GWyTvRMtUyyId/vKXzh1hf4e/1VGOISyQcvj4D
0EOd73BwsoovS7iaT2O3crqfb/s4+j4htGRE5kp/9KYxuYtBAIq1HdRtRPGceib1IhfvLnUi9MOk
4bc+ELdopSdCt22gr8PG7vjmcPtoOWg6APUxg9eBEYo1KZAUuOOZMRVVJ2BcvmHN274H4rVAUCey
UrAeAkzIRGPI9/kcWaTx7pMObV2s9Lp8iuVxBW72dcf0p6Dps4c+FAu0jl3Z2/izLEPjXK8CC2JO
eCzerQXVyYKxYgBDcnqzWfhBtIDuA363GTQS4HdXbp9TmJ7cCI/+i+uPl1owZRdkSjjXbKLyKZNP
cZrN11kd5jte+9lRYNpT8S3lt2eCQAJiKzg+7Vl+FEZ17DkYcjKWxDwHJNfpE0PKbTyOcDkjd2iw
M/HIaq6JzUvHL4c+KQDgM2x2cDtimSJS/KyKmfsD3La3B1QftUhyxg/EQCXrcdw9nbrIb1JGb2Px
j/B/Sp76Sakagzq/8wqWBbuWpTHdmzrKMAooJcK5bi8bJhl6+dVi5KRmsn/Ot8t48KgDEw5j5CwQ
ZXYEGtaZYPEwlMywcVTjnzKIw+50SdNZIZUnTJBQvCqZxKuYsyCIG/UMzjj41TUae4BpCUT1AZrF
CyGRGUCOPPp9VtryMxYB8owa3jOIzvkmbwrnGaLU65sd8lrXTj0QENnONgInOEhZmWkxnPinFYhJ
prXmCApFOLdXcC2YbaB8JhiUBs14ST650YNGCOowZPYJrPp+yL7YXv1wpGz9lB8fGSVaf8DOTnWI
W0xuqYeWU+DmoUGikgXdJlz+wNi9pwMJWSnjXBKnQC/EdVgC5xOF4gsr6wvDRjlyKYpFqZdWoVC6
MFXQDaLzzLlsyiOyjIEMy5sfEGx4D1KmL+o2VhKmHKyk+8a4+6HShousQ9peCk2xQuEjNJZqWFdt
DbYGviYU67hpZHaJ76CRc377IXdPLmpTAzaZCG7KHCLnWP9d6Vt9VxVveMOgghRJ8Y6WkGFDba1i
7iBOQY+lx4tPJh9Ja6f3vyLRiryW5rltX3b9jY3f6+HjWt5Ir8gCZAtW/IfjoOy+hrcUASFfIGG9
u6OQFYtYD/dh3BU0w7WG81CUn1WjqEoOoSGNsNnTwAZUY4w7ALz7CvGyKVHOGe1WZ+pGHdi1oS1O
5mqKM36X2on/epUHyPiGWuj6FmpYa0mGDD7ooGfer7v5O3EcruIznb+NR9ldXcgVzEdOOT2PJI7W
vjZQWsBolv3Bi7t9Rbhna7my51DhXfwQAct0WVxCiuOAdiFxgMr96ixOmMkyELZgYYiT3NdyNnz6
8rb+YvA8u4rydw1WctnN2WuGPVTNdrh9ZRFFChbcXIW+c0ZUTyqHz8Jz6LxWSWKs2fDun9suqduD
/Ugjj+s8L0fAvuVeU0YK8oqAj3s0H0+ncs7SM4StIyiJQDuvXYUc6RzEQNegZ4NKyCBTkWrY9rev
A8tKsWi+dOtVg2pg2UPfwIO/NwrRMtYFR5co2xizQmQoRPI2H3YPLm10P5RzFpq2lo2WEqg/0AKi
9Pzov8pZ0kZujX7o3UCFzbm1s+JvXcBMP48w/PVRU9APII33zL3XlNMb7Z25+OwX6QBjFQztr2h2
Q9LvVrfpn40SZSsPs4XF3W3pYgj/hE8sDS8g3DxvRQI1VYpsc4W7eWGx6HbTS9mC1qb/ZX58xRvc
w8L4gsxVGD56c2rtMX/5RJegheYtp+wLtheILJBj6OiZJgHjVGPyX5VegceE7sjbFLpGbk071Dlt
G+GhQOXmksfPdiDJu764Ge8wjkY/W65zTszIAm5oRi8Ydrcmlvhwn+z/masOF1nqLRDOMotTrINq
CO2wt6kCev/KmmZqE0h2Qn9g5aMh1wp8+aXA7FCSw0VlxczIRtT58+2HR6Wk5IT6yvHPGg9gIk7O
5GSc+QW/07Q2H+4vKnagfs4dLcJKuNGqNsCybVOOoCzKrus4zHdtK/IJGi3YMlk5wzK2nYgOwDrQ
jwi+kEoGw4IGwnBy9Yp3XY0yariPcbibyCySrDQPRqW1I/j3Y0MyRYD4gqgdSayLejnJVeEePw/y
sfeXV0CTAo6AJzW6r2MGLBw5ulGLGdd+RVmye7JKa6ZVPdnhKmmuxQmMv2Q66R/LZUpN9Is4kQ9S
aqIFHJBwko6tSMeRM/Q3wZxQVHmvZqrRir/i7pBvmhZCDHvyYCV76cjHrUdGOus7dUHdKMR6BZ2f
xCTahnT/DSMJh8HAMoXSA54dkR8PCTi3i8I9gsHorka6B/7S8bR7BJnqgRV47bXZqGxvp2kCGaCZ
kTGpM/CMKzR9tkZnhuZmyeyzMD3UPnPwFU9LiuI9SgbCVFG8YKUIiyEjAVYAZ02ZD1JLCNnPF3W/
N4vj7IIqihqkwucP3pC/YyA20eCZved2dkBfeP2+Emkzk3K7Q2GMbY/zZRPpLGRwuJcvZtA1Bz/A
9MsUlR68oRCy4LZzkFyf8VMIl6p7t+f/CxBOl2m3c5SiWwfMfYkbJsGXINor5O7+//vlJo71NX0F
L3tFn2jGr1qrXnIK+1QtKlv8qkgZe3TAnv05W3c/wKVbZ9jwwasSBLVBz2oDhVR4VLXw1Q4EwrxJ
pLs5UdTJ1s6tDt23CgbkF1PPX7b5BUXpQG53/4PKzyzdiDd0sZiNuFSUSdIE08G6HmziyvOqCKuW
sRE4NB77rn+zeoUtJ56Jz7vBgTxp5jfdoVoDkCjmw4TgOG3nMeJHqA6cMp4pNdP/59/irFCg8sHx
J0/RRnLP00/I+N24AnKSfNFVqAsSjm9Xc1lYMnyCHDfNL6HB8CHOP5eaDiQLvWh5r9W6vRrqUUCW
loXf9zmM1Xj80qVsoypUlVF3xM+WsY8kGeIudZZLiFGeveZ7yKfAX2tvDozZNx/8fFn0SJKkEthW
fDv+lels+46SLwCX1DeqBOENXIVpttlnNrARnOqB1WafNEELmP+GpuE02YXMJU9CdtOKIogOeW2v
CZ8XUNEx5KPzUY8LnuucsK+1FfmnK73hFx60aMLOYCMwdXi8jG6GCCYL2q4HgmovEh1XAxauUTfA
KfmxQN/1XgZmNlI+XRF9XIA1qprS+JZMYgdV/GhybDni54II3xQkIBmYnfMK/W+Lm4Nr2z+pYqfa
/ZrK7Pdlu4AnHVWrlM555Ao8ZdNc0QSBhEGmO4A8MtqLpFp+IKkthPQ8zOQoMhA4WBFoBIR66gJ6
o+XOP9LQE2LoCLFqgrlVgWm2TD9kXBigEjqQXYWixVI5Mcu/n7j6HMDsobL4W8hV/eJvoMwXkFAP
xbFqw4BiME+675EQS8YV8Cc468SuxZZawzz4hXjcWKJVclTHbOEPSp5ADqPBzhXngiNLRCBxb5j/
IvWokdd4X1vzfQVeqU0Jdjv45KzS/m5ZS8Tx1BHR3jRnY3mfln5Azxq57nu7+bZM7jc92u9whx5l
kbGICkOLhXGV7BmoIeOUQMjfdTjm5ykGscKtp6yPiN7/ROFhYaYkrZa8wriWnzQq/MiOrn4DC3sC
P9VZQAWT8ERdr0vV/N3hmpENnh8naTPZCCqdyRR9z+ra3S2HvLCEKgZeFtRTstr+nHn4/axqq0oa
ZtznP3j35jo6H1/C9kAYdlK3yCXdVREgZI6E+YsKf1xlgvZWRPX74lKoO1pCn4R8FE3HDYEm5P+7
Nf4nwWAjk+meXT3Wl+vB9SEG/tFkEmePYx3UuTvp2vIqj6EFphr3LUsCTZdBvpwGDakmGborIFl6
Cas1Fbwe3f3hMZqw/OHP2ksjc6Rx947dauOc9HZTRWy+XVJ70wuZm5pD1GUHI1nt/uUvk8VgUaHI
RWh58M73NTYGC6oCNQphJaEe2RLBEWVTZVy0ZNGM7yEuDmOq4ymFJsvxQN7CFHbqSE0V5y59+Kl+
o9W67wvXVjPN3ML9c0fQIv3QqItfpRBPBifuoORQkOhdEQ4EBxFCYVKyfC/6GpkwM742hO44jPH+
Ycw3CVgbPi3Ig17TwE/VTvjSU4lRtX6uZX8/Kpoxt2wORBYuR22Wbw6/t33bXfRT+TYOcshHjrAI
KNp6Eu36zNKXqwWmeI4dTc4QldY/BnNr0XtJIiNcF83PS+owaENJqQvR9CiM8YXrl/NuPgu7ut2y
mGomHclNWx1rYVZ4tvc+DOhn2KxCSdFzCcefJ7FRyWdEWKqYbvIK8lkM1+gcW8JHeCaq5tVSr3VG
E2Yveqj3tEXA3XO4MyB3aj1W8H0wv8RSkvyV9enSJ9nqTGUS+z4O4BrSjNwazB2R0+gAQOFt06r9
KSAN/bG1l82/iUpf8rUTH9ljQTYH8T6YJD8ka2BWVX973IINARMlZKFWcAlPWR0lItFrrd3wSY9W
oYMBBABcRkfza6KDzgYkF/xKhmW2OqEe9pQ9wm7NKJi3KMxs6gAazIcqb4SiC0yHXjULCBG0q0eN
BGxRrVz/lgavwQoMlNmZwIdZ6jnlmkI48GdDbb4qMFDDefWzcNj5kvoPtgStkuGYgoNOawtLeBdC
cy18+IxuSkRgPoC6JxLZcCoUZROVSz57/OOnnkwO/vjBYLas2602mpLHFNbzIGw6rSeefoA4uahc
iwS2sh15PJoJK+qdBT/39kSpm+0n6dH3lzzmbGE2YAcsvOj4hnEE0IkfU8I+S8DZ+bjAFb2jhDuo
ymZF4UAXxZXupvYvaurCHJn8oJJZjjKbFbop4w4tCj8s9Fg9deJkT8Xb5ghJZU9ueNXRD49r1sKy
wHxhzpP71iPwDFA/o69AbmewdvbBBLBmiaRcqURM2FVKhhe5Uc9e7Yo9Ac2Gkp2uGnimT3AZma1t
B2XmRDE47Zy18k+lgDRTUYT5YcVf0xScgDAuSDO29k/N2tGSBFYATEYSfvLGXVqk3dxVuTZ9axv/
tfnQNJk1RCabzoO0/HIq3DwTZmh+fEuqGmVTPB6Wdnyoe0ihdt6sNICIzndhYS9d352VSlJEiVvr
GV6Z+XEOOTwI385kTkYhYlLJpJT0op1UMJeWBCcuV1ZHqy4JC2jXFRo3JfF6O1edsf7ZG8awG7b+
r4P78KSu58JYa0MqRZNlieQG31Qn6WZh+6JTwGUM54ZaxuAnK7HotH3ONqY+wQEc1lioG1uZJ/1L
j5lVFNCP6Z27vqWBcvRqdIVK2IEN7gkmtnjiJs1imkrsH4/lBIaHUfjLC1NPCLbn3Tdnl2ciIsso
XHRRtDF7maKPfSWu2KFazJc3a1hbUr8Zu2P0Ne9vySKQDzEh3B/1r6FsBWf0Ac2Lo2u2FhlO8EjJ
MqSkks6wwURi0ROxLpr+UIDcGwvui8qjeTRqaxOWd2207v0uoqJYrWpOc3+6I3kCfEW293bQICOf
ao+QM7qnD7wjCxVO/NMrr6tz8kOh8y5dS5awUBeq7NO0FekO3aEb21wW/8RAvKj35g2oZaHfe4uD
KXyQz4KSN2lU2N1GMAsj7RVgGRojw+6wwJCvPdR1thKpoBuChXmbZIpbe6gSE/T4AlcCWKeVMKIE
1SGi5D8UNnKSYz8uVYKof4mNUln9P+YqKUbDTr265VCasc72JBKwSAHdXvoO0PgVdmwXeI6FqcVo
ORhqRkxxylRdNnF1m/1wU83NyHWTin7ncv2iAyTfIRGg6POeU3hV5iNORxIBkHnSyXuKgwpsPza+
/Ka12b8LSXd0XlRzORqrO4FL/JWzgTAjpoSJXWM428Dc4k7UbjZk1nalW0gGlgN3YIx4afUum/qk
25s3E1Tz+4+y6GidtSA25h/1NHrmC95G/nxQER2Fm9JN/m9GvxUHtBJtBMiucEriZwk741AJBFPb
bWKHsBMlKQeuy2P4bcJSYNuMngWUYmOpLfTarI0n+PSiP+PHemavD0jVxKuwj6gdSFCWEDBXn9/+
QSSgZL4c8QcTtlacZWiFa+ZSutnu26hkVb+dHXVnAhq+AOp/zLFS5UVLFjpN/4CPTN5N89FrcO06
bFV3lRr23CwjhSbIgwvIoCwTwwytaClPIPXQLt8W2kXM7kBc7d0XPDeZEWhiYB8BxrdHYXIxnPnx
XmiBNzbj1xh4qpNMOHYsyjjta4Er7iu9k0V8eOzLE7aR3dzjX9vLDTfc8oweza+0zdvackQdhKFl
k4cPvYtgGyxW7ce7RvJySz7x0ZVhYrqJ0Qehsp1LJaGOcHCJ4nIZQ/QrY8UXHl9O7LkkdrNZsRbA
zWsT3JqBapHOjDmkzMTjLodTQ+H5c99ht5gqwzkYb+IdSDMGU4KVPIaokbzauSoC8WI4oKJUgA3h
r6BjxlNl9DL8EXM9XUyoL+o2X5Ou22MidoapLY6Tp1v5XDIYKarEF9Wjb/bc11plR3Ixp8N4pQlf
V0tzrpzj4FDzWq7TTXNUYC9qRAXROX8fJwmnl9S6i2WNInqvIQRMTjtSKwGlLxaZ/2DdCM0kRD3y
QxRurI3ASaERCRuamlDlsKfz++jFweodfPQ7NdYsFQSgxa6b8pF1gy8Kb/6IWu8i5EAxlxyWhuBs
U+BPC/BtnUOS3AR9TORTaK0Ikg9Icp3MFa5ioRKWwnbEGc6NctpGdwjMSKrwToR8QLfOKpFoie7Z
nubBypQBnIjY+2aufi0UJyfBFseJ9PVi2pzaVeBovcgVDb/d8r8payz9yGSiPN7EfuiRLc4E0kXX
qNLJbOGuRvx4VVaW666DBBarmpGPXeHaZ8ohT/afDI+LxJi/mHyGVW/kP/YrMfeTFLfjYRxxFgfJ
XO+TwvBwYPKzSZ7Lgr9iOnC82cshCChi3uTFaezCzxnA+92/2ckXttWEr1UEy5sdG71DVZdO3cdr
65CTCHdAqMJgy9V3aBDSMGpJPQ52CDgXUJ2NTf9K9ITWtlVQ0pAy1nqzwmSzcWH0p9IiTASNyb++
vH9OrW2zBvIETrZb45b9lCTve92140ye/Vo7zx3sLOyTeiihyrqCqyYI/HsASucC2kS6tyREP272
0lT1fxKl8DKff258JyHPTRjsjIXTG3hIUUzvqZq2hLeOf0uYeyGpQ5VxQGqDb13r2EL5en1IhUaB
OK/rDE2NcoimMaWAVva39aq12osvyC442YVaTRYK+B30dWNbASJbO+kMgLKd+cx8GNuBLUqsrXdp
nZlLF0b2Qo5fIqZUaMbTVCx14mI9jrDIMMZ7/v2A7pk+0ksP3t2tE1s083FmtLJEF4kAeXqzu8Zr
0Pe5aFaOOuR3/oXwk2KcHSGprXz8lgfvu2d1GPo7dlPP48y8xWlpOI3peL9IzIGpIaBFdMFjICkw
6fHD9/KRDp7ukgF0/ryMjF4Av9v0zSCPXD8YnK0wKi8rp387oljP4np7keNT42Zn8wbIZFGJ8K6G
RepYpR4Zb2g63HWGVGgHhLpKVsnwkH3AcTh7CC/xdwcmiVxRsdbAf2zA3rdu09KlEHT7z2BHAhvt
oHpl0qdMLyOf9QXg1HNQgh9oheBm/O5epzIUCPPiUJJiPi8X7Des/pgv2EXIo395m+tmj+1wQfz9
/8Lt3wFvjbK22VJwRudOsiw0DqwZ+OV6cvGK1cIAq+myxeSYJTY3IlYqMxA2q/XjnCXXeKpflka2
UmG046VCoFksBweO6tIFaJsunOzlKoW8LVt8T/O5Z1D+Czx/QzfCzi499UGF+E6aF/zGN6WeoHG6
C/xJ3i0T4UA6zAK7CnK21CQeQgKeRqDD0Y1D2C4ZEvEXyKY5RnWeGldv2QS7KxPSQ5PxjaPe1fik
EBjiBYAilM32xXJcYhgrl4Uaz+lMOhcdL5587+bKSHVf9HZntzS3P/TKQS1x0GZ7s3CYIcF32gHO
1NnqEE29X10VSvvMge9I5YnpGnzmtnYQ1RA2jlUQDRpCUs1uLKbr09h6/2rqaQZEUQmIEcX7YFDY
0J2kAQ+jqV0UrDiL/xvpwRjc18y+Phb+PBC2IMSvK73gFJx/IzT96FawApRJCMwDOTVsFyiMerV0
WCH13F76jmHImD26rlI5Fm4mletKaKAsIAuiCxfU6v3CotORmWX7qnBoHz/HG0lGr9xVLogAraAC
edZ1OeW/MmrxQEh65du/Vt10QEEicgmTBm2lU3SssD9KE+tLl4DI+qQS4Os9oQThpBFEczI2D3S0
urlrgmZ+b1bqH05z4XIKRyHzYxsQiCmCB7+fbSteiYPZFmP+h0hopz3EBAsSowcKjn1nwyEH34dX
YJjvWzafAxiGN0fErxrAxNVocROGh4+F80NiOFfRBLLeQKvO4Wd3YSs1xkDJcLgvwTqN+I8ICU6+
h0IYjOZnYpmVHtD+WPzKFkJvnyRhXuU9S/nYL/S7Ev7oShZkr9y8IR6RCYqW4SA5GpPQqmgRMo1Y
oc/CUExWjUqNkWpqcWEwhivHb1nG/C7Ukj1OR9eg8STguFDY88MnG/wQ2bYCANqw9YdHT+BNJGqi
bsQQCKhibCn7wsWG4uukJQsB50e0XcfQv50rE3p7IdvEfATvnbo9Trq56XnzlnmQ79ZoHq5RSRgA
4jCrDydgRf7mTN7A3tBjLPiEcmT/VKmNn+fNyiMViVplXkWhRs0hQ1LTP/ItQL7Xr5phDE0oqGoD
bWLncdQ8tGhQDHuMux643QxMfnwND9pixjhvJfvDr4Z0Uf0BxGFoOF/iNO8R7iwVBYA3nTsjM97H
Oh1nMm7R7pG2sQEZeTiD/HcOCnVrQvxy6JnWjeeqKP7HwNTkr0nu3HG8Snq9+HwJkprfHEqivAJU
Mbta6WADovkqEo0X+LnHgIDv5cM0JP+d2R0WNAOvg7lDHZess+TwQJjmVRggrWExeVOtJb3sZuzu
KCatsOEynXpBq3M186Fo+oAkB5MCaYYCqimpbHgjJKJrrewgG+titNOugc03T4S/g3oeEsbXN2aX
0dZCVzOJrfTtMQ823ejAzmABB0NFRJudMMqH32hB+V30zyG41WHIahwcLVdyWd/pIo23/5WaW3uE
rK1YkL/02sJmdLjOFWqzJ1HoHKVtmV5fajfF0SB1Qmu07K1o20+FsBPFxfeDxUpa9/nGp2N6f9aA
3UmcmvZcGg7+H50QYd/0B2n3Cmi+kgUKzsrNTV3ZcCEWlwxD0ELVNoLcv9hNWDKcbW0gfTiJcpAJ
E57pP0xRH2u9AOljzefFaZd0Vl0XWRBtUqXkkCSnBzDStWkEyGfGac080hTVp5TRWZ33Xe3l+eLI
L375T0ex0cFA1Vyzne3BI5pCnZ5tjN2aezo3X7CKTPeft2tQeGjV2BOqUq6vrR0u4nOtAp6ESQh7
wT2AVFplBQjkwavIK87OxYtN2Z5Pc+EdPDWssMdqQbSRZOAvwiU7RxkV6MfpSz7x7zT7C4R/NzUP
nYyPnot2ks9MXSqdvGW2SeS+8aXWZfAYAMMqQH1N5/fiejYAXLCLqZO055o9vKzJ3CzoxrV5C2Bw
Gv6o9hsuTAi5OCcvhSHEHprv3pxhDg4+mx+4qGb3NWbZTuFPGExCvhxeAmf9n3Ph1IXIUUAM7c/D
/vDr5fpz3qB3ar7A4RuDOpG5wxCUekKYVxR63tGDsre1PCxv93C7jUGzNCicHhZpVMRbCJLTeBVo
PwK+G+iASBdjqFk79biHgaF1jXp+w2z8NSpdHzIwo4TrgKs08/BpuVASfXUinT6r2e4AMQqAHiUk
ENGioHSBTrW4SLnAm3J6TIuSEJGVkx0tZLaXR2Wy5AbpGpu0NOVkVbag3Gbgs6UOb7LanR/ZrOkB
X1lUJEF+n7sOGNvlhTgjyyc3R4Eo4h+OqqrtR2X20roMyuFeIgPd8l8iIkT2NNaWox3ex3fnMYuJ
V5jrWepd4KeTVOayQtNfec1vBqNOuDRioJqJnVXeYOh2njkKf+1XJoYn2pWxl9qPfcQTwt5kVsVV
ahFbz7CVk55UBR0On8P0gkjHY/vGzPOjsLZiOMGD5e8wGHB1b48shTZUGu98rBHZytze0EMkbIWN
PVzIUE5AzzSFixfA1KwmgAHqCBA8N4ENn6gj2bvqaM6W6CuTT4qnjIMVwiBJuSwXrQ0fvwrpoAYV
Hqo28blL7ww3Gjc0qA5hb5b9hcozP1jiwCewINa3OzdxifQt2yS04KDgViK/HUjFT8yIdgBPotRs
PrvrfeyPvHLt7nN0xaXqO+tVFGhBdpp5oLlZJKLRZOMqXRrLcyWOyQxcZbCvNP8l/lSV/h6/ahyE
992konIYvFYHIExzrteb0xH1Shsvz1x70AZYqqIbhOr6sLTHcm49GKOW16p5+s5vAq2D4ESE/GGx
Vqyve4z8SfxLcc+P1l8ShupfyD8USQVwIyPM+ROO6UabPc/n5EVNorcmjHoVHPzuFG3r/iXfEZ+b
F8HYGRXp/WoFE8Kt+WZRz7JomJDMmt/8rA367ezkFXwKcjysKcBuUc0k88wGKZFTyFKgV3RUGz30
ECtXvvvw6Shq5f+VlC1Iy77irZp4EmaZTdyXqFh6l+Wt0K57JbRY8W19pdY3GR+Ly38hehPG4pYg
p2MrtS6DSHcAMdCEcXbAmgGc1OUIuu7YgP+7PRwHDzO4zMtqdigfnRjGii5K0/tiLlBEhjWRXfVA
U9HXGjr8q3IQVSdZT0cbzLy0v98PImqBNPuUY/GXZYywP8/fgOEGNhLqEZoL9CV4n3jqPq4RpNhK
hVhuU8s734qXKv10+7zU2Y1CohJF8+H0cixdvOcZBkczHLffQLE0lvbRXgr+0/M9WWutqe8VCDMC
cnucCuwg3mg05ICEwKa3eewyscghFOXBblypdkVTQtz1RQhqysS2AIUAlKCiSZwRUbrlOARR02FH
oYT08Ypv8e25x4hIaKocLkJ48clGsS7wccwQhzAS+lDROfTlpVC+fn94Z9hgogH8lncWKi2qkJVe
Rf7NEX9aHfAZ+dlZI024ncIj0JqNHXFPxoD/rDSM70ALvuWW03z9eZ+qAX+meB7e+rIxN3lti5SU
lT0sltA4w8akZRHrL5pS+tCX4ZnNXQhUM3zB8t5yy+xOItDTBJb+hV48rreEbUju/a7vB2hL6+0t
n4GRK1PkGbnnfXwdDDTqX9ujMrrSZ3OIvafApor+0EO4wERROBjGT9jIqSF/lmOJ4rp0WC+TKBIN
C4/3XAwFC2/iAJHN17/PjsUrnjiG+ZiTdXhfGxZ0ULRtpORnSlA7FEBWOj7XDmieKT7DlA2J4ulQ
SdPYBvm/+Sjm8Z9PRTqVAVga6ACj70gWG6Luwbon9wxsd3zMnPJ5eCAw+X2x8qwlz1mBgNJAZqNo
qszD6JTjNusFhmD7uzjVknlSmAaWbiXb+GDlE2g5LMchBRkuQF0UwcX6awDxfkPGPAKNriALA7YV
rmnm/oBvYfhatJ2UQXm3i+6hfqmluMiG4Z+pRu91dbYzflfgkR4I+/L/DHQ6qGEFME2uIpDvEjBm
/0k6J4zNEd25hzwt5DoV1GrQldCMQ9IHoogQ13S8wbrsC4viGhvFvpfEX40uvjOw1dvOpRjRiVxc
+BTx6OmJygrgifESRMZ1LBSV027TAO2B0NJzViJm72Na0um4UMha7T75Fe5yxAN1q6py9HcqaSAF
UDMbVechKsdzJhbL2J/QGA7LmVdYPHaoOTDan09UR/j/vfyBRUtK4ngTRjg+YRYIeA48jSH4+g3v
49lojkrVZVyJZ1kgTTB5tNGd4zIRp+rjPXyXkxUScp+trEvHQQAztb072sTLcp6phgF+ExFF/eze
M6S2MCUTzjOXzMeK9amQEl56AEm36GShHqO6t+O21hTWkV/QYDddl1d5N/K8cE4KCg3dFJeiSYKL
zmMBk543u+Dxnowg7UpZp/PRg88M49xRXkEKp7yLF5W2lUTrh2PIDAeUocfy2YUWGbn6T+ihCwb+
OdsWpfyAyrdlL66gqEKNXSpoj0dL6m3EXZeVdzyO/qMWqVbpjPXv6LomAGxJkmOU1c3C0UcpopWN
6ag3mgl8mZpmoNLvPIlB9KitZX5LPi0M4pE9q18qzV77cKp3bL82R+zfCEnup9n+V9gFCrlL/i81
5m2Mvm0pwkWn4GBXlD5YJsOWA5+hZCUPfs7hF3g7h7MCsS95T0RNmvw5Nlb3byBMKwIMhPOtbJQ7
vK/vxXfW6BYmGKmcyec5vqcbRn8DuUYiIU7LmCtEFcS9TK3yOi8dfvOaZB8jT3Ebx4X9/DKLkAuj
OPDJwEOfmG5mDb5cfviR98o1VJi8SIW1/PQkKV7GbKI1nPHVX0w2bctZg6IeGFa2ZlGh3oJmXKBN
ajl0/nS0JdbxdxHc1oAxMnWVBPrb8xt5vZIS86Og3laN2X6jutmvd9XRZncC1A8DaHsGFmxAFlIp
6Bubgvt1nreMPw0B94RrWFebocg1kBt2bsaREPGLNW42i4cWAd/eg7nep8V6cfgUSVCn306wn+IF
wDf/Dip53DABaIXL+S0kZ2Dwdx7QINZLWHzQZPZoB/5vbqVV+Q/sLb3TRQYiOm/GVUA1Sj7kfsEX
PIACitO2wNGnbENB8SKa51dUqPQzHAPmiVSD45mSKAkVhuNgQApyUwsyzwV1O//MY86Scp27iB+7
XLrnuMp6I7+1sQcyy0c0XKjB45j3nABKqG0Q4tZZjYo4tOIn3XEjUKmVUpMT8MLGafv+ND25MRdt
QN488d0m6lqlZZr7tMGjp7uzf6TJHITfaKN+2X0GcR/Q1G3mtXR7JekQIkRbf/eenvBvZEHkpgaV
Ii7tpIWGRnw7760MAQhNdSCjDjv0mx+h7LTw7HKH5CtBY1N2FayGzy86DoN2/3dafyEqjV/wS6XM
740YKAYJ4xQqRS3E7jpRcKHPQXKYcLg7U/yEW/eEgqzu9VOSgVuCTZQEMQ7p6RZ2B3loq1x7KrT+
uC7ZsmvxEyrH6J9KC7FLOk4p9LFiipU1c1MABYuVzFASNpSnFiNZsaVm9n6fh6yomoEM/FbxG6+0
4SNHoEobGpH8jI4oo0zfmQ1GsFIzjaBe9G3QkCOaUO9s6dDHnVSknTNcUe5lkFccbcr6RrsPsA2e
/S9fYmrCf5RY+61NrPwJn+ZO5JBFI5Ahfp7kFWkFeZm/C/BaiEgu0hrRKRL2C6BwLQxO+L76ZZMh
6SJbk8M9lVS4kpbh3zrzzjGKjIA6rgIaFH13vVbWcVCopn++WUUxsUUvs0mx2wTIbhEj8ja/RH/J
0yqyvyJSko203NL+TpINVfeQ6NbyB1nPPbwmBGskL8VjMOIo8BEDRO1/NzP3rVH8jXPJuyifjBNI
1Mj7Iv/eo3x3RR+Ia19BrIdQoaUDF/ICCJ3Zb081TlSH0fLO4RVZsEda9PovwzhPg688AWThvmra
py+ad4ZP47Dy8YS0ncaHVvlFEYV2YxSv3HmevG8sxFRCE3Q+PUtamh9h3+vBEAfgOZZHSQ/AfFAj
LHyW+z8zN/QScd5Ks2PJVP4WZ2XpoGujsqsowY15FC2EuNcJh39oWQY+08lWLMFwqPQQYFbr2Ue1
N5TZoyp+zoQjSzMCeuuiYhD682KuYiOHI6spX345QLkDNmlBeQ4+R+0THRUJAu+zksWpYDMs3Kuz
e/b7E9grXVx7M7t80UJgmJY3dM/Tybh0nPDOFniOWRdtuSeN+IADyvw4qR0h8a+0FFEmicGQ7sIm
SRUAISr4/BmgAPHk9JGHN/T8iIOKYyMCtCL5rrg0TEuZdWDVuzyt2mRkeV2x/QCbepAgvKFVTUgv
UJ3ybsvZgojBdd2VEXtVx5WNmlE3B+xbdAoSAwA17WQBqXTH6GseHdMUdyqpvkFzjP/sbk+4qNh3
3DryATTo3x4467f4x2iuCa5dNMXSI6mye17h9F43kiFV3nfh3J8AISyHN9QQcyAwk1vShxaDB9nw
GBwRJrlFtxq7FGaG2RbuE7PL68tU9WET+NAhCPOS/j6G1VydDAdPewD9LZ0iEsF8j1BmW+be3EfM
n/D/SZs6WyKtazYR4b34tIS6BzP+8qKa4632KEoP2GgRL7rtEg4S0lauI0z20llCZYbB5yVLZs8v
rMWTi9J29pl4f4pp70Mv3ziqr4ZbHwEBUi12BmuyrvNnAy4qH1+NMuj3NbmEw7hDEBzXb8VAceFy
9I3lBvuLJGOL6qGC8oWoeREDEORCzgm92j8Hx6L7Cr91LBTH+xc4EAosnJuwIs9HfhuE7yjNbSVT
RTvy6Xq2c3bMcPhXlGse/YPGWHVHwHw2azbjvAB02TQj7PSEB6A+pAUyc3Jsz7l0ZHfvom442Ytp
yfmuYaeZYhe631bYpAdUQCQfFBhmkMRm6jMDWhObuhMFyGkFO+cUc8mql5ryy/nWif++JSoMrJcf
nA6i9nHtm5AsdGo7uCAaJYa7BaX7lLjVLADDcrvJCOVQxPStCqOhlJZ5SDInA1GGrfOyu0D8NDHL
nbkUMqdHbQvokB3grTPIq9qoOUp31SgJHnHdJEr2Hh9KP3qWSBmzaqAoEtMh+kPXtzBYrmpdpJvk
bUen3w/l6itv/SI+bmt1SYN+kVbvxwDFJ0ME2PLhhXlx6rQky4zOHdgQ6q7rLXcNYIqMTxiWtjm7
67KfGUp5isDoMAeoiVzTqV4iW5SaKe0pdVfvAlvJDp7GfehfSG6tpXGKH8N43ZbrdMXxpRzxRmSn
u7CyHKNy7fonYaoRz81ONRc8DVUExZ5c+/4kWh4cfCYTP6+ronwQBEcIO3Qy7CwkQ/RKJeG8+Sl7
JSfef+58WFyYPBBa5/7vah/g0TvGJmzRbrSb0YwL4DHNm9V0UsRcg6VFWRRc+KwSA59JOtgujmHM
j38ILRpIhC4CxzhdaJ07obMYw7wz0eJWjmlOgtGJZ54vj5vNYG2s+vQ+w9NSSdO4tmLbj0y3Dl13
KOsJoRx/GvxxFemug0was/+spYscLQi1jV1PenJYZclJjk5QHagvnu2Vf7wAyUMESH3L78c7FSI5
ttbdx6W3aIgDuSGOB9lzfgOeaeEWMZgmeOGkKdgCO2K8P2glAH2U2g7mhn5e98ZFxgb/phSU1+4a
73fDM22jaVOdT9qqR3PlMIqnFkEDeNpT37eQzjjOap0ucPBLBdM3UCnvWVBn/Q19xjLW6VV3SU56
O4YxI9eV2hZ6nnNm4nZ3q9x8HuhtS5xupkTJ7AQ+2DcZSTJ5b3h03dZNIT6RY8kgyYB18G0bUFvR
E1geWRS+t+YJFYBItuZOJHsuoLmU8xiYKTE7DBFid3kAgPUgpz41Gpa/6fk0dVWprTaBkuo98gNu
p//xTU2qF9hRHKlux855w9C1VaY4djbKt1VePYv4cfFEK8gsSUEB6/5+WmTI+hw74I+HwumC6qGz
23Qa45Fatjyz7Cm7QCP3l4SnAgw+WCltjYq2TD9UDd9VvKYsgbaPeIuhU9ZPxwoHgQL1orglpUBh
YGGpkOX5NTJtjuRDwZzevXrIs43GfBXp3vJ1DldKdO+FAphZ/HC/OVVlViEzfanoyMHv/YUV0jka
QFbkPIvy3vRA9j96+q+OIWGq0pbP6iSgIbfHDlg0Fj/o96sYob6muzmr7biO5cqSihD9Ccs33/g+
vDvvcICvuaAb6prnKORTA934iIAw2ash+SmZfZnhWJNEkOqDcyVC5L1L3DyD7sUg9vboezAGVxHW
6T8XyUSnwD8eeVvYzMoptlNROVq4jbnxywxqP1xjB8kA1JXJ6CccXhELPzFiGN9f9qbeltfkC5QT
zhtHP6w3Fl16qPl98oYX0JGdc2VDbADUGG2w8LQLEVSRN/yYLrW4gJ7PqspJvkIkdgzIX2JNJNSs
iEmE3qnkKkL9vt1Jr0tgvu1Z+F/rBqADxtpzc5cjkYEW3IMIvYl/yOHlav9hCLM/xJ78eMjQZ2Se
jjk+jajcCFZwQIgwgF0I6XI6wRzp1t+2cqOfO6TFrCl/FDvAWyXmJ1VjIKKdv6+YIN14MmEjoDmq
+7lIGx+zvQ7JvDXuI6UGDRySYKc5e9EQ9ZjQcI0yxoeFmamJENRiZiYU8UfeZOw68X2z/TD8/uUo
D6AahkyrlyTusP9mRRw2zdOJNENtaqML/9/I+pnmpEX4Ru5sZAtsZ3JCtRp3jBTUeEjXRoJHlwXx
RgJIm+mt5DjandFIt3jej40fgUufjjKqDST6Aif4Ms2zHjXOnZyP//RHkUqPaydYsg/mERA3GZ15
XVEPdS/ZI/bN5tDJv+/bpt1jx105+9posLGDRB2s0xV9HZFdf84FrPkfClEh46doMCrhE4oh65V5
bv1sSQneXfLvVUkSj8HGkPOgrVF5iJW/fWwJI+4vGA4vKqIsxTXNKUP3d8GqiQR8YtqPyld2YuLQ
47aCx0fNnE1Kr+3J8CLlWqgZe4ulN+h4MD7zli0VXva1gUbei+sfTEPYYfjQCP3V4y4puyDQP0gc
c4hIzNNjOHUXzaeW+Oh0bJIGljCXVy9dboSdF2HaDRR2+SO4YuqcMAn+//gbg1eSIgLD44xUIbBp
BWmEZXOojIbCrYpY35FHXQQDzKnBq4UrqasYKQPND8qNVtaRXGNezvU4LSTGzH2761AgnjZS6I30
1yHTpwjRioGe9UDime1/X1snG2vTVQ7HtL+Cd6hOwz3wAgHHCMBMQdlbmAiE+mLoXVATlW9sBVNk
6oqvqhKWldTd977Tqo0Tgf1smPsIsZHosKZ3GucrfjIIhpZ+a0iAfUEkBVsI7+4JzEfAVnSDMDwJ
62UHxXHbYXeCSBOrClSSi1fifM2CP6eTn4PQN0v+nbzw+yuYQVMHOvB5H6tsm/TxTSor3KeSaHAQ
wD1YN90QbWfj4/vqVldla1G6ne2nW2t9dsExEuYuuMA9aUaa9RCbbpL0VOhA5XpNZQY1Em3O3nPj
zay8TXC9xNKWR2B1FiafwXGx+XDdouFt7rMUu1F65bLmpz0BG6MdwgkaHSLJvMPWWrJ/l4Tl8q8c
h53MizY3EBVKH7tDYJwbHIehZweQh5/kmVe5+VoG38pzJrapEUc0XuncC3upUH3h+XwO2Zlc4qtk
j2bgktoJufCByppNk+zQ6sMvGlEKMPNLW6o5ixbbo5glfpFY9r6zmqRIvq1aQb5J72jMOdpX5XrW
oFqM5jiaEkExmc9ID2TQy9m+0UDl6eXNL7zkC0NlfWdGk2T7tt4IuhzggPZg6sCTYG7AtCpt36DR
72mK8oN+0QkrxOFUSvwwm1Ecatv/3x49gDM4mO54Vvw0w50mlXXY1PdgiaJsUw7DI0CxCyGq+Sq/
6cq4X31dtm/JUsIK8rCqSCZU+ZkIWXKs31TT20wH0vqatNCWdrXum0pj+dvWuiFUWvBovDABXRwB
+G4BsndPJhOq9GYHwtJ5BMP+Mw2wLIWmyq2vM1HjEcf4TsFY/VNniNW/mcYAbxT2bRcTbE9d0U0n
bZ7h1zx7nA6xA1OeZsIQgQWYs0Scr3eYuIraN9FSyNWvqXkqn9tXcm68Qpfj6ARybox/NmErZ5r3
0rvxvHzYIzNC/yFo57LIHRCaNoky9r8G3x/jvVCiRjdYQUqjZHD9kD4Ev4DHW4fzYll17vQEyPag
Q32Lt0Xfa/5qYsfXim8Z0zOtk46A4X/5shBVNMgHkFYF7bSz+NOcC1SwM0FHUWUQB+EDQIXhiqN5
aSK/ltwkhScecvAMVPRpC7fK/DU8XW/ZCIbDY0wyCkmGzbobO5igwbThHZz568qzpv4u4ZliOesj
f6Bd4sAdj8dE91gydt7PyANFb5IjpZNQjR4FiwE9Bffyqh6l3Sjn3UXEzJSWijavynJRp4Jal/Y8
JQ5SxImKv4b0/u7V8KA78X6lORpHYjcH68qE5CCmTj/agZp5656Q9GlEaaAR8GKCsutgkJIRy9kN
bhWX2WhwdOB89Drr5auqAo2SZLwh4CuRBocfLSQJXp7e25s4HrwhAyuNCWRQMfXOCPQpQVf8Qxlf
BUSuh7B1sWcQFPbpLokaiPC8/slDX3oZndEcVtgV1l8T7SdTTwp8YkIxq5euJmPt2aKYevjgr4CN
/hhNL66eg0Fi5GbNMa/sfslGpVwynOm/QmZkAsOBxNspxurfleJikxSTUXO4uqu3o6E28YRhh6P1
160FoV3RrbzVQGAHBDwF3FRpCZcgdfGxus9uJnxNaIKVagjKeCDpLy54kvHMa+UzUR0lctpuKArG
pKN7nmwVvXY0foYwbGNXxSsGGEybp2kyDY9bt8uk9jrz2flaFJDSMJr+py4U0lisDgQj4cMmAMat
/eSApBdrIBoU+CxwM2ugwCKriEW8j043j/V7/74q9iAtD1IZz0Eiswem/+z0EwIZH7PZvzqXpnbU
CdIL77H788PTW0QW5wuAV5njaFOwG9/RsbNMC5xewjD0VhcKddY3Um6WjaYinKtS0JGJaqaF8MmK
BtAt8i0AC9xetBKDQvt2TcF1nXUo2PYVEhKi3eO4ujW0spSRtGb15AgnK8vHrX9kcugc7+RmEX0b
Hw2mskBEW+tb3A8btNsf93zpGTDqU/wilu2sjiTbHBqn0wfFeQyLKkuUyB5gPTJRpxOsaXEApwte
zdU6R+ert2ocDq5VzzkLiTx933bVKCMYn2TFwrpvPCIko25+ezeI7jbkudVoFnHkkjj9p4GKNtPM
C51eb6vaAt8IHZ5KQkCYdjcWRJ3kdoeeLeGIT+djZCCScdh+1i+C/OuFycS575BB6gHjNgtTCUNm
+JZ0w6AjRig2IaF1dTLXfR0EK7BPI3pMwrnmh1MlA5uL5lVDiiWBrskNVqHdAzzgc4pV+aNjzS46
BeKR0ZtSbVdyZHKsFmMp8WRqg2/Exiu0Kk7PvZNhoW0MFSfDQ+LpTwJaMaMDsoys/1t4/B+m9/5K
0SdqbkoEpJyHO5gG/MIFit1wGAv0tE1BjztRmoiwqAUcHyOVdj3Gm4Pkhl8EImpOCqjhX0A6T94p
wEU3GyI2nb/cwVAlA22DVEwATBRGngGiiozQL5l6Gwmvlm5CO8+IXGqPH3ptYHpUmNUB8t2G+KqF
yhJVszm2hmztn8OtVq1+aIgJeqRPtD66IzxLiGIHXFz9vbKLvuMtiddcH5T1AOkLPcVkkQw+AFJ/
RcISgWgWQtLbXSIK+5V1NUxmwD5l4cAluasmyQfmOB7cLtPGh6k56nhKBIJAip01tzKqXapJC8F8
MEikyCWCMjGpSkWTMecNvJvLwBn90jE/RjdmvCxVHLfb0R1uswLbYSov6O/b9s39sQo/g+Q7GS1/
modaQrWF6cDB8l4qm5fKEYhuTkZ37qUdqkrk3T01DfnOMPB6hDyngg57wSH5iPbON7JlMxIWZ5Bi
uPHhyMVTAdmom7N3lB0fPlhrrIZZjueO5oXRcaq1Imfu5Ro9Mbxu/SguMZnCtCs0hiSEN0R6crtx
IGjZlbfpFYj/5Tpd7YPJfXv/Vqx0X7yMycY/rBReTc0GKZywydBLM3XAYvktmaBk32V9Vq+6AKT1
ptkkUT9W2NNkxHfFIq9yHa0huAsz1Qi9xzsSKhdWheSPNqHnlbAo6ouxEW5mL+fN8Q4fsBZunsdu
/acwf49Z2Tn0G4NXTgiAeZfnRiDa5BGY1fZdtcChPMafjUcU99+KFYTPksOLz5yBGgWlNdXPXtCk
18BfZlAOpIVMecSjf/IRCYVuVKWin0LrgAE9WxEl1ojrYfzq4cehmWss1KmLo2y9AAPvBCvRZitJ
Q19jMf6vPMMOpVN7J3QqPVC4oP1RbunuriD7bNKht9JIM8N//x4W5vX3noDjrzJhoRdWuSyKcf1t
sYNKzh6AoIiDfHVpHW8sSamrf/Us+UZeqPvNDvZd8AbinfOk7tKdc+ojkNnwA2mRVMxRDgbrScwV
QhHsSrBcOiH6QlDRc0zqmH+D9B8tYJV7j0T9bsTLcPJ8yzuzK2LD0h4itMJpQ5uON6nA6B9qjmId
oMe8Y3HKQZKDbfTe0T2PgnBT2gXJ25M99Sj2axTdjPol/gVfO/JNJ03QNnQC3VlygUSYBsm1Ke9X
hNZc+3JCrBUVDRAeg/DFDOha/bTKnWcW+T+Nwbf/nvPh/YIH/QwQZPMPBe7bkXFQu/KFSElXyynf
XV7mfj3CaxZb84+KK3L7rXsTG3Nls452hGJ7TBdhml8fO/EsZs0QovNztQerz6Z/DxFB8A1yyJF5
QtiGAZlIPuHCWgMK5Gl2NMi456yTYc2dygc6XdCSOMJxnwK2P2TjtnGqk/2+Iis3KlowQHDFuz1L
DzI+SV6y1Rvp8Jt/fnTHhEKFXO04WTi9CRyuFL056fA/JMO3Ynv4UtzWWx42PTp9f41zPVVSlm5t
KvJBOJEkQbvx0iGOZ/hCBt+FV1Td5vin4E+hX7YX1KHLgYe1X1HV6F2sS6Lu1RtcHG95kZ0On3d0
b/MxZJPk5mMfiDAgKZDfL2o7QrszsZfPpPVkEfq9cIa0ESAajM2Y7O6KgJDU2VC0GZ7r/1NmCCvs
JlESkIbTT4dAqpr+RTMcigf4qrVB1dAVIV4G4c3QTvWHeLxMLhHLhMWTRPEQz6jFhuHJmFuvVXG9
1xN6D/cV4JSL5oFECYHuw7eatvzMbIgsWoesP+BeB/pUFRRyarTXKoYnQz1eQM6/UbJ3OAFFFoJZ
utnb2f481TQHmKs8tDnrhG8a6XQP/zZXoKNLXZaGwuyOT2hNJcB9u0jON+cf19HvQXQph7G0MpPL
Vdeft2+vC2bKcQBR9gcUh1Dc9YDtypZ4b31PRPMKGtkAOL/wwYHLK2f5maf2ROwBjUwXLry/XcEu
5bPFJtEBLY5VGcq0aERJNbbk2Gna6V6PphKAu8/1FsrDidhRMI6RqsGZiZI5G+Uq6zIp9SWMJH5o
xo2EvAZJV+y8eJ6KIksfQUH9wsv4nDI4/oIBXMnoLUydqF260HVeX4zz0KkcPiou3x7hfA11/AhF
Dkuwa+dqbIyajCU1NGRdlsrMybTZJEeCIJYfISTYsyt7RbDHExNQLuWUIcqePs2h8oYAae7qPps9
HZLyzS4f/Vl4fjwWleIoWcRrCPmxsYSbLPWNJec5SHtYMq1HRBDuJz0OAk/oYdZWwwOiIiDJl8RZ
wLyb5F3SRUL/AogvLtWaLh/+7UqjFfeAYnOSm3QFfFbzeFCRXLmZFk1IpOeAx6jziel0Zc/340MC
PIIlbEkZ/daTc3Qr6M38SG21b/j8298JxIPrQp1M/imkMjhRPEPwdIBQhhbbwucUEq2NMuK/lG4i
G3L6YRv8YENTJJwULdm644wrHqq9laIFp66a3oS3PHbHSZvfmU6kPm49tXHtc7M1oc/1sledCrPv
WZJkiWJUIUhTXindzq3DgwkwGGIAdR3FhDGv+huCA/2kY/l4NVk4Poza5HF8ZrKIOmjhTr670OFN
5TW02NE0t/nz6aVpeHWYlQ7xcqk/D6tU3KJqc4KiXhq3kdh1B6BG3NETMJaTkePrARl44V7FjcQG
fgqgfzmxJzdQjz8IjZH+Kdoiqqg7jeP8dwZzNFeKYb73ndI2/qKRPnj3fLkYb3BsW/vEEZ+SgWSR
QkVZ6EUEnDXOkGBxaJ6B9V75H4RI3QoVSDTR6E8VUsw8mpLEpjMM3Vv0H39+TsftQXUDmakhVMra
GtemYgiZYGdEDkd1xwwKFTSacigNYi5RC+jjIMZfpaATkLpYEA6a5WK/KgarrNBh9DPNHgb4mJ/H
qyMA8Z/IOg7N703ZmIco5r2jparBOIjltKiFYFCQkJe36oeuQZiRsBvo2n1MQqGfQvxsPLIJtIlW
drShupNB8fD+ksVbWGuVVZ7Eth6rcxwK7o6qC8221JDOWu46wbClb9z2yzpe/pKEP3wUmT0YAwoJ
fDsSHP7GghxvAQ7xk7NcxejjKOWKtWHx7sQt8sADMiX15F9Kb7LoRenFbzRZ/yJIbGOznXbkX3Sd
yBy2QVbr6zDYrxYq3qhuvBYJgXNG6fPJ0rKH5+IpqOYtJHoOM+9k2ztEOw2ZAuRWS7ldXFdxExFI
kH5OsqIwzMV7OGU9G6lFzCP26rAFIN511QOL5ApOysYFxlEiaPzPwqij1fcjF3xWnc8FUr4lmFKO
y8W1fg6hzAJBOcmJtScXBcHW0QHJKY6RdaZRz5PB2SgbEBx1E2D59pmxPFll77qldSCVmZjfrslJ
W44nZ7OZxsjmUi9Yecl+gnX2BEnTVvYMbheVAZ9bXrajyQLheuLQm70/UG21Cq0qKrMTQWhax/La
KBsg2WBat+XaSUY4l7qkKRFyZHY9bii/2C2bwNc5Q6Q+sdsTRDUC1XykM4VXjU82LtuX1Jvs4Ssw
UyKZ6d904/tGVOeY/51Joclfe0Yd5ramrHdHwnyyI6pIQuTTPVMYG4jyP/3Fr3eywJ03OdTCaoiq
++QdTtOza6mwZARt5T9ONMq9+4ZjM1sVuRndBjTzEiQo80YRJYStifu6RFZTwD9Fh3eKSD2o0wIx
6YFQOXR75+Qllbm7EEkdTf5U8zs64rNgai0o2LCk6p8PQqluQhqNsH5B6QbIRW54DcOK6D+E6VZ6
Jilew7es5oYkwky/4Ew+YRc0d957AiJPQ865JuKqwMwLGgPPoPpIso5w+DBSgnNQ39e3V4ndqh4D
EV5FOFLUmRYWTFBw61QhE6lxE3qOGToOmPNWbhILEgY3Y7YHdh0ji9fpYX4Erz9RENlhZCKrts1w
4PKuIXpQTS67j/oQugArcvvKaUr5EatLzvmYdCeML9Zdqrkm01DphWq1fH3CwsBlMPZyyLesCt9q
9fyq/suZDlgHKd27kzKMS31USuF1XWKlTW441zcEXxzw65ZQEaprFPoZauh6qfNDpSrXFvQ7eUII
ZgpquK8XANwLN99WjIELgZUfFhLI8gvnuyMX4TCXWNpRr4woXYqH0ST2FgxuH1WAVrD6+EAoGftR
aa3wvqOuEqkdlaVi+huLktAXVd+5fgty0CpaDvu4qHcOwYqZzc1IM5kwt1dIc5hTZYzmRI5gHiRW
Vb0pfako/VzUuwL8pJ0fq4EAK9CvsNIegeZhUL/0k9yDqJ6KNn78UwZ8llxoR/mlDJ8iBHBWUuju
WjJvPmfxYfz1QexWxM8SjS4aYXBQRumflMddWTFmm2Y3sAV9bf1qJ5M5Ittv6LMTAZuKnxygFxUn
5HGdhNHhg0gWUv/wcSQQkgO+nQJIiNfwUVBcFzvWhi3eOiiIydpeoRdLNugsoGkib/QKzjTwaI4a
jQTwvQtOS7GY8sEzHHHhGhHFicGSrpURzy1yt63JxfpMm+RW+bygY8rPT1c7DYja8eEmO2vbrXS9
Bs8vDvSMY8yqi9UHXYgvuxFj9I9NPQqdLt1Ws7wf4vZ4z2LMlO7qdDsVmkXYfR3dGUrL9+maeeMT
Wi1skcIZaXyryErttf4lS5T6tg+rq4bgLO7FJI93bJLoHFHPUdsvC2CugL7gKMgHY/E1V51zhGAU
H9WOEL1iSEuw81YM+P+NggT97UGRFplpgfGFvuFscMqgIMrnXA//zYAL2eC7TuvavpsQz7kbivxN
OiTjFpcAIKC/nLCNBbUFWlBNjAyjVM/hwKbiQD1paEmyJppUxHIAg6zZbShzsLSWwXH7BnFZ1rkA
AX05ZW8XB8P/zz3Dssi3jULmx37aRUrC4SjH4jRkmFdaSSX37cVisjskI9CaxduAYdfVE6uHxHkr
uCj1CbIIbWjL8SQraR9oduWEouCJzzDsKPqiVhCY6nS/Y0ZFhap3Yukc5271dsi6MPhvhoVi3YvR
AjjLR/ygVZ1HjYWbbz9dSjBbon3dJnpCVlbWs2zzN+h9QhKu4Dzjv0wWH216FhLtSCn7KpLJrPm7
4IYeyo9aquWQtApjzSaNQwVfH6+I45FSgmxdGMFXaWenbzJPgmALpyHnPfuxs2G2gefo2dqDzNx2
cwlEzPjgGkp1bQIvQNOATY9b3eWwA4PN6VAbGtssTITlbZI+m3EMPZug/X9PLDGWYvQwO3r5Skdo
/E4UQ7wTlPmhnBc761PtHjyzRtaio3Og22WIEk11A3e/DK0U0t2onziD7CC+rNiMKqUqis6bflnd
6lAZdMglUzeOmE+cXAAsKupRqw4BPy0YBVr8190PtPvvAkGbNCQsW/+yFgnpOYcHrB2Hgm4I4rJL
1DmN4j7v6GN25gOHPscFveF2CeLieTugbSCrCLs5S038Wy0iqEfD5+My31Hpow0dxCM3NJiJXCgm
gtSWhWHcU1OIWxtKXAUdNWaWAKIhAMwjLUj6oNRCZFe6HfuDQC8uUjIyueWswPBtL5+kzPFyAwVw
kVQLhwIuv/aR4h88YpZwF/V1SnPX2eHHtUUh7Eymt5Y6FNSiSqZevc/+6+1oAlcvrsrfqJpFm4zd
5Yz6hepINGGE9c2CNJjbjz3Ff5FU84+cWK7UmyxgNxJiMUhp9P1hJ+j/pEm2/9UpV30MKj62hlOs
HNw/TLzTIRSXVTuWt2DQVO5DAK84Z9Hc6V2w5uSUJulHn8QKGyxjhFjNTlY0FpvhT5apXzrbLZI0
/tfJ3k/Ozq8646hFKlt0rmPdnvm1Yr7NGaN6Bvg1GIU26cAWkr59opb0IzmTTTyFsuZa8k1oCwBJ
K8R9X5TvISDpqkcWAo1DBR48rrZDLyf2DidzObbPWQm/MYhHjyf10KSvU5naQPtCiYJRXX099Lfy
aHg7iK1s5p6uCPaXUbsbSrgZrdBJD08nN4EpcyZ8rztLAI7wrdd0vyuiR/fist3mRIFjvB/6lTUC
qNzqSqw8Kb7LxYoMI+uKtrflFdslt81ZSPfZUleQ9vpxodCQ5nlfVO3ZI/aD7yZIsvgkTASWv97z
kAhWnWE/oWjTTybXlgbNdf70O9HsE38W74ArzuQRCHQWOxJoRqB7ikWr5AdaDeOsdr0f/AOhfCrn
yCwcEKIPYs4FNd7pEET6ifBUQzPZewjqYOnMc9boJHJBPeBrR9+Z32H/6/wULI7Wi1dx1mPPP6F5
R2XZashfV9XcTpDvMV5boAQuPeL5z5FAyu+OjydTt6anwcbfF9ex3UKI4JeRwgAEhG5kuiNFeDTZ
Fhvkz/VTm2zSWxl61WIcu4w+1znZC68GdY2kVg9+MadneVDKOjDBPWcD3530W0qZBkQNeDuvSCf5
PrgUDMWKvEuxD9HaFezmAowMur472Nq+Akt3MxeEm8DS+DA7HaAfcyul0mWYY9m4GpwA9NjkzvVT
E1/slzTUTFQhPx7XUu2OOIgv6LLhWM/u+tQO5qbwX75y95CRvsaqNEle2EhXy4fSqpIaXcsZ6Rtk
NHjLcmQg7KTgTiand7XFi6xTV4CSNPsycZJNVFmqGL2p+k/VFimfTKuOAWrEHT1zrnunjLRvRgSL
8sYIV9ifUEgdH8NI+8yvUALMDwegj3UkaB+wYDGfszCe7abqr3ww8uj7ryNvU31tj+5I5bJcfCEl
0/RheDGRub67l3V/XplTTtZS+cwLnsyE85HL82s/xXbBshvRm+5zybe/OBqwlgVgiGSE+8vfYtSS
F6FzG5HxgmFwajxue0D2Xo0tsKbl7MrSwCqkjJnw6QCd6DU0QGd6GtV1w+pc4N7qkbEXdtfeDnow
AXW2daj+k6XKaearQW+R/usZGj7ZNB6UG4hu0KAIvI4gUF6UydlZoVOU0iHZqZ5ve+8xSzwLAAi4
+D0hWSrf41fMayM2+TfmUVXJAeEQ40JGzc5u+QFUVLmcuj2hMzsknZXsjPQV4mU3ziezghve4ZM9
ZCGs7OTQk9FOh2sYbON6ak+8P4SeepF2doO0xXCLO1+piuKeTtWMTNsdVKwPhyXwUCBC80u7FuZP
umVgHLgVNFZb5nxNdMhlif1+EuA2cy41FUg0N3S/EmXU5Go8C0LFlzm0Jbx+QAu+Z3I/W6QyrI3x
ye2llc7uYZwVxiJvU4X5mp8pchCtnjkp1RvFh7meD8lk4YzZjJHPtEbPY79cYniHleaOtJ3Nl0g9
Pfg0rTVKyY9F1VvlohuTJCKErPS7xJgukdo/TnnZrWkyth7jjG4Wfo/IlazJHiz9tYjg5l/ydYgX
EIgQ64SaZt+V5E8ZWIsvwsfhkzTN0fFeLyIEaeZMsthwMc/SYQEVFQFm90hYct1YISFDqaDDqQoJ
cv5LkwJFgMtXUH9w7xytFy3ygIJ8B1qrSC/s2PcyDRLHncvvwV0qbuKPJMxq4axxXubiQgvK+Oie
9Ao5GpBBY78W/KiLSaHgYNH14S7023ZxqDWt2JEsvFVGdmnuiPzDGRLNDZfBU0JVl4VdUDRdbc86
xzrt6tb1xMouFnSKOBU6MhH0XGff3AeitV87oeEKv3KfhWZwf0ObfQeuOkdD8LMCqzencdGps6oW
Z7FF7gmkerMlJRvgNcVIdQiGfm8qJQ6HjSgYTNxgmbkGKT6Uk689fG+lDELCSaNOuVxsr9Si58kZ
XMxcpGMDaam4eJKpdKZYx3Jf1WVPm3gSZkrnmlB/e9zVR1nCQop81XjcAxV9faStMLo3rGKsQqdt
4OaYbC9WcmMsRX8Xem//wtiEXtvbOWnzIzRz7LzVSWe2WyhJPiaA1d/ri6b3ykmTY3ELD7TiZybX
D1KFs1cIuXjY+BuSNrS7/jdfYlBL5zi0ixfPqYEDHYX0RAxxA2/GXRPC0kqynbbwUQde/HPkrBEH
QDoO8yTTKqNwFuWWojl2y8NK0+1k2Xt54T9n6+sqyq58Er8yZrxCsY9kBcDGjxYuumYXhFsztryF
+1eWGUdo8MsBtTuPsJRpzH4PefG7lLyOsu1uKOdgM4xLzKcnYKoVMq18uZEYykurVFBcb37CeKM3
dI3UY6skqDrDdyPkuvOrIi+TXMWX9nB1qlwH0q5pcIs+I9LsGrPkJStS+ZvLxreBMnYhP8705zxL
UmpeIF2ecf7hlC2ojFeaIyzPZOhwJgb1I9fS1qVrxwU7A3Rc3/WFoD/59zvNj6mrGNWxLIIOL2Kl
pkUV1jC9oslDokG5+qzm3ELp3G6yjWoxUeGrGJwXemynX50xZvcnSYPKYNQXot/Szps6PMzAf1er
Uwl8L88D54WtiOEmbUt0b5PBDymOEwWFQrvXYSxt/lXg4ELIusUOsZGTAusXyqjUvEkpIHkcfxpV
tuvoaiLqQBqqQa43E7ocj/4USm2lcb/T3WW4ekYmk2lltdKU4xWgyQw862GmJdcQYYL3Qy0dLw5Z
qbTWSnqsn8fv/Rl6IiNXXd96IeQwSbZTXfi6nemx37wT2qZ9XnriucKLY/Z1SoCap5cBdEMs5CQN
qNr85tfuDp7ctrXhgfeVJJo9kyyzQw56JyI0KL3attxO8p9hGLowXuZMvFqHLG8FR/X/WZVEUoNq
/aafjHTK2350mjXCKq+UnKpDjDSlLcEHJrYDOhisLm0Lbb2Q+AnLYeGDHPpizOk/xqbEcKqDvSWQ
6xhTzvCyvYSh8mIWsQ2E6F3AA09BT8EMa9Ktbndv7O5cp8gxdCuRurjCG1clDGTgBJCh4Y/v5BhB
EiCd9Vp8OXZ+yqaiHSgwQYMT8C8TynSfxMy3q092U/nRQ1dZCpL40GeooUrpdPp+YV2KzRlEGbCO
98uxXjakRNt14suPW6dsTYddIeN+qWsgN3eJGgyDZQ4lV7Mjh9/uNS+2e7PMbitkB9R8yTm75mJ0
qSV1arEIDA1tQTPwzlQqJfioPRusXsEZGWPVFsoN0evwWJ9ZjujLD/MZS09zDT7rPQsdmgsYn133
jzOvC2laVzDstNk4MNilcUFAhyyg5o6EUko0aXaDZJzfGc5qi7oyx67V08OYFHd5hrbDRkNgDJix
EIxRCeeCTXPPYWj2CgK1xdMxZ76yFW+eXIkIxcUct+cOXI4sEJUXR4J5Wlk38abL8XTBUT0G9i5D
jO0xbbJpTVJ8h+DTUPtqZf9nQh5ICz2NoNzO1O7niIIUp4pmNG3wzOB3c2V4dZFo2RP1ZSvzRj7p
2HC/eKUbov2HlpIt0coapZ6Qk/5rl3QVux2vs5kGCHfHhYFyyaYoC5vWBVVXvUEf/7irYSUYoQXc
H0QujMcinqRXSOm7bh6mTz8P9HcYPRcs2YrL9MzrwcKJfzJgfI1ySABVVaXq/7priKxNJf9Z82Wa
ejt+HtA/0Eb0/5kxJRTd5wxQQCd9CMpA5honJK38heDBIuZixjg8NelLQ9MA+595cXsJYq0cXhIP
8zPJNUU+QlwhmTbKAzUc8qgo7+WBsGAeH03ro6JSJvJiaB0kyhtUrcdXsgp7z3chCMXQJS0LuD4O
RBkn3t8u33et5w/uxtO8ZDJgralBK1zJYgfl8bKZ+NMO7ENtqGCOfKX+pcH0yzIG5R6S2Kx0WJ+K
WioiPXBNBYUXLBhGH4lXhJS1LYcHSQEok3rfdYq0+9Yc8+tzXLphDaF1psKsgrXDKM7JO6tHOn75
IF8dsWWKCO7W0hxBQ01Q1QTXClXWWPKk3/JPwr0U5J1fmimCCJqbiklSwQAYpNkeJOttR64zEC5p
IfEWz18ZbIDzG8FTstvCAmKZiLKcNVCxzYkPnWJks4MNDH1Vgy950IfrwbGu/3zEGS28BkKryeNA
kV7d9KOrK0sxTX1caTHsDkCvchpaaK1TnGExRRPMksYUw+G4N8wEy61v9ZERCa4ZQ5moE+cbyTSi
GaW06yH1YiJKkc50+GH83eXoIqnymgNypvzSzBw7tLnqYYQHZ+v5b/CduO6inoAfGDw2+ZC4d2JU
PCgTN7kL1w1LTgMVJ/r1Zo9AZ9Rt0ZcRt9J+/y12T8c+OHysVBPLkMNStWl3mANZMgf/AWQcdtjp
rAopeO5+Temxo5YYM6KYHBQTgg3AhRnNwVXBRxc3L6XbnaRpWtNYSC0DN+pjADYbLhTzOJMsEhCt
ap1r/9yn/X/cmCqR0OwkLxOYtfVDqD6n/5TD/m+xpGMA5vdnllTytctdgpi/3WIjeYCkFUTWY3uf
5BN6MrmuSwto4pgr4rKuyGuBrornzF1hajj502JRsT8EjMC4/DycmaYjt78pa7SwS81XWPpphK0X
9xqHqSvrucl2iVqEKVk8vNrxHLHWh1jAESdssIJUmqgVM50gcMYZgWM48DQnnLEpMjfqInSwMcKd
CduFUwZ9nFcVXoQ6laeOYyudziD5SWLq9Yp9ZZx5zvbuDQ03AxuydYTeUTncCZWG+YetzKJPCIK0
S8t5TmQZHns8ZUpuevfApwvoTzMfDcXamJwl/SvkKSV+HmvLU/CSFRlAhjiq4xXw/72fyjcIWGfN
LyHfML2HwuXos107mcCdTyk/jCS6fkjXEqWvu9LGBXmm2TApRbgnWv6CpuqBTSAzkyOOZL1V8QYC
THbS2qlxg8ILMohqJTgHjiGSx3tgFfCQsU6U2jq7MRiJtRvWwYNQcHCE2uP2m2iWO7BFbJ3p9W3v
rVRoUeCefXNiK9c1rXhAwaIQr76cI4FXf9+vOsoTUeE9o75fmNmhb++hF3iwHMspi5yBxj4hTKF9
3MjVFAyt1lYNyaaNLyLASi7yZI3g7ctCTwiftVoHioOl08PggV9/IomF9vN/pK6c8WD76RzsXgNv
CJRSXve2tNrKCg6hORr2Lch4VqMyCVp1Bk3GrhVJ7+K3MS8HVeVUIQ0L6hVkGdhfuXd1fa/BHlON
Bxxo1uHIS8BiPvH23VWzuuKXbjSWQIwtd7ePZ9i8Ubz+tEBO1xK3po4X40pCKa/E4l675mfJeO3y
kzJul5ELnP9AoYOP2eEQPp4wFZ5bnVMNKIqoqn2+8TC2x5O3+jGLlL24VYfrT/JPTFMkTi3YPnuc
O392xb5RlKU0FxxnsIrefRo4SSElW8VvksPbsDWaTHYWR5lvs/jNbB24uvXZ++HQBzzpXqtI/lEZ
FU9jwKbxs+SmX+NR+AQjsDp5CsvERVsJZoEYd5DB8WXzIVsqBtAJ+cI7bNS9CwxoSXGsNJGNljvC
nZ/8Ru9fIYx4pBNTv+Ziw0QH3xMFVYlXo+wIPxEpX49Q89sFsGdB/Wwna6tq8h2Q29WtaSh7xBEj
LqcwWjx+lI3hfmvdQrh8DDg8wBZ6Ze/zhbCJPk2PQ+smSbieKl5Fir0UDX+/QdEaKscrwXievmjV
2YbATYLtSoaaao+/VScoeQKDIsJFivEU4kgjb0FmNcKfpzKPaKjlTrLsggNtZDWpjCS5bWaBd9fW
Gu815IiIGCXTc3I6/vrjfDfChXfsI1A+Z+k8P/4NfHNv6aHzDzvhGrue7tiXN3mOwWmTCD+dO71i
HXERLtoh13O1sjh6evP+OM7C4Z7OiJwbndwIxT27Pt9fqEYI3FPH5qK0eYiTmuTp9nYiB8P0b2Ab
l35dVjHy2eJ+ICgqFrog3tOzjFA/vfAvqlulgN9x1AJmsNQkP3PE+tAqcZTPnOquXRaIj/K6shv+
PPhcncZql7Qo/bu0WMXEqiPw0anrLmel9fi4FvNjjAuTLjTlaBqjBUij1ExnU665C6L8NUHbEqWv
ew0azXSjkK/0nEtpeN/CJryeCnh4zsukOH/TnL+IMCAS6wivohdbiBm/mAY0aIR//qKCZ7lzkSEu
Vq0Xbf42tTjLUWdt1gPDiTAAYTGx0MtVfOrmfRXeX+gBvViiLc8M66VWzJV7X9vDbwgH0H3SA10+
9iG4RiCROKo2oOpnA96HN0nRG72wTyU8Uu9D85MxZyltgKBuRSNv+zNqz0+N+xXqwb1+HnsEsu/j
Qvz7IOiu4rwrLrbtqQjJBXT4mg949BSSwjnS8MpNBNlQ8+NKLyFJfmGpDdrdzv3Xt2aWuMMFJc5H
EGcQ9IkDFr/Nc41gH/qvFc1XXP4UIbce/kZlAn+J9aD+XsNjC4rxSPTXA0296pvFF86Vkaf4Kk2y
14j+fEPHHdCpERxR06tn6iuGEaMB6Vb2FMPZss6ULNI9sUpNZVGOpVD1J10D4Fsv7bRkkX+41tji
FIQxrGSPbJoviZUmsZYhyiOnWJCeauF3Cvr98JdHhAS/XscnSkjW8cGfU/qMSMDgAVSJZJ1W73hY
p+pWUPdwlQ6hMycdpGCW2s0M8FOVeK8e95JmhGNhRk2SK/nORDYqaKwUf4DgBJHZEuWZx5e6hB3M
wpgKcLb7UQ0/6mABgIkGJQK5Yt3ODjkF6481kJXA5FaulAT7we6BGAWcRSLBR2xV24Iqfgb8aLDY
xKvCvV3N4svrefSxqK+sqIkzs4FBL4lrA3jW2LvkD9dpzw55hthHZJkxlcqnflkBzyxOFNyYUkv4
XAV9HcsQX/IkRMh79FE6z5hRZMK3fP+e/geVLrJAdRAMLImNiO8gnpBdzAqJRGotPfO0W5NvJ1mX
xMdwETe7nF50+QWtvgXamDR4sU8Wllskeu9MGOBXYWV5a/obzsrH73Vd8cMBALgE25XnDP6CO9nw
wrK1GjzaLVHNT3l/5s3yrKgRnNfaxbIckl7OhtkSSso6dQfOX5o6ykeqFnv1Fssa6hg/mCpdfoji
bFqiS8QOaFnuiTdywfEQ8XKYM0pPCMxwVbvXsOhGuq/BiC6Z/5AAb9nUljB0+ZxPvr+MC8IhWVz+
ko4RRNW4llEv+cYKDwkWWwy5EZW8X9YlmlHzivz77XjMcJZ0+S0n1pD67zaRlNqVERfJEwufAZfI
CnIxnQc06ZeugH5N/Qz6q5D2saMFyS5dv6+K+oEVY2ttPEi+THnhqGQUI/SREYshgcxijiy8rd7F
c+5gSdD8LcijhY2OT1fIoUezJ64ZSPXDC7RAek366D/cNLrMpL5yWNDXIZJ0SEResUnoGnPWYium
W6/uuPpk1BI3y1d4Jj1EHj5HVntU/zMdpymm3XaRCVY5i4BtNh/BOQ8LO/JeAiz6wpz0MAm9hSP4
Ond30UvQTY4zpV0ty5rJr0CCPvhRLcue+FVibjfWHnXkbHnFuvevTD9mJ3xXmkiM4QJKchUjNDBu
TiSVssJSy8ItQMFRV3UwtFKFCkRWKLwd8WHNjzKZJYQUY3yEvhY9G1gozcj6FYIGUmiArpCZzjC9
phNr2Ga6k0TWx75vVFIRh8BXa3gIpme7qKjfq5gHrwOxNaC05HMlpGiXr8dG8WuSdFDiAqBm/eBZ
e/9G+XjxTEc4dmhRKc+fQzpJ7IMYQdsgyGHOGuj5jX9ahAcLyCkKSSOg9hGX+elIG5k1Iw6spYxt
1KwFSeVZ585qGstD6TW4xTKHiYVktxgUjLPLqBL+A7+OEB5Mygs/tBWTdhTCqQEQC09/zb0Q9XTz
J2dy06JO/hNaiZbLN72YCLDRgUbqqGjPYVAJj1fqGBHb/EMnPQPK1NY2scYhb/9kylNPI1EP2Yo5
OBSnuVWip+jFXjR0n7GFmJF1ItO5BGkY0y7XSvPfKj4z+LR7+GJlEQgME7kxxABCcY68+8IMjU9O
8HkqGEy2PJO6tQxMVw9wVq7sfUs1z5TC+h2VthEDnCCgAYOQVwr+S9+OzxNzKipFQK3I/YkxZ66U
welKXRH78Dud2l6MjcooPxFja64j5WJ2b+3gTZyLI75SpiNv88TDszRcflU0vB9uEGlS5JQR6jeF
Co7CGAxUmLNhRo/xt/YZ71DoKxJ2A0AoDDUa58jPJLcGg9Hh+rlDqwO8Gj9CPZM5bwrTJgJaabtb
o1rC7wyZTdo4wfwbUSPhQOB0DQvWaOk6dNQi6rS9XTpfgeOFbEFrS0dcaThiAmcNaaYLrN87Ounb
6hZhui4f8D+Emx1mTYBirYVpwrQpooPs+PI3DcLx3LtWkEF8yqOs4ql087neujdiGg81RiUQQbSv
6OAwvuE3mgLMPefx3zz019REzljIE5/ouSM2CGgIhrC2oquW2Ck33Fp0Hc2VnN8p3AXM7DYifNbv
5ufPZrpSIpX0dxjwqLB46e5HfGhDb3UJYhKL4V9NYVwnAOd7kySJ6+YU7HW1HJmFl4JTXuSuBt2h
SyjPWnBs+tDEnBYmZ5ZtUCqDUL+3KgiQi14j3uJylyIVqN1HBEuI7+JLxG7NzQJT2IKdiHhNHYfn
lC2RR/LW0YcK+2YvmF2i4nZP2/k9Yk+TQC/CtTLsocu+YIbTorTdO+tS2UiDSA98WiRgl56Y+ns1
5cwbrfSnOcg7WY14+mhvLoFHTt2Xj4RFtfZ6kR3oetZH7E4eOFbe/ujWrMw/rMD+omaGmXAtqHyB
xfly1WnpaFjZW08YEIleVG6WOkrew2Q1YKE/OOGYog85O12Bj9vT/iFhYQTJ3fw0Czl0QcI5VHuM
vGg/HxITC62T0THXlauGFql2PmSVO82muzIKM0AGgZhkgik73X55Mgyg5KKlS2w2hoyQXK8Cjl2d
5GcxXcstvjtOJCgKhluNw/SsevKEMAAUBgFqKiF1mDRPy7JwbJj/IwfwWL7Uw1voAY0QxmBaDZ8C
P7SpLzajGXDlWDTzarPUF8MRV2928ptaeMqu5MoLxaCoWZzvrwimrSj2ZB+F3HoItL0hsAXGrkZS
Oid4CKkDOPQcL9M/CKopJVqxDKNIyEgImHAUmbLRLKQLjseH3ew+RpSbKTA1Nd5ORfPS3ABTsrFN
J3Kp4WAOmev2mlGi+FC05PjvqqA0f+XuRYH1sja+2Bnf4f0oBTZQ5ZqAZCKkAsgJ15INQP6cvf4f
RpXOJq2kwo7iZTLbhKTJsoPO6meeA4YVM8M0t17jKFVzbS2IxUWkuIXEjbflll6BYUwYqjM+8/sj
p/43/4TI3CBgnj5zd+vi/6UmAH0CVMS6NzfUqPh7vTi1kVHE25qbDMUbs6a6IXKeN6bkLP7+QKtU
XBlpwKlx6I92ZBehGQKEpD+EffLg+LCOXU34OsJIurfcKs4uyjWwhMezp4mqC47+PqJ6NvD0TVme
vNzFzAXX0g5pxg3yKmhJcmKpVFhLo0oxf7FnyHfa/MrlRIQviqN/V6Z3T4601PdnuQ/GFWhQC9YT
bE1n5H3g+qk68lSRJPuN4Nw8+c4c9G7hItVbrnMXUhzDtTWwhUMMAZKDteFtLClUWLz4QOU4a+t5
9xsWPAMUNrBqlJD575JhfvcJ14WbwOwJr/3JutjTIqiplP2xzlCV9ajq61YM6TXz1u+cvA6viXBI
yfcyW1V+NaIQm+GOfi3yMRb3FoatN3eQg95C2576s8mhXOGPDSMRtyE1ppGISByU4YtpnsPcK6Ek
426wA5qI1VHA0zGxuYT8XXnaXcjKWp6A1mFsXfwc8cMexanhwi5n7oJLzgwdo9b8EzOZFSC4fgj6
FIG/FLnwvxn+F/an5JMoXNExLCZCoXt15xgU95kZvMaH4ppox6YdQ4/pzp8xHQyuHBxkHa+Fim6c
8NuQ7OeEdl+o/EMHiXSc9ixY6XflxuH65lyfwziWAL6RwNsjxvaHmfAhUWAjtpFpLeJw+OuhZW7H
hkSfsBGcFfTNebI2OrbjJVtPlRME1IRDfMdLj3O/KEHVjRvAowS5n1D7Sm85Zd4h4r0sNFvZoCkl
+pprQWjCnc6MVPySSSwQ9GxsKJXUAU4t73guCoAmljHdaQ5KvZumQyq6fsWdG7M2COZnjOwqDANg
o/4JYIYTurgZdVVTf67/T+CnBqISiuRUcfqKFclQwzr/ujj/HCCb7a3+i6lhhdWdXEzSBysnDPam
DwpGAlHcnsiMvXf6hUn1rrJpWzAOof6RCxDzrYG8nwdbTgS1SLTtKMrBSXpD2AA0Fo1xsdM0GzqC
pCBMXM/FdFBakWNjmidXp6MlR/10PKZacuNfGCv6rVPjGUdbJh79phXIHuFXvBHGf7tZXpcmjQjz
RBRtc4JN5cfPPpOBBQaCVcgegYT/Lt+ncth5ri5G6mC7iQZOK7WNPcad7PX3+R/hLl8JkEok5+Vf
ZFZPgc8RNf6v58QxOZb34TU1k7KQuIipM8LOdPYdq0vFWy8Bx5/S+1o8u+hfJtmgCgJqynCyuV73
/f1S+/q+wr0dYHR3Uk3I7sjscRKE73vRfM380v70rKohkNcuD+1oR0L/ZgCGRVqrikmKfQ3jOa8S
FZBIdskG9H6uaUxKbt/2rbnLs5REAZZ9qDahivpBqDmwZ+7lOwdOnr1fBXOd1qpT/l5z1OwG8rB1
PSV/7Tq1dCRRDgBU9+P7yCn3lYRjn5EJwZfN/ei0jztobLnu5dHXyxxt8ngmL508JXOz02STKshH
gWGoEaUfnSDqhhzo/zt1289mh9dMihowUPFokFy3TODeRIvKGPIQCw69cnPH+zjUoksd9gbiEp6A
iwm3uDW9wigK3wCkRLt5gaiY0wFY39gvwvNL61uoYnUu2UD/eg6qUwXZtVzm+UHSLsjD+IvBsu4Y
B9JOX7HCQJC86YivSiRtpngQE6TynTuetMEQGtfqEBL2gSU1QQ8dssDD96hFe1wh9DX7et4CWBgo
EyCGPrOCLaVd0bbCzBgrfqVbpZqrglNpFbShYo5u8pyLP9pG2dDzncafY31p6t/zqqR10mqZXuoA
c8SAcnwcQSzsqT2wioVsyGacYtTmyZFSb4dJlpALRSJA1+/qa48bxtI8KZwpPwmjwmgMVMw9QWtx
gcfac2B6ft6bb/tkMQbmXLzhRnR+54dE/lzeeQdLAsDkUcyEpRy2Dh8imQhmK35ZndIyQZCj7X3r
QSRQKA6w/yMmRv6vXVoNNV9xj4N3qwvZq3JPW5GBsekE4crdoKnlQj+ZDY7xljWWxWnUsP6RfVGc
18JdS870A+NaRQwrS9yMznN4dCsvFXWSEHQISvYA7M5JgzDd5rRN3op9o9SsTnLfGZHiJzWMjaS4
acCcdXEUGAnItwqzADISYuSGdDyhKe0lbnYty/7EmoP9hLIW7BpiHxLsjr7xOdSEUAZ6KUKizE4V
sQiS5EmHcT49cu6feCam4gXYe7KLB4MMyRhDL2nOvNmZx6Cy6orA6DUpZDi2dMffa/W4ervPso4b
ElPIna3pVD4Q+KDtJ+rOGcpKw+Es6XCE1nc33OjUt4foo70IRATMMKYH2VOiTwCbm3yRcKGQFaVn
NcwB1rashsYbUr3PiLrhr+pdc13gNoIxqq0QOYxy8aSfcjR4wc8xpm/4oki5uvArwuy4dMPgdksc
xpvUCN6t/xqqpK5WT7LaBoAVRCamWs6SiKpVXW299i6DuI0ZWR2EwPnMPbIv6pGH5oUs3j6ZP7tk
uFm3v6o6KTPfV1kR+nceqYoinC960a7QmK76uF0qAn3VWh/N2llNT8LDrne4/h49cFek0FfWgXdv
M/oA1+fxyu26F04Q3RhUL6gj7CNnlNOOpKHhPRQXnJiS3Nuk1PgfL6UacDwkYhaeySenU/qCOqFV
Imp1iGiTwuDMsY30m7xYSBK54YduTD6Z/ZDhjxrfDU5VGiRU7lOKdG69huGrqsAAaCXbnUpP8baI
DbnmXyJI2OrfQjtMkpJSIjkNiLXFTxcYZHOCIANEpOkDY6CQfTiHURP+avPuSUa+ySYSg1HYLZHb
luDn9PzGXfVn3noKK3TF8GWZTOCgQ4ubKRupvuSXN/cDhY3rGXKu1hII6PqgAJIRNjRxus4c0XVV
puLMRAay+6nCAaaA6i3/w4B/i7Myh/CnQOucNnayXb7YsHJyNw4aDIsKqRUs1p2+PjNYue9xCz2i
6gh2GXscqJWwvJuwRY9iAc3HINCwljuFcUwi5bMq77p+3RZ/RQpGPXcc5P9y81WNHEAQ7UaWEDiu
l67tmF/EAY92pXpYJ2raIEEtu0VOioNjUIH5FIuY+oxaCNb9o0/xOrsEGPU9S7kaCtjHk/LLOoCz
ehWJlQsVOv8/R1R5qPllNsXMYjp5FQmtDOOlgyEU/VM0Wbyi+UxYCq7BF2CgJ7M5LTK8ZWdv1oXu
IwziO1Czm8Dt4iKo/Pk0d3Rn8W84YVAkiwxkkrcjx9/uHgQxMg80gTU4Nuejd2nYZYO/gjEW5f5I
jAyz8fKJ/PLTbUMh4/hPbHyK6/vwtN9MrLBP57rGvKxJJ1aPiNWuWfdSoWU/VWeyYeNQy5jVyg9a
+oUjgDGVZBwTpBDfLjbNdBCgbkzQDhHypt9Lt9isfEaOzLuAd5L7lIbiMGzsuq8Ue9x8c7/1bm3V
h31Q+AkhW4GOXGOSHOwvA7seyW/aLCenrxtGZ5uecGDnOWReCe/cib0lcHwPw7ux9h5z28aaZV85
TAcoXEd0xXZl736iR5mvwSftLrjviMdombp6z16WoDb1LYVgTIsOynmGp5AuuUYAubfGGjFjdymR
UBS+nqQVOqaNorJ1BjmGvPsXXUTwPINj5hY3XQHJkafBuAgzY2n3lKQzMOB/jM3ncKjjQaw6G0bY
W6esRnWPMaLCZa3mUYC12cZOF+EfUJY99u7j4UaPI5bluhTGdwEy99pY3Fqc7G3WZJKC1b+pp/c4
ETOVD96/TnirsUQINmWkWfnBXbxLTZyficSOnMI8VDV3Ye06UmtFK4cHu40N+KttPfmkRd8f6DHK
YRmpGzhYVPYRZOnGAlMIbeHOENH1uUC1J+lFHZC+VGOZ1oSwmEoKkOozoDtLQWEPfFF5EW5nMOOg
D0PEQlXNQ2PUHxQGJ4nDrmWhnyCR9XBfuFvRSAk31uFinGsPfauEszfu4S22UhOVglf4xZTIWmOe
xgdzAMj6B3mLsEsRxGtdevWc7/Ps72R0+a5d1DruPriqK2sDX/lVuUBH/g8LMTTAkGsiOi4qhB/c
/11ffzytTVHX5IQNC6NfMCfPO1cPAF4M7QFlXGhWgZ93GkMu1HoCSG4Ux1mUZWDtwI8coqs8JNJG
2eIIbJRF+T45Q0LXY521m0rPbwoJ3pBKdyDVzXCeyBElyZ89wUNQyPRxPH+MXvv7AZhCVTXoJ+zQ
JbuTs7kii4luNfvVx2fJIFeaSSUdEB37t96uf/1h9eY49Plm0UfJ4oyvZoYVxVrqDF8PiTd00OtH
yCZ8mwuBWO7t7QWMeNikIoxE7TqFCI9jaJ6bshgOII69cT4VMc3DCmCqBkXizH1T9OV18mhO8CED
ZBdgPU1F7VvvHnPxMGyz7YR6WE5eZ/XFNkJDYUAwW7W9FLPMbp68HifhD+A0bF3PTizRJgxLvKMT
08io/hdb0Mpq3V9ZqKj83OJLxk6WaJNB20qF/ycvZS+1/p/K3mZJZX0TngAdMkHvWwwg7WH51Z6S
DYr1AwFz6EhVndJujrmBkhzzwYhFkEOa5sW0qbv51X3pKJp3Rvk+Sml39AJrEZvh3fPLpHJi5Q5G
0X46MMf9650F+lttUJuygItJ8Cc//1qIyfHlppG+yvX+oYTGm0YHPniov9kmKKYAKKMMyw4CuADX
4EjV7PKfeDrEU55a8HcTHr8UqJwk6lDVIhSCI9ahT5KvVqNtqvtxHTSRFsa5daZH7Vl/r1DcRVSP
o7uJlaoJVFVoXtowwlYedCeZDccCTNiww4MbTKP8w7wtywnO6J7aYgnkGzj9SUq6/f5lcnWqdl62
8HTLhxbLJuW/cYL6u5jNFpoPxiTk2Re/lJ5eY/XVShduuFRHi6zSs245JGYlLbiS2HmyvpAKhD5M
ZqhxsGbo4Mfk5NllQEcRerwH/Jwff3fya9wkAym/7MwYs9lbGX2RMlTVEqTtZodHnrA4rZS8Zc/p
9XgRl6JyjFSgNQaj8j9aSEb9eXe5IXnWr4+hrsTF8Nvytjzz8iB3egZzLcIPJMrflm2cq5sgYYeD
qceOlG0lfj1GsBDM+g2WzET+ZGrR0xK9qkpjiJUP1pJO4HtVTWWqyTVhGmRoO+Nm9kZq9/uz25FV
RBh/GBuSvcwpPtF96C9ph+oCpCD2Rbt8qua5v6t8Ye0wJYQ6Rx9MaCkNYTnFhHzDHkfuUIGYdYjM
JPkzZ8Iioe/xzI7bNq7bKjBhOIDuxnnmIoWQwvCAyd6tUAKc/4781BKVxAk9EAQmY6euHUotqUkn
ddhRGdtPsEu9YRqYlxZeGx0SFGKY+AgAivgq6kClGTQgzsUgU6BgaFqcM5qdQSbKZnjrGkR2rC10
aFHhIpUWRe85yrCv7ek2FqkGh+IiX0TVIDQR2p81UMWAPuqrpz4qVfVFKvh5hIj+DinFNow6aiB5
pVUWTtCy5ckB2nxZ5Ssnh6lqB/0nM/og2C6ebGWn8VOWIOtscI4r3Nal4yKYfIOS2KRkW+Ep2qi9
W7d+GTYJmkgiy91He/w5KfQRkLJZsKm38fwZpCPjsrN340xLPwmfWw9L4XmB1OIh1PWJSRjjOcyW
QA9MSCXO4QR8SNKas1lHhruRBAR1wV2d4r/i4IwCdBrN1WKHu4LEpyEnjB9AJlBj3JR3Qs1oqnCe
Ev8JW0w2cPk10tBVa7iiZpDNsH5jTSOUh/n50/5I+4h8C9BgMihMaxp+R42G5r/C+dvDHZ3X0D6R
jc1sA1bIys7G1hjDq+G2ErtlujN5r3MPucwbFyNdAR8XJAJQhOSqhugV0CQgKiCiJ3LAdwA0AsHP
aL1YQAlc1ivF2LKxvPV1p5B5XjsDb2MKUi2J8L5zOPeGuEwpa1v3AYedAmQ7GQwqH3xnv8DRNt9N
8PLavbHbiRXhIonWEZo/CWYRATxr/LYkotx23GvjJFtKjhnzNpouqHkPd3EImQMh3r+NftEEfIIi
euFpCILTgF11O9AbOFUK1LE2NjwH+Woyp29seRmWGkncu4VUKGDY5SLBIxqK/UfzNvWP38sg04zw
VyG68QhlSr1uThXGYkA7uxsDTbH+FDw67RtH2nnT3FWfSTiD7jXFCoK+MT5VmyIQzbVjk5yHWD1q
UUT+0Lwmp4dJ2xRd3oM/J6g8uOtrXM9akSCXxJsVkPAZpYKPhzARNq2ySbTZ4DSk3EitnUW7rKdq
rDLtKt/KJBKj4BBz4Ooh4vvnMPl8+lVc5As09LPTA6cVkNqoz877vrcoWUc0A4zTU5EiOt0Ca55z
Ggzkz1SwbqsTsWqUodh6giaxr08Cgq3vz/6DcN9OH9wFw3VefmlBK2tyn7W90KUEbB2lFFTG7L/w
P4B7bnW9QHun8texcGhgoDvVXTBDKVZ4GZGR1Qx4DjDGQ0DpED6QOnFnOYpK9vmXAt3qNsQhNrXD
DoCz+4AOjwIrVTXSvfCjdYoZpai6TLsWJLnBNl27aFbyYZ12nBVXEvEScGEb3+XXleEO/4qkKHMw
26hIWLsa/SsYlIEYOoPnz4b6+zKbsoV9AsHYhUImjiXMIE3HDi6wtRpe4Fu08YfP2dYBLIFDXtuP
fcMI58CnGu/GmfoA4UksBTN39qDpS3BYlKwywBZ3QA02UNBtd6uCtVYArLd+yKb3UhOb9KrGWIPp
RCIKzRSB9osQWOC9JnpBCCDQj2Lb2LbuVHErKZbD+uooZ9Aq2Mjcnpp0ypnSiqSNuR2pMssE3D0A
MSr/jTbl7J8V/t2+hna32Ip2XooVbfkN4/W+VZ6yTCJGzB5x+2oGx3xw4n/A+EpanLYkm1gQdGmC
QcgUge4q68Rige8tFnQOH4Q/ngmRRW4cA582Nr21APSPVLDVCw/IwqrteEOm06UssyPtYKwUohYn
O3jFFkJmoDO9Z5vM4P4jcvrB0F+R5yH+oHWOJGY9sKJ2tyU/WPIntM3MHL6ZJRLBfi0AJdjERa6Y
OogwR06ZDZF+BbFIOExpjiMcXGoj6yRuMXOnbSYeQP830xeL8KYAeQOdDCqaE88h0j5rqp34WMLO
As+YpgZQXg1PfmBGvRrrPvD45MOUuHL5SuO4UQEF93vq+1w/vNUtLCW1b4sjIuJKY4vnK0iwQHmI
rOILkQZ19OOvrJPFu9YaV/wAFLMThCzVRv25feF7vG5eN3jciDB1YvQeeqLwy/Fc0lOgYkC1Vqu+
qvN15K1lrhW+SQr4q7Yv82EEOp/AE8euSI53UWUkzpmp/WRxsKanwbgBE4zahE7qsb0DsJ3Fx2LA
bEyBnrhgqb2fqN3o0qshfDQC5JpVigC5K96pp9JBjXDH2MvqwS97Cg9P0hcSHelaiJphbmA3z4Jl
ggzbqNUm97jxzzGR/8grdZwZB9xF5WuMI5NQCzy9cTLXa/YZhGpnlzgrhb9Gy32N9+y1zw2957Pu
A64tQnUuK2Qn28FyUZadSicFTtDPHS2bjCpojBlg4QL5wgO4bpj3mLluf3H+ClbwtLzpiHhhumXk
OgqR9xckz0b2AXvPsCONH42LIBtPwtM0+knnsbbiwfczy4bndePO2CYbSr5yzT0UUEVIyT/mMQUI
p3awJXKeH+JpBIrmtlQFQULKrDA0LnaDlnL2YcJnDuNbkX5pibSMQWNDRDQ/0cJzCqQipWWDQhYX
rTHVQPEHWoimlY62A4piYzaVSFIvOZLrTwgC/a3v+YP5kHpy7l1UaqtKh/2niOOAyBsL8p+wWzGv
lgmWGFOZFlriSrynHHiKViJU26L+mp9uKiIBRAP3eHSwVaVriNohj/7M+DWFNQVymUBJJDnI26po
8Tovpqgbpyj6Uu5tmzxYRNizKXtBWEWG5YHJadyp6DdvEoUDWhpYiJd9q/erhZNwxM6X5gTaOjU0
krMsrv2gQHYSkfUWR7A6pNAjXMuGHWdgdB86u/C51jmeMk17Q7vYLQZEfs2bnYPvzayBFVhSIPZl
mA3GerYtDu6cDgzONU9Vm7lv/MgYfwZb/hhxOhVAUeSZ+wOfQWg4pCod+p0ygq4aVss0e6tCeX1T
u4BfYhgYhxK5m+JOmPTiE2bKvJNGxKD+ivCBzAGsoxmcRmwafQqVSfxjuF2fiPOpJvxJMlBn2qYV
W0JnnqYe92b0XLmp2zxeZqVb5tZBihE+Mjdh+c6dqYV/+5jTgTRJn0hyF0DQMz4BJXE3YJVgysh8
2SCNuKpdtYsb8Lso2Dz5A6qv2yrFs/cFdlmaljWv8357iUu+aspGUCPfSLmnhqHeiT/eRnTKMUmy
DkdqO11XSWIP0N+Ta77ceKyULLif5vQxjscjIUngRusYZ/dAzr+qN6SDT3yBFnIG+5YRuPpxxvs/
MtgtxKg3V5f5cNYXrrYmCXm0zBmfAM+m75uDUIYeERJUl+zPBv+YNvwLIVRRLB+3p7sizzeiOUJs
QJ8YUHZlWWqS8Veb/MK9O3kjFqslBOYJWdvfOotnlEddYInvp4scFA6hfR+21PO00YZT52xsEs7N
EX8GhJzpZhzV/UDRcWwGEsWUsDj+3ozrNJtZzVegHd4SYua+ft1uNZmK/hfQLiyPLMM8zRHXgc+b
S0PZtrKZYXLmWG1XzS4LBy0WQq5FgIqH8qV5lxL9wgDAg1K/AYy1bIoh9uvTaUYE87USHGfllpNa
yPZFPslDFkrZ8wmS7Hw6IA7wp3BWTXw1aT0EnLKogbqogy7WpBloUtYYx+hJIXC1AQu+8hyVGeSi
Y/JduTWX1GjhC6s8jKfhi8Ekk+46/LwB5OiVekvwSKXjHOegB9Tm2yUmWUVk5DlUsEJ9b4ahmIza
wuLk4nVSf0hKnI6Uj/7W6VOYs7wwhlj/nV2fviOdCNqWJeegvF7UXDd0n6wliv3LOKsrKyBh0Eja
QciXl8YbegVXTUW+BT5yoENqtk620wt1ExzVoZlkn2hZuXf92Q1eMIEu8gHFLfzIMSwcTTwSHZX7
eks+kxO7qyHvK7YPSapXx5Ao8DPf/WWtEDPvTqpRf1ZKWjP5Aw33G25Hf2Pe7Xp1lbywD6yI0jQF
j8kbALm2s6MEiyLtRpl74ma+uruBS3gXUiT/YrgjhugoJ0XgIxIaM13pyMZ4aqDu9+nuqUYE0QAu
OUK+84ffDuncOPbmBO0jBLfqp5WiiyYTlbvMCKZXSnDsjBHH9wfb2OfWbjSr0dZJGVcgt4Slwhpt
Tke+UUNUD/IlZYB+x+4pGALY4NbIeZF9yu9OXdCbBG41U+JI7axZLj39NC6R6rN5fMLFKjoAFghs
l9Ih4zxcfbjP2IiA+/V8J5gUfaZzbARfC9PrBa0GjEzpD1eMr/GwM5LcQTPy53us8Ag/dgByTY0w
e6yu+7n2fK0+xFa+x4cU4bmY+rtwfaUVcrI0P2A2VzvYawizl/lVLN0ljTTuRDEQ/darnO/m2Xrg
cYzZBjHFyO37/l8EWp/bwUpx+huD4dtu8PJ7GY8EFBhAYcXYmPbEJSmCMgdTVmX0I9twsEma7mYN
hKw/yYJ6CM+d0233vGbkmQjf1P7/UF0fXNUKjykPTYKtTQmkFqoSNaBBPmhGFdvQ6MID+tLvLgEL
ryv6Pm9Gnz+fFSJxZaZb6s5TPn6dg1ZXA7M3cWTdHSfvYuqK6zQeeStDvsu2MjG5bj3Row/sZGgv
nL/gZu0mKjG7d/NqghGxIaRrK+pJaNp+H5VQ2NjcQ+ajpJ3uVrbc+omBDqDCXHzUYeeRTF8rWT9k
XEPYnzSxopgmWVuscadBEiz9yAH2x8NCK41iGXG0JJgGWqrTKpINpwmtjl0O0lHJLmeP+R+MakF7
h7Zvngnyu/6OjDUhSS3gwIttMscghbIHrk+EUdqFfqoqEHNcMk/ddW6NKEG8Czk6DR57vhEViD8c
KUA0CQp1p5zvZT3a/XwJkvP0iKN58uFpuA5kmrESiRGds0r/9J0lXzU/O/l755Gt+yWGW49HwuFN
9JiUrRx9+xXcSICPquan4B2FnIJxjiYv7WcP+0m+jjiDrNmXO3QUTue9WRv55u4nDFf+1fpYAtC7
q8P0tHlEg0tAQjTGWQZfNusFIT6p++rKPphICngp4JUj9j5lqm4V/NNLcW9iZhBzM1blMm7uO7TX
FqOInc7VfVA1wHCclvwSCuFbnQwd/czS4J4U8KWotyTN+0lJF5Qf7pHYbCa2k9viKafzMnpxdF0V
D6Kp3W4S7bE6UcFc53ovIGItDdSySa3v21/75Ls2o27VRU2P2Id3PPZPRI+j9y3FmkXztugXQYKt
LseC+iVI/cdqF9x2uTduDzPOJyHTW23NjiZVPataUTcHUNg7prYdrE6g5CApqSH7wzFsISUsxykm
hPyKbt/xkpkzm7KDA9nFl6qhr/FF9tBSNPWTW4+NWfalos4Js/Tj7OU14/e8h1tLQehEE35Ey9PO
o7fi9VEWRgwreAAUuWa5vGDTlLuBV1uWgMAIC2Qp0uDH7c7djLV19Zz4XY0tn/N1EbcoWE4A+/DK
gvWtXs4HRxRskp4hiDEi0MKRpPj+OkbYOaspiomLfq9HT5Cm8/zpoItu/mRbrd6XSu+gxY6aprvd
DGXlRCRcd3sHJ3Haf2uGA/8nE32+Gm3Ik1zj0f40J98kvDBBgNUaIucaAOuYT25ahfnshsYNHkbW
fo/gXGwPF8//lbyZYB4dFeyeBUwv7bJ9zbiZpy4u10qgwvsC2Y3DTuMZKRp3OaBHLfw1m9YQANm6
YA8xEx4OrTSClJrvU3ezP0kds251/cVKE7xmCNr8yUlq1D5SUFPZnQVe8XhqpfAjMEK0VPq6ksnM
gtK8qJM7ncVdHpWvySF2cxHwOy7j2tTujgZi4ZhAfyUMqUEXAxEbLqpPbVFxoWL6OtWZdkHOUwJT
ahX9rDi+iacCyKtNjGElqJ/0TW56mrMQmq2PVcJGheK7vcOSES4UThJxdAPvPPKn50Rh19eNenE5
HdbwzcuQbwlhpzzeTepno/UkrHXiMKrX1131kMJ37yUlfxkCXFu+HqUjSvLyLR5k/Kixf+ZTmteM
Bz/MD2g+paMAQW5sjQzCdW1CeHXyErJ3BLP5uoO6i25X2VxEnjHY41+mUNG+EN/uexmewlxQ9hyx
HtLYP8Uy/V4LQquKUa8BmA8g5NrREQBwc4IuUSA2YQXeUMZFofiilMWIdQ7rp4seVTBW7HQm7jGo
1qb+Zi2a8cXMNykxjTqiBXE+e/XvrfBQPUtqu8VfAzLRRkCoTQqmdrls4ZOz1fGqVEgJHQPHM09n
ioyyRxETI4BUsQKTBeq1hU21Ij667f1ZcmrPqSGnRYkyiqj0NeoEB1PflcIFBAjXCCr+ySzlqqiw
by538J9j6ZlYIArntKMMhp7erBdXMYe3kQoQB6h2p8F/+MG3mP5BWR1TD1B5tGGGVAZ3NarfqnwQ
rQE169W5Bo6kNktghg+Ion0tt8o2/0NexyjdxSeIJi7FW+lViQGfCp2TJ/3WfmDlIZo2sxqQGtzd
dnxuuxdDe3PTy2Ix5DR8nvi9QQS2pzH4r2Rdxs/KLkGpYbr3pgSrkFZSQRLgg7AyAJidWAXp4ETs
Paf4U3qgKI6Aj6/SPQLzHjFYO6NOv1ohKeNFboqJKSXW41QOm1xiqXw/fVso2QfAOVjv2QrDylaC
HYdfOaVAIioXgoSgp1N+qfLBgy2GO4X0gg7fNg4rAWpOMVBcUr1sFFrCwQacCylDtupQJ4zZcxyX
ehetVP2suuZ13arI3Asift6ZiSVhTCk7KEjUCrR9hCEJldXtIC743qyu7BvsVpVlmEpenE09SnYd
FD4SAiqoyJ+uCspxlKOIkSNOZCC0h6IeKWhXzhMUfl1VLIDa8HrbtPRXsOZl1ciVsg1i/6RIs+Aa
eTi6GYV4od8/bM0/wztEOvIepDOxz1Rx2mqAxU+B9vPx8NZs9pbLkAXixgpx29DUi+ZPdaqGcOMy
JaoYVcWc4l6bs54KQtsJ+4jYvYSTzu6NXDCVR3DfvdteS4wodHVly8TPvdCCOB07/7LG00cehgC4
DYAU6C+SdNl/qjXNDSJX9ppDiZ0jP9GfmxFN7JldYNX2XGA+la9+T3VnsV1Ua/9dcV3naa9eH9aG
e34NSCwigp4aQ8urQQse0Y+L0759H8ZZif973mPViswXQU1mOlpRDQitTAA4yYi9oGB2wnsHHHq9
P4Fug5k0pIDYsVG63qrtQ4hRCugikCU1Im15eeGD89MdUyB/b+Z0JHnkJd3f+mfLvbXVWKo0w2TY
U4WrBEN8B0Oo1K7V5ayR3EBuWcdoPMo4+DiM8JRRVNOyve5oRrA6cACh8zywUB+aa7K7l2DH0F5z
vX/JP5zRFQo9WLywIP1Fcp0U+SGZU4h0tjMC2x9/A/D+NBJYuq4FqjAk8UABbzt0yuAp1dM3/eqj
bZd5BL4tCYl3m3psCVbtHidrnppQLojrwlJHWq3t592Tue4kIHM+FQPGo/Q+eMUfzYbfFAGH5Pri
qNUUxiZRMNo/pnFONM/p1uOgEWLqWw4AJzGVKStAtJMnr+/hAsYwjj6XZd8qNaYCKVivzT74Nya/
VDqPHbSYTyUJ5sq7ayK2JSTgqYLYn765iSh0U2of9/1tseeIe3jLvsSRXgDRkn60pIfzts3fHUn+
aHZNENssnGyTA3N45xYKYfE0yRH9k1khefdoZAhFWSljNwAwZ7ib8M7wMy7YVW4pz+sr5tVGzKni
haVAIXpM3hQNDBRiQiF5JNFK+40JVmPnlBTuLdvvEaEAZIhygKsaznsjHY9KJf4eAyH30WPp5eyM
Kqmn+WBltXhx4Zk03kWsNFMyweXBL/mhoJiz60a5Vgxbzhc8oeg0uv2vzGQrza2cYMXJ6PuX4CcE
s6ZclI/uNAZs8MhGEoP0bahtcE8Sb9qVFztTM/ZOQA3EbqtIQ6JY9Bon267gGxFx9A2rj4MsyOhb
506fHs0Her27a85sNu/c5EbAADeNo6ApnfJN211ftl4DFwAHtpLSSAXhU9BP0tuzN460rLkk+4/p
HuJVv6yiriCVMFL3RPIKHutdspWQEvzEpFLPvhMCQ7njPczud4YnUF7DRQK0cLnetzWld23/E17p
hy9bD6R4xpHfKBOYR6ZABZQkQBbTxksMGnwPdq54Ksb1lRWuRpaDdIQRfqdRiYFnCtyaQBzafUjf
E/DPZc2YGqZeVLj2v3Ce/SoDdrxECiGkQ2ldqh0PGzM6FmUbkGr9tMLTWL5y+bqYPCuXTcwmcltQ
mgAV1uuNka86pWiWeil1IHcMUXubGIn/hvZgzENOwoi8Qd9QP9Ni2I/qLSeLZ5GmLuJPUyHQSgcu
l9R7HmclAdB6n4ckbmdwWK60JUmZB2RWr+xPr87Y0Npm9i5Umz/J9GBjiAbt1qYRqAcOFxxuVkfx
EtS5a5xyJO5xKrjV4iuhaojVnTXAAywIPnlG5eQp2UJtuCHjOCPvnA0RtHcN8z9xqy91bYQ7+kGM
X6+MeuTbBY/1/AE0iV6uWlazdIhY+hFiSSR8Y//6r28bE5PuwwadU3+pRqLBv4yiROUm7587FLGL
lXiS59Q6mOHTvAHyK23F9jrzFsEEjmqd2W8kVkw/1Lr+hakHk5fysuquYJL4bfHAouRKNXP3HOXf
Ajg/SzFCYLivUz/BLZ2oF+4n7JKBraYHkjk7JzfOwMaC3/2kM6bGylorpujgPWmmZY0/DpPqx6li
g7i7aD77yMeHd8o04Qc7wIlTihnTPGxbyEFFEpWtzOo6rDjwV68a/PCjXTl5VA01tqLWuQPytZSj
1kHRtO2X2h66LnbyOfce5Y+AvQfUHCG878dZUuZ5KYCGw48ZtRpiPjFNNywgMbco5QE/TLb/l1rH
OzrokpuUaqDVuLb+P+nN7Jxp+PptLRq1nNOH05P1fn1foV8auRc6ifNq9JZ7gwqsKUiOXiEnILHa
UdUFW4S9vLGiHeJbuV+WTqFHq7DjE6dQbU5ptpyjPy8MHl3m0odvaePkjEyAWvAYrVe/q7EgYNWW
7H/T6SNJIsLAATvhJFmO5hwe5nt2MwOkIIVtvV1HzbCOb80FUafp5EbaM/M/Y619REJe0/Bhy1IJ
TGBYy5NFFCSUkW1+OUlGF37mcGI5Mgw7Ryd/tK5TxBsRt/44NOmANCYix26PFCSeqzZGvdwwHm5K
KPM+uWzHpAx99WS5l9syrO0GMPZMEEdrtouaPGDLfzH2n+i3X6C389drWPZLGlZp+I6K9DRI909C
Y+Nqpd6PHhF1ltmnfv92gHbHd0K3FWTC7csU7ibaRh0LmCbV94TjayOcKALD5rt1s35AcIbUyw5k
ivVVrAUJ6z0eF9qQ6i1/Gs4woy69N5A23BqsY3yQ2c65W4p4lq+gucrH4NVA1GJjvIgFzMdtMTcb
dh5oPdEoX8pIEPZsk6BW52gNo7OorL1WWHkmAtCtSwD61OQxgJagytpqmKw1LR1I1dFnG9AGnKKD
vIVsXLjLactgOjrds6ZfNx2TvvkYVYLPOA5YqE65prDEAGoE7uiLZ7w9MrUv7T592Da+GYj0YrI0
/IXLM3C1dYsDsjeHYJu6MH32GCLF73uIgqL300uM3SMyQVleR6JJju9d5UvZxboLEWfLWSBHS6sI
y6zer6EPI7ENs9H4WLJU+YXgDMWQCHk7xQ7wT+Kt0ilrGDA74KeToofTtoaXxUXQu0d7FkGbIVws
T0eSIJR6M8JKOidbEN/0pcG6FYlnlbTGq9GxhW7FfVN12VbTYlzvUShFJeSTlceGsZZag/eAY1/I
pXqM6lzBQov3XKHMBjP2PhIHJmWjj7tz02ihNRU8TJQUCweCSmSpV/GuwDYJVl8tfp1gB5SyxmDo
beAnvo4/pMsWLkWbbbT0WC283AwPKQkO2kr0fnApCvmbaQSKWiyxcMAzVxuvWhJ8MQHtzvtPRa8r
hHueK3x0vOmxD1ybeBF+HrJVQkyZpyVXwq/TQ1u1fKyIWBc1jTmYZ8Z48gBAjzaeuQ/2kShVH/xl
/z78JpI7NHWHHl+07N92SxvpDr7bkpgib7l/ZV76Jaxjg1C9ts7GM/BceKDWaC+5yiMF02Bi+/sP
HCScjId3aYLtMhxqd4pDnqDkEN3MMWT5bJpPKs1kCF5edJWUQAnYXFBLc1E5cayGQ5VDSNTw1v3C
hG2mo5WuecLvyMN5e5duZRHScbG9M/AKsLRCt9UMO8SwWRddzte2XwZSJZ5I/cDyoT0Mw1wLVr7k
ejYpRc+6dZgkoV7gZlsFbATV5UL6FZYVuHdp5Q60Ubu9+GgOUCkn0Y69GhRhn6WI7VjW630k8YrO
471sZliKXPJ99Al+mYBPlXyDzD/dezHhc9ZjEnTLnrQu2roBkyPPzGfYqO8B1O8yyWQooS060YMS
yHICWddq9jLuEef6d9OAQUX/NYqauSeseHwA+P4HN9SjlwMWce9Twbe9xcnoKwY622uN6AXdF5WU
xKmakfY1p2DxmTM651up2kxtrDIqIww3hAoBRNARBfhQ81UnkP993iB6eSg6yD5FTnKu8CX59mBu
jkFOMDg0soUUE8cImQekOfZzfwHD97s95sdUMiDIjVhbUGqbLe0T89q0PnvIJxfi8ggo/l6s5hDF
CaiXfFbe1QhYymZDjwOJ5EEqB/TeiN/3qnrBV1zRzB69dxKs9wDuIEIQjX5TmnTf3T1BH4jlZEOr
R8bULwp2XbT7MthyG5mTSxXS0dDn1pxHhVU8vKduVilgIGSG0ZdwHDmI6vkL/8o0JPbhypGacEoW
DmjWa274Abv385fGwJ784T1iJeCDYKgY6rCHffWrwj/bQAm91wl+jv2ivMelA719JEXrAHYOVSoz
bHvlMMtQdnIoVhT6yWd+EwlUkGILeWHfSM+uLARI0fTBcn8qUvJiu2Hk7+QrmzHigGnSYm42Rb5k
QEwGhbi3W5EY4YmpxQTvWnJZJRsmXjJdfVBmaujyrEIMZLYbCXzg3sVsZtdhAec8lTCXKGXKMceS
Uc+O63wJwI4oi4x0CvT4bwlnp8DfAbo276yZgrZe2oabgugpQXDwEhpmcczr0tHf+GfUJn80K0bZ
U8d3JJEtW9+flOBYB4cDdnEw+hzi0/MNaYKlqV793jjy2NtVK0lnPdDnup8B+Z/S/fQFY8HqxC7c
8viafEThu2JoifAwiXiWwRtBYoeasSbEJOBKR/WsURG+PZ8vr5GQu1W3psOpILtArYVVRP7TCaDl
x2s7bBOPf23b9VYZDIvd5nZ5Noe3k/8zvYSYN2/KbsbjWNwy387Y+PsKap9dr5/4ryg4qYrlGESH
c3FWIY3NwNeXONyEkXjHBLajKiBzr4cfbqwkuT2h1goN5RWSssatGNROdBVlXTM60Sf+VYUKB9oq
TVk56sIVGOJWoOeL2F3EOJ+3cAQ3U7xTRtRtCwK4Ua0WA1PVGFrinUjxpQdloKoN/9QWpg5qtwbN
7OYegQuMh1FsPRdlyX+Ylb8K9gd8GzDxOlGBjJLe8gN2JLCtyfO7kFe8m3xj3Y2Ej/He/Ic66uaN
yeKDDHvKX59SawmBsw1MAxlgtSqjp3pGWP8o3ZylyAQ5NnFU3yt55OVxNEXOVjv9mhqKiU6e2b6j
EqdNfZ3i4m6tx249/EgpSNNLHDOH2I//SYCVpLfZrvMjgPg7jqVieUBaqw3gJTxJnCXXT+7vQYMs
wHOTH3djWBVmTZV+BV+nzJIvl0mFTvylpm7fO4MIkqHl4wXZE4+Y0dsQdNPiN451hGy31WbZj70i
Yglai7P3MX0sTsLZIV1Cmh/vdxgswoQDwHrrtU0kRRQKQAWH+qdMaibNh4Ofnror4maJbL1sUCed
F+rqeGqyOc0n8Y0gVtYjSLhxKWMJ0/m1nEhSKwUq8RxjfbcOAZmmWXlLn7soU7kf97sbpKeHfnc+
CDOO7A4Qb+1wdnmzhhrA52vsbuxmHgybPJfFFf8dgPdFiC7o0Yj6uIikHT1waOoL5whYmWCsX8pb
YZi6YwbiT8jOYgLteCfpFTl9LSHWnr0ZOcM56ZKhNtDEHiuJOr8XXlC/FyYYEfkz/wgJzwecMAK0
aMBu/BlSApkZsrrppdpQDSVjjKQZ4O4pEL2kUOZuymMdigQY3TDOZ+Gr4VldYwf4VvEscInE/r4W
gNQAmiNG1VRnhJLh4DSSUQ9oiSYIjqWvntWlP9OCTe9Wt+flLBHIiUNxSytlOViJ7f5JCyIxBgdo
+guyWeae2uTem/MIr+pRrg7+zDNCjeg2yuDynJ87GzZlWpzLS1gjvixnnwnicwO9no+vOvL7gp0R
bWjhkxWClGx+u0B5+pTlL9eflGNGgNih6XGpxBmHIRelGMxObcQ8B/lvKgu36XoaSD+ZFbPZw3v1
5NdYwJ/m8cs8sb0xmpcyXPO7iBOI8TRXRcJorNlbIcbXdZ2N0qKtWqli7mR0j6qsB8CJXQ2oTllk
J90CO9f/jNHWcUR+oCp2SLoff6feyi7fwTJ58qHNGhwu4qgjLCN0CF0Q0pqgqqrNyrhHDJtXf8A5
87885sZBGTk9dmmn9KIl4AX4ossURJGjhaiDdgS8G5rni9XZtKKzyHuJswxr7e6u5pZ5qtQ8ih1H
SC41gsGLWN/0jN1S4gwXK+3iop/niPIEfplU0ug0B46VY66yHNUB0r7uCh0PgK03u7emQCBnPvP0
2f1AT6nTk2JTiMQcrM2jkuR99ZC7mlWlVA/gJuTaCXMIqj2wMSqwrrsiXaQQQ8uJxA4AQ8zx/UPS
ME1Iz0HpXlVwKMvjz0ISDsWIqwImIPmbqkMR0VeqU0MIfQVS+gDBPavq+4pZS7sJLxALeyR8TKzt
DrKr2Ynh7Jno/9TwokT6+Dympou6hMxLyTSUdVPnQyJlP1Ky4dL0hHn/k4+jMYjvGAUA7PTfFzz/
b2cmpIEBE7pmmk29gpSBoQtzZsVwgoqEP3hPS+uaODgtnC8nJux2Qw9UpxnACs0O3ENS12qUCpZ0
cybLfuaD+UQA64/5KC7FPpHL19+GSUUjWjiH+usfwmSujqfAEVSt84m0KHrAwOrIETxqvP1mNSFj
nl4KR4n2/p0r30w/Vy9KTTfaylVlCwNqVRV4TEcjyUHtte9tSDkFJ0fN3bNiP4AeD57zso7ec9gd
DLZ1cCCWNIPtDtWzckBOyc7FXj0lRiFmiZ3dbqVmaLhosodiGqikQzRxPjZkJyjr1jbyft9VJej7
p/BpevD1rXz5bo08P0RNgIIxwvcz2NotLERK90Yrp68XwRgWi/IGl5789lQ9Lucc13VfwKedDn8Z
APJU6z1TRNAbBsfPx09sXLyTiN6SMDXPs/PUwaO9PYaWZTdMv3e5Ct6rvLE+AtZ3dUAKv3iQ6c7s
882bWdMJisqkMpiKlbVk1ScVzPmdkdpg8fh1nNcM+er+H/369QPhtuhgSD1k4kTQxAcnke74njvL
zvDXXzyKKQFy8KPO46piKSIdQa75ySUyY4rGZxa/2/P+7Dmo47LGgCldUKRuA7RP+o5X5a/zEdmO
HbTSHkc4uZZvpHJp4GodqvzyrUPgxqO7mHVvrjBXVWy3Gt+bKSornMp7cyCTRgqz5g4rDIvzy89U
HvVv7+AAVndLxsNhBNfJkkGNUA83H7nOPR4craUMZC0MzK81Wiul2Wqk8SaO0kimS+34YYx1WB4m
73EVbcB24G3iUNt4t6A/ADuFlVD7XuEO2ukXUC0a51kWYWfCYNPsFp5emWBn4MKbJeQw9thhbu7/
EgIjVOhCK0sx9WwTZGmd5oJlozYgpF72tF7P11i37YpEC40Qcr2kR0lcZ14j3vCP5Rwl36biWSit
bI1XIlh/wn9kR+w4ghlXFtD3sAUkaTNL6dMdcgoncxopnwrT284iq6Asx8iYoI8qlh0MDhf0VzaX
h+7v82v0TYWGrQWOEYCTJYVtSc+wlcFBfucMroQx9jdu7K5hOt3E5L3wKjNl00fnAT9OLUvo8P+p
zv/EjcTju1IAf5IR4HQaXIH0od11+xne/qBEPoyfG4rhQ1v30qCaJaHmVMwdoGLJ6YpecSyG10Pb
qZSFtNgLO7dEpAgb0YKxvSdNmTdSjVcuiE9sJSGsLdcduzUPvytNTI+6cdeTrbuzNHKgp20k/1T1
/2DVvIHBn2o34bJCeds45cdfU27TKZL4EuoD1YKLhClHWhXmg2B50pDjTr9hdfxzSqfL+XIdAyTP
ocgjm2gF+Hki+RqgxrxwRtlPSeju2UWrvYiDynyeuQDgmUcDpjukbKy0C5fnp4Y6eYelluTdcB4m
4PRSniAn16sQ3V+/oJHXf/RGQHUaXj94HqlIkaqLAJxqH8tviMo80WvSVjEX7//oClAIs+Zfxt9k
duz4w+yCQ2FkckSwk0lMA8+vwe1lpwXsKroORZBVKL2P3Gb+AzNxTWPcXNez/jmnl66y1JY6/A8G
ECeTmdrYRqO/8pKmcDoe/DA7+qDVMA5QWE7Lbh0mGZ+NP7k7nx8svOze7+QroKCXQphBMfVhTkJS
oJFo3/1uhVihS1pVcg6jnJzZtxcUekt9SXhAVGnnUXxhskkS2/Q0i/0JGdZVH8Gb87k0hLUfujn/
jUhsNoS3XhmE0llSCZK69B7Zc7MhUTH/y4pDG8JxdIfY1ZAkK6HhqXLVEkwkGhHic9NuRVECZvA2
gg+FGIDkGufUJQ7V1D6hp7uC/7RYB7THoa8AAzeDy9G9golTLk6GaNLaND9I/u75Z45LeIRskTRW
ZU0XSWVx9+NgmpqvcISOEjmNPidflPEUKGPFZkMnej3yMrxw3YKVhUIfmfjueTO1cloOsijy2pZc
q6lUCGVKhGkyPaGBHATtltaIYJvTlA9dUv/poE8lRsNu+F/VwNl5rGTQa7K7c7a/cVNFKXHKVxIz
cHjIm1/0KF+7GeUYaVyUyiPXRsUeLHo8+GcTLQfCIZzrrHX/Cr1LadG5/imjpgBacO8B8btP1TPM
SK6yeSrIL+SchiWZpZgvBjSgN7bolz4Ctd90RW/fd4pE1sKSInRUp17YjTiR7Mx+Xmipp2PI3Zh4
bJJNaXvuMN3t8OQ/p2KcusrOP4ep2Z1yJQl4IADkO2tecK7+9WhuDrJGYSQKN5XMelOJRqDee+AY
FJg3xZMmu7FEt3jOOQTY6oMUfIi1+HoiP2U9gVrnLu18VHJKw0lT0vgbRcsk8524U5ejZk/1WDmt
QWOV38UI5v3iiUYgMLFVTVUbhRIvefZr6N8qeKVHwSvqfv07PIXiPbkdivjxg+DIK8vFI7mf9fMP
mf+MossHcaDlkAFk1Pv+bnuiEsNYGOPGnTgiUIrNFSLbnoaCLGeclm69p7xmX0qGzQWG9+F3mCBC
XYWzEBGLTlhTJLnJhLqqzNFNeFR0FICvsBNqXu5mfnn74unjnrABybNQFpiX8bz+VCHL0VanZIUn
ZjZcgqEISSYvt7swYbLBSMHvdNvU7zRh26klxqUEOm1UD1v7/nWvLRDRixWchC4hr5UtSfLfCHIs
/ICiPvZ7BXAbCJQXi5y9jP+Ld2H/1/kDF5f8ylZlwsC0Z2fZcf5Vt44+GME4o5kUv+4Q3BrcPue6
dh8MxF4EMHhg2ktCMra8XBxtfIMVhswsJWbjfKMTYOkW7bqbCwr/a0dB855b8zIci+GgeanG7hqu
y9jgaqUi+XmjC9CvBto1a/7dCpBrDKf807hksj7giPCVTIO1ie6UQ/J5yRgjfQmLSEJhppQeIN3f
oMFQ5hQi5lEIOhem/lqSuUVyGzNtSdC2SxBM6LZjxHwIAatl+aGCYCdbG6Yt+QoeDgDXokMGViPv
6XzdWZr2psnViilj/19CCM2OFyECfgTlA8SjLwddPxMNMApNusJNe3jgQuoFQU78ct62yLSX253+
1UkF9PhT5kJHbLlLku283BbeY95suYYzNy4RM4R8uV/bpLSQx5Jg13WXxHXX6Q7cbiGm/TO5Hpdz
hDqrkzZeKpy+tiFbnjQB8bW8WLUDPVMNm4LdHLA64X+c4XiBVJG9xZXcJbQpLjTAswPxXiVPSZ+h
rso57zY4kG0kH9453/LSbo22l83ccQDk3czEmD0vO75TklxZAv5M7Of8aJMBL+Tb7PVivfwxMnHN
19obyKdq/yr4uRHKfaa4OnRq63JVR5v3xtVxRYYRg/kiLwXg4V4m+BNrU5KjKYUH50Rf8zVsWlrl
ubPujrlEA9eKNCdQQAwip+0zE5Q6j7a9nHEhYQP8CLMh9IejKzYufcEtqZITOgCmyk7JclPl2+U1
9pw+ETMYr7ZqaTUPA+F4W72aIBVIoGgMU1cjgbwUuD4zSjpOcWKfWaSTuV0n7gBjhif9dx7oPzRr
q5xiqftYbj6bVvSILPWe1haGZGwgq16kozEeup8hhcmK7rniX52KaM9eQFK3oBKwdX+5Mg1SWKf3
suARIqMKv2H4TPwVsyvFpQ7MTxd4n4V4/ne6RvzfoxGCX22BFELsix95kPV7E72yuZDtlpQO9VMk
Oz/2GHX88iFYcUTBsLAAjxxXdZecjlvV1FhVCOacr1kOsMZWfbNqWIr4LQi/h7EgaH0jMEG7ExN8
lXG0cCudCURFPoc+izd9v3UgNquhRvxuNOY6BNJakvsuvNgAOjrdpD6IbQoRkzH3HmYqvkrYayxX
WmVpxBkagIOpQHGL2aO9S+0sEK8EQhwiCvSIi334PMl7LFwu7D3Duv7YGdXOVJ+Sn8IVC9F4sup0
8livpUo0d1tmrQrj5HGeTgqZKSyzYrr92veORaofG7hMYjoGrzPWozsEIKvfpwrt8Vf3LXvhFdak
0QEIgRvbyFGyk/IcCkqrvfMBRBgkj8SEHx36zOUFoOKNm14lyqwfbrOFNRooJ9ZEzR0Amg2lWoPy
HoEQqOVbKQZ0Rf1e7Q9DJWOYGVyrytqR9Lcc6WApRyl871S0e/WMt5KaGdoBVQ/y0obwObzsQahF
90B/yI3aAHs9N87CLrkr5OS0NaAHkmhkMwvLDMYVNxK5yie4De4T00iZTE3K6I5qX0nUQfEH5J0H
Wp9Zkyi/PNj7KN7vWanVYHZzaD/FFpdQEou0/+4Rw4uqSIuZodc9o7iVneb+OAHEoriguEMz5nYc
zQmX9XIZElxmlqhnZasERmCt7JvIdGTAUbCHqBs4kyzRVARqcSaY3Zr2zVJzxN0EzPu3MzJJXF7v
SGa1IPOxTvLcim4zantivyjEgiD0gxt00bVXSUjDuh9IzRiRYtAz50sHbXjMVNx9vBwpDDm1WK9B
SZWl+GeqHZSwUvzQ3sfYPZ0A2hj4s65nFElj+kHr44G8Bpgi8VXXNwJbWwAuP9VO4/RBGW3OjqF3
D7PAuw0oKYgeuQwwSqsVaCF20mh9ZVL+4or6QCxX5B45JntjOgWVfN+eYI/6iQEkdW5dchDCN0sZ
pVl16MfbRC2niwWa0nd+JlubXrQZAo/CbcjmnDfjQu9X9/A6GyWuuZi9Auzfjja5AqrGoOjdO8+B
mBhzaaQNd01xNh1Q1Mxj4aHLcahx0jEBgSeBGUhOCYJqK221nagOngT/RR6gA10l32fg1jDydQSI
ZHL3IPb4iJ4lQsg++vE0UuhdyuKt9VXoYKFmsJKTsZX8uTa4bVTGLOIjJuUpgg5PFStUulY/mVb+
1RBoTBenZtYnv1BeiaABkBLZ3EtsE/CT0qN0ZuG8IgfO0+XcvXy7J3BhhSC7MUFUfcsCO33dYbmA
CbO28es9R0lH+RP6PhrO5R0xe9hD+sdLLTyP20FSCoWnkbwCKNCfuLBIYVqVro+nGDONMx7jknsM
R1ns4rfTFFhMnyI/VLRyY1Ja8gRd4EBHvJZPSG/g10xjlUcT8qgqdTi5hFubEy9Dm2WJtiq25Hdq
GEHHu/iBUzsEbIOpdsGEjOJmyhig636qzQ8F8EoMnSmpkh7d4tZkNuJsDxfKUlS+fL9QugWgzRyH
fG+eCK5k+VO9ZHhAoI8MT3SJrT2f0oBD/jeybQoeP72miBdIz1Efrzlk0FU15KFlyy/JUI73JWpX
AHasyLAJBiZx+XpLA2FbNhedm4Eu15DoEpHHeDdIp8JRdXJBHhMBqrv5VtmHLp9Kk8G8n+d+SN+1
F1BxHakc2p7nr7H0PQXLs9T2/rBJ55lVSmbvyOEfxXu58rIuXtGrPE2rnThGGSnDhePjOA7h3LSV
lxt7PybseRVPPTsFY2qubjVSMSd2S3t67Qzf35UlD8R9q+4rIyYQUoMV9gJKp8R410z3pYRCLiYR
Rwg9LF6Bdg6vzqplE4imQUTKnUbbQzvmkzRsUmEJnMfcl5+C6ziuRJhTLl64gLd4tNvtmoU3771M
L9xF2cZysdsK0mK3YMR0BU+9fV11bOlIks7XX6+3QBXykXQOia3PnK7bg11th0qlLP5QC0QGEK0t
1tD6RgAJBJpP78kov9/V0VKSbcuwGYqCBkTDlkjLMRg6Z5JwGUw0LM8yinE0wDploK+FAoX+iSUH
6fOFq/OZ6zjMRfHbT5PRERdC3Wt/yP8STN9gv8rLbfZLOGRt60D65RC3xfInWWdcODt68XTHCMBO
tpOTeiwOMZcyEeMxL2iTOOfmdHY9ByCxfwsvzYmHsOeBL/RCXdmbnJVNbkdNcPjNcDIS02qOZLIm
lMAuN4oKBUuX+h6M5PAzZ+9EXMpERR3suSLwmMJTNzMvkMf6LmvRfQQ61hQyelGJwFjhX3BKBPea
EPF/mV3ZLAWv1IlLy/qil82Q1SnIJ/IQq5mJwRwo14K0gUBcvdo7vzuPsTX+0hS7ucBMV/vmMBYc
7Rq8gZdCGsDJoM0VxGnrqzeX/H8a12n+ZkFclSGYti2NxN4TWgL00/vnKL2WRVKXEytO6vKSHpHG
niPuvFWd5zSX6f1GluCRy70sWXTzpGN1IynYOBcqpPYi/IjCJdw5+pxs67pAqjGyeqiJ0V8rIz/m
1tQlK5UsPy0ourCS7jlhjEu97FQOK3hfziohMmHFIhPAZek2Vi30ZCZVEcTNZWkLZesNEWQzhIXH
PzK96OAsZ8Z9guqUrg8t6NAIO3Xt1Obufz+kDrR7DrgkN1mWu0bGeUyJm7bwi5L0zZtpRJWAbCgL
MeFIDElPM66HURrctHKvTJwIwTHodt5PqpZECUsg4bgpS7YDUThP805s5aKPYQ8QI5rquFKL9z53
+QHlTdfQn45JSvYU1tBD2sbEEAN38eUH5XNpE+ccRuqFreE1U08evEyQWemreqU6JIHgr9yR6Cao
2kce5S0JqQ/TaDWfin6OpX8QPFvBa3lSz0zXHIrPlRGOnYP9/Dzue+TQuKJa72EvZRDN1qoJ/U//
aBAazJU6dWE6P4YdJSNz8XnyIGVqAKUCKM57o8fPE+oehn/mhuCyGZxX99dP/BqAOpDZ+P6vo1tu
PtWuMlAFRHjaJtOopinysSbc5HYB8CCaumVvgfIjX6jc8Wzpmza5dIfbBNwoAzIC8W6ILGZb+YDj
/fpYW0P2JOdNAlI45ZyAUPrguL6mvpDjzCZeyZm7gadjeS3MOAA6hbpjurrv+bIBbnFvN/Kpqic/
dnS1/BXVACHM8qxYttwO18ncf3ors9kLkRaHXZhHn0cgIi+EBG3ex57EL3TrYQdj/Jg9iFaql/p3
STymvcUEgkhZLzf+K2YWVUM7+8HkPgxtN1x4653BWKzhSy1mKUoNp4eNXc2NIdVikcyan7/Ab4+H
5uCGEQMM/SKcmLTaae3GVumNQcDAzRETgPGMcMOn0Fwh/w9mMLnJJjyF1sf0xWleIbapw7ecTTs3
DKrCSs+Wf1DDfwR7zA1biywOBEmthuOgnYaoFLBX7Jne4kKqx0to9BCWAgiJbZVyXYO0mxxKgQlJ
oipUaIbq+MkERsukRD6fzuhr7CJbL01hEx97wlw3MtyFl5MCdV1cMWAXn293HCxUMmHQj1+2LxEI
veUUHGQ6jwKMRv2/ugNAR9RSU8rlU1kLDTTTqf5/dbJ8NkedpBCN3Y6L631yvSKgKwMs6Kf2Qvg9
OxAoKM+1QYtCBB+DPIQOTQnDCowqvLItIzyYQ0BpeIsFDefE6SedqgZyGGRUKn82hSO6R9tHM/r0
bAa+6OVaHXNoyqHC9TqUyKBouEg81xvSL/mSVn51T1DwVuWvUv9TGJgNB+ZkFv7wHtPgqZb0k3vX
YZ3JE98mLypux9XPWbgEl85PANPwtvmdRmOZp/stLy9H9TwSqsMT/uR86yE1/kVe2yxLZFhx18+j
IIbrY6OlyuLXF17GD7/sNC+ZLbBun0+nATmGvRu0+sD1LQr0c95qbjTkvmk0a/+2qhfNPQ98T8zq
/jW+s6vHmpedmyRfqu7KwWFNmXLS+EXEejd6eSqYXLoqLYZne7SUNexPvyNRfvAVGdh9F22UQi2j
9k+oXT/ZZfkSDbNws3YIJ80PU14QUbm8Oaw7UHuJuxkifEL/eqnXrPkQMm9xZDdoiYBQpH92/7qX
Egt/eRGZNBlrPqw4hMm3uHw6eekavAKAMkrZOPkaqWHP6QPLduYQb5vYqXSRmrwhG9TDZ8SukTHm
r1TXN8J+GHcOlb9ZABTkN+CpizQ3JVYH7zZ53hWFdKaFXuABEWXFPSlBIu8C5xq2+bDHXRJB+Zzh
mKRA5kgY8uqOpRbatRcFZsZ9lBSzQqOW1MiqXSvTbP0viT2nvvRg7+6EumRAcihZ8XU/V/9Eg/3+
Xb4DOgE4rDGGQAehKZJODfU8VS6p9fTyC80PByZDsLcvojWgpQbSsXbeuwKKCLFMs48b/SnZkQJ7
YTaryvbnLHyZyhoeTZaaUdfpksV3kucvSkDPuqwdHrp9IvkSVeiMCVh7XXiDZ/on0rrdqa7EEZxI
3u+dYsIIdrK22dw2kRDMcOL1ULgLfQYAmoOS/W5uTBGU1McVRI5JH22KYtdeKVHjDvUoUi9GgaGH
hqP8gjpEwgK47wVdQPYg7n+snGQFyW0+qpFZWbXC+AaFb33QDtpxQ31jOTB+6nD6ZkTty7EBy5vk
OMPseSod59lRBrsXi5o2xlJJiyQVVPpleYt6JRZ8euOA+oIhyhJyBXyhz4csFWoN2L1MG9bLMSTD
Z0hQYdu51Y99WBdHr2WPUeSGh0Zvh0zluRFwXngyHxgduVsgBansu+PQE1ui0p8cieMxmYZvv3Qj
VMseLMoJ+qirroGxs/XBSvINe4Gngcw7sX74cdA/8Yfm0c3F/ewhM8a4eVcAINdSYZTHxD6XrKla
y1XvTPgaPvrLWI7RB5o+q3yb3XzilG3CyNUs8t2a7TQb1sNJmUWelb4gfM0yYtDY+6gV5FY2IPcs
hRYr3r2D7BH9qSJ6rwcqzucMNzm9fByku6Di8K4HT4s1kRjTV+MDICj4kK4HwNIAXEQQAs8RSf97
XCOGTKVrlQDBm52szXDmzlMx29iU/wBudB8z5TYT0OfMdijVHH0eDZT/IcR4QrARDS22KlVLnWyh
7z3BLT1XF3zndW9ZY4eRuZY0tShgydoNPBDcJm/6SFWp+bsPrddag+xyKPppCluCLSpS+nCd7KW4
2ywPOcvo29bwLshmiFrOnDhM5L/ZWOAC2OqsBKYzlpzqxyYXTibknQ4XJluQb14i579N9XsXio/D
w73EJAS19huK4Ue+zjZS7JEMpzBDl2SdVTOfv/PME1qxNsLs7eCps6WRQwXhuSr2cbThYiKxUEH0
gS0ZVl5h7+etUEHCtmDBwNj/Ah0r7IUepUf+0lIPzxdMKh5s7wBhFd7OkVcWHF6dNZk9DtKTcUhV
UTjhlLA6AhtRRyBuJ2S9W82LPOvmtj2ShDh9mpRJOvsulH4+D3enYHNOtqGjsrF/jWTYKalzAG6s
HkEA2ygf5CsSb52lc+wi/xTPTSl3VHTzR/NMKYekHM24l8wkPyq4ubzCzlDXHE1rxdVijTTm7ORC
ZCbHtTVFHPUZd0Iih0XDbcUupJiOczyXhRQzoP0q+uokcbO9qvyIZRdiaGwVs3AQOoC+NxAi1SBU
jEZ4itzVxnxvP1QT0kxYPmUUYMKuids5CWVeFWKPBaeXzsjX5OYZUFc2bOosSyZOAMSJk8QY9t+k
7k2f3DsjTOs3+jY2sJyrrcfbyCil44Fom47TdUjMBxUQKEu6WjlxZDoBbHoCXXrXVux1AKOe4Fcy
C+JoR2FnjRaw+kAZ/6W/UmpN+6eE17RMYwdYA9mHHOSvvqRkmwwasLYTMSnjZq9cvCdXEijTrxRc
5igJXc6FZ14eujtViTHnYLsFiQBdZf1UGfjh+KreZGSoMTN9/KbeDrF4ycpKuc8aHgcvCeGkFdDd
+tzAdKUDt0STdFOWmgwCrFVX9HMbA7wzvyCsJVIhfVdbnUqz/KTFmoE3H/Sc6To/AnUoEoDkAkTx
CggDxdLmiMAFOc6gPFrrMy1M32s+v+gndHUiUx1EI1NIS9lAkkX0zoRm/i8L2Oz7aOtp+AhXJeXD
qBWVmcjwVeyom5o/kGcC7vdwPRtR6vWWaBn6mNKayt7t3kCReXFl+QGV1KcZEQ4TtvPouQJvQW1D
vBlsy/QIUn5vpJG8O0nz8nPgEXyG+EL0tONnVwqZtpFACqvQ3bpGRgsGRHaHyiq28IqklK0bb4pR
FDaqu4c5Tys5r+21FGpkA2GvsrMbfIR7AaVQwrB+vId3aQBa46SkBQKrSKJ1OgmgxZxJTzykAO5n
cdhIgfq61NUUE2qzG8oKq+VB+NfjwpxQ7Njwv0qp8MK5Gmq43X/i68m3QfqEWoQdyH6qybwkyXvn
Z4cUgBj3z4NAEFKPhBH574w7SYf68skIDoXtMgB5qt8J+UubRd3sZUcSNAVGlP82iCELfBeepKug
E6uBabWO9/jdMKRyyBBQUFUwvAp6obEezAjMUvzPw5brTEv+K1B9gygODSHGauefOvlFjiUamNfV
roe6NRKW29s5byzmKyUwCRBS0hi3nk5PacGbAwqzZCBHOh9lehsPMY411goJuT2Nddtgmh+ClyaK
DQxYKsL7X/8tz2BO6zRURmffM5xo+tmVH4XpsSFrh9gyy8ZjrDGF06TI8YyeC2gVA4rMEhqh+uz1
bMka5zOhCYAzp40xI0pTZcvLUz9cRiIrAclbCbm04YafdqHD+0ZDHo2B22ms41OhRthvPAZVEvFq
lWf1Y2f0PmN/PNf8rYuyEWdst+i8ek7//R67AohOoQWADNtC3nc+I+TGCMii5xZRkaBQrwrB6NNf
cGEWXqKHekW1FFZYInJfdo/84IaiyQ36sLRE3LoF/wSaq3CB9yLRhP39kGZB6No8fX2bcxRTyjaa
NADPrm5JXnKyO2lL25s7fejdtwmTYhIdlERrzgmYHF8otU9NMa1ikCtxdm3Y3qtIO3UZdiVgrRqK
NPGUb8oJgME4e8661UU2qc7kDaJDGobCRR2LjQJpuw5S79YYWt33vZvII1lPsUHeQC7n9VTYRBN4
/HkxoBk3SbOTQasSrFLDr25iaiHz7+aHkk9qhBNGR1K88jqMdRS7n0+/le7uC8moPzUC4OBCncog
wZOJMPesEaQihxJoEftMVmY80DjH5ve5FYW7Rh7L24pKqLcs59pb5GgtJ7H8XYLucM27yJCCOOJn
AsbyMuWwB359FKbVPbTXGmHEdy9lEdyLPcSg7ayAhabIr5gchmdU++LTdZTNZaHYa2/SSthQP5Sq
V4VhJxS8o+M7zLKfKwC09gUWLTPQ0RclasUKxwLyJlh8bApTm7vq3KK6R8OoKO51zlYBK3FpnmQQ
e9NJFJry1WPHd4zpTuJzLDKFMkcv8NJrSG6Bwxdn9f8VK4aJqENH0yv5vchRDUlAvI667B2/i6Ci
rhaaGAyJL3/+Xkl01JiNb55cHMlSeEVBLShPz2WMNK93IQ0QaQrA78V/gqhuRCnYxfQEEd0cTBsl
omgxbTw2QC+IQ3BscolQ2DrrJ72awEScvceALwv3sfJaoijB6qRP/aWZ+qFrCPL8dvm34fann2GR
3hq2yUlAI6Rqi7eJXgDqxcwiLWfVwqvgJKeVOU8lJerA+0xEbZh+hTUUZJA6GC/dgaQRuA5pJZVm
qXu0XW7EuAym+fv/yTU0Ru8sEbVDgljpiTk0TxLvq/b/lJoPJfDEIbcEEuPyOhvHseJhBVvHr0z0
DYn+EhLa2lS98TzbHkFMXoy9n4jemcO/vJTj8zL3zd6ZhvqR/0LlXjzISWt4gVW/q0s8s31TcXuw
wAC/Cx2km76NSM4uW27KpR77SxVjDh9IUzX6IDlSsMkE02XKhZcFAQkV3TtW3Mtau2chn1qkXiIT
NBnbA7M0R7UDKLP2YVraEqIgsuujW2fS0lT4I18rRGs3eidi5K8dRVk3hv94dkTuCxADto2Xrtst
c/oMEwh8CTfkWl1CsH+OiTSaCPnjnf+cV22HIVkfFJedhwE9zwkIBLzQkqSTtWZUgBBEkGFsVWU3
2d9r6JxXG4royJUlIeSkNi6AoHsLbSKDbEIb0he05SZPw5/+XWP1gz80rwFNAB/EfO8DGB3+q0MX
mPJ7QyqoZTdT0qWPLGMXbK4z1AKyA/Aivbl30ConY1F/8YulSH4/Qji9hFdbVJYY0R2ex8Alj3AN
yhv2yDz8rj83m0s8P4fIcObkiHMXZ3SswignS2JlgNo1vHibVNAdDgLL/COtsfkajnTBy+OGDdb+
tHUrLCDTgCWnsXnZyDWfJEu0xQWmY2vWAe1/gTQ7V/vpLXjPn3PeelsWnW82pzOiJ1rLitORO+Ia
OIrzzxq8K7Ff2+esl0HuyL6A3Y6P/hGEZUh5kSoJFzSIfZvtX7PJUzMWTE2u9GZLf1S6/sLLUMug
UZNIef9jhrVnrT24ipWdXeygfALFVBBj0UwwN9XRZq1v3xIerAdEiLg8Q3Hx8CEzG37F5YrLoZAh
j/c2k9ye71udWFlG8bfp5azW9N8yVII/pJnz+I8v8Wk6/Li6jwOJBg8TDlD19R9Ama8L+Tp8ZRKm
npdJIVS31JUEaalBaxmM8nBllEiVApzxpAIuydQFatIdqauHsxZQR2bZ14kXj9VoUIAor0t/J2zJ
p5DXnjN790Bp6mj0zDnPYfG3WDGsZywxF8S4s7OjvdHhcLVTiHi+JYS031xIUa/MhToR0GRi8kXM
4/0qte7Hi0VUxNoYih35jeTenF6ke9ET+leCcr6yD6i1R8T+imVBaPzSOFs4NHiHlg99RGSxLOEj
VICig7fG19uvvamns9RTQWebryH9eejpK6yCk/sMlDAeh3G1+gy1Lqz3+Teny1O0CGQ88jJ9xW1S
+aTxfLiHFgxpuYBBgrpt2fnJM5971TFWgSVxQzmZ7pdyExaCudldkKpr/QVXBUrxmBCqMWjPPaCe
JsCKF9MJUIkLQYpxWB3vdGFTyd6tui9PHXtMjAh99Utd0wpGi0vegv0ohwZ9OPDM9VsnIC0De74z
24jFH8UWzbixLMLCJ0ln6G6FgZFDfUGrDvHpB63DWjbi/Wic385rcOTozrTcc6bIrYOsHthKJdyv
ru0zZEFrm0RYeHZKSdOKTKfqe+gpCZ4TvvH9pkcDp3RjfJanElB/S3fGhVZeknou4iPxIV+g9MJ+
SRHGCb5iD9w+yc+nKZ4HKZmykZmFAh5YSzXbLLjUDLQDe8+2MEBHAjOZKzjygRWJbRyvFX1kN4IF
MZOGuanjLDSPiqWaqGhPqpDVmIeXZTDvYRBrzK17wqQd5dLOJ62tEFn1tjQgsaKIGUmfSLBQRVDV
Oj9f6edSMhRfhxEpysN6ThH37/mBGXgoppLOZaOuX2zbz7ez/vPngEvCqdYfuSPH3PBgCE6yeYhz
pWNfTw/FC0oBVb++TzdcvDCCGTta9YiS1hgJrzm+buiwsV1eA5wCFyyeZC3P7629zGPqDSOzBMIO
5Ob7ujt9eMKCQIyQHnpgsCNxKfu3QiMgASXZNgjtoclXK60TtSwQNtSCqXube1gaQsiDsbA+xLEp
X8STaFO/nakokQc6khUxMCAL4f6DoWCx+G9SYrQyc/pBVm7zRBtKr8p3zVQRjNOvvB59qEQDXCfW
e8fhOcS41v1CdfYNt8ifDa1Ubz4pkNkvfGzyazvNTo3EZbcSdmRmRp9mjkZbZbVQ9xibmUaIpWdR
bze7t6i2vPz8nhHszfatexW6wzk8zV+7Szk7TyXO0JIjVKh6Cypr0UnChV8a1jcncYvIZJbZC3xG
MIWroN8y6Np87ZMXWUem8m1QoANnZetd6JiFjdVxT102SmkVZqIbTYMjtkbrtMRIRewosuRmwvIU
i3TlHM/D0NRxALzREFXwnZ+F4KVgzUDRX73WwNHM3wx4VH9yZo8hM9kRC0mBFnP9oK8bCdCtXq9S
/80Kl6eVeTHJ7JOJTPodrl9dY5giUprk/KYh9cfHYsEzoRF2rnJjXdi616LtmbsZoz8yXmF9xxDt
UoF/88C5bcDDrBe/3V3yffBix+pLEohK/v0NjPAz7c1liHKZGMlDjOGGg2aangsH6kNZsjQMTYA4
ZQ8rTb0g2k2SDZWvsECU5NT2XCbVjVuWL5Nqjf/yuYg9IlNc+MJm66sYypmJyKm7vnUkxWD9DE/g
DfKy+/EVOFKmptUChyTy+Rq/0Z0nUFkMEhr4OPJUjvf4YOIis08Ac6HaafGrX9k0S4M3dAhGvUpF
5URw8KKj5FydLEKeCQN5zuY9Dq/gh9ZT5EogHrtDVAQzOOiRUhL/VUgvwLghXUYJx+I6co3IZ1F9
0OsjXWSfe0fp7WNKe6YgqcvgdAf6bCPyiwjSJ5zC/hb+At5w1KDucnPvDnZsa8+Zj9pUHVOeSdSe
DY1Ff1w0q2NunqRonsTJiWmKbrneObzgTwCL3Xk4Sq3gdsZzpUblXzg3f9uEX7JPD8gT+2vHJQKh
pUAtl8Ac6jfgEESugCEyHhk8laFITk3R0Neq/DCaO9rjPIKGk0vdUdCWxpCD38jJl/rhwDyyEt+S
ZaJW0Ml3QkCjcnzUAe+JZhyolbrjBU4NHHFB70AFz4iQeUejzLgeu4LSFCpFTR3xkFN8f0FrVjO0
mq7/VtZM7llUTNzqNcZiBGy0U07wU1laQsdZPnNdGT9UxnLXTBiWLJpYAXsF7XSBEvNbJCrqP/OI
HP4tPLw+L0AQV6ZzmaorQqbg6xY+ROc+jnM7+X3i7uZHSBMP6KI+GuUuu21PmqVWNqE61wTV3t8e
2Legw0cqfC7BeSvErfnFPiQzom/Z8CHar3co6GHxno0DpvCrNsWN2n3rT0gGPZtzlQ77jr+tXixu
2sgMa6Ch8cgbGvgeRjAQFPjlvXiMEZxTF+0bE1N7aFBZsHsn2/bnzjcKa6OtGt4igDsRXM6XCtxb
s5W8vMhRmmd8zuYivY5S0o5vTARLbFzf4EX2h8A/NElcxnhdxsIfo7rxMq7yKvp1s7OHMXQ6MpSF
y71WvI/Scxqk6EJga3UC2LUisrHwAE7dsjF6v8ZGaVrBtuA/GcaNVyfr+FRQxclLyo+/NH3XgDpN
VtWu2Vu7ACQvRVfjLw9F/vd/JSeFKQQVniJQ2BASBaSEh/bofWQfMHj6SNiaVI2au5tu7CpCc5QP
WbVlrfHzV1PJgZkxwxk5n+OEFuNOVsCaz+XnniRTspY6LPKOy4I2XI8AsPF+TVdIi1VzLAwOj7TN
h/gjuFxVpUSvuFP6EYP8veScxLdoB0kOP+714c9tDS1HgYYa/c7Ow1ZxTtCTPS2+ccUdh2U9gZTS
IRHmRMC72qPwuSNiXh4rYDthT7MM5fRzgJDMM3Jgpbwm7lN19sHF+VVu5Fai6rSvNx5C7xM28W15
teoCg7/Ep9Co7sg2ZrkunwxPv33P2OuE6m0RHt6kvoip8yx5JA3V5wdlCSSPClW9n4uqRfvFsNYP
vUAjSa4+uOgPIcigkaF8rCYGMNiBjNVxvqcn5QkmKXPFAPTaTPYREoTgeJqte7lUBexleKFkhlYG
X7loSAuO5Lopc20hqRWW3bQRB/AOZFK/nWNJ9r6z0xHeLG5Dx5ymvSAULVzqzd+N4I/wF2W2qYV+
jZWWRrJ92ho3yjjZTsS6kzlmUgha+VQOczs6/biaES19e6OcN3hg2CPY0CYgWKHGH9iYTq3MA2fY
qEzpoy2DZ2Mn5y1tr6Olw3usRbfKz7zuSVn/+9yY6UCH79usgLImDsnpEao/3gbBlQTxqeqrcL0I
qNGfzZtN+8WPp0akAk9MRGgVgB7gkNI7IL4Bx2qr81AhuVNZ/AKp1gIKLccG6WeKVikvyZsNVjH3
3gfMizdZl86LyfzK3YffcpTGxyoxShD+beIW39JzfZCvMHRWfyvmaVB8MI3AgBf3iCyMiWa1a6s7
M8wcZkjzUkF/LXprA5QCgnGLnWPtFhafFO4MNuyC3k3Bn3zqfZ4+plywsWlRykTWcRyJMa45WMle
uZ9xLQBzVLaC86/fBZZLUWJI8/jJcY8Em1cBlpSj2XtvZvR6X2EPD2ciPrf1LFE1t5bxxHsr+YEq
xgpO83/8mW0KXd25EXvLP8sWqL1rgLlJqdwNBggQqxsyPGPlV9YZlRP/VZKQaBvtkavPPSZNXlA9
9aAuc48zUTzFKk+Zz3wo1FRWFoDs/s3zW7rk7wXPc2auak8FZ4yDY0+M+RESuVedUA/LCfTzV2ex
wtB1H6OOQkxXgd7LlbkWmzS4meXL57djwrp46eZjKhsrA5EdK3s4wefdF/kDElhlsK/Sw7pwekxg
w7ShDzTxknkqiweHn47CX7hi1QVRmWSw/rt8Hk6aUU0OzAZvRylJT6OcXEL2Dky0sSISSAjuIoWk
gxKMKLdJbIvn9Y0aTiPZ6mvuNMTXzOSog67FLz+iXFIcLP1+J0dZ9LvzCPv7gYgmzAcpxhdYdGTn
6OPvpe4SFw8wqBNwDu+1FMV1ik1p6vCxS/G+ZalszRjNjbBMci/dHEVJuBfc7NSxeKjBAsmkd1cy
oHpT1r77jWxmtx/EuTOtXXJ1wBzmpelO9wn3z6aA37o2rSxKSEm7vF9g334z3hdI/hcknG50Fm2A
w9EXAple43+2BhJgVe938pCXq3m7KXzYO1zOrTOKiZBRaVlLHUzlMEk42eSYBcrIcotmvBeUxbdb
lYS7K9opoIX06ZBeEI4u0t6+OLGvyruInaNow1N7CNKd9SIBn3BdfkxiOJGHKU+IkT533Yu27VKG
YevjmosU1n0tsTtch+1DfvYe20SRDy89B+uVwpSlxPV+zUIuIoohPf35scfMEemg4ktDhKXFIMz/
PTKiGfj2umF6jHs9fTF3XGDPHE/9fo95HBOO1u5wWLIpdJAEZaQqy04XnGRo0bOEqK6MJyqcNTpR
9IpkpCDi0Jz7NPbQIHiFlxSKdOdygpHBpTid1PQNb20599CFbc8GdQ3KbzqjjD6nnr7wRD170Ecj
LlhM4HI0KvX2HQ5nAiwlJ5shlMgSwzXRvU9WDguxgRj36/lhtTdjBSA+dwIRvvO0VYH+NQYw3m/9
MDZyM5v2wtraf88eISeTNuc7q/uOPX4PqZzSejoGYVXdnhNWNJDSfJ//T0MWD1gJiE13aNHV2n3G
QSFJOmdBAG018rXWxA3uW52Mt/QgL7dEHm2Jn3xxe5B8LZaYp2XAYLE99xdjAFASYYjl959ADynv
XlfgXxvptG8IVfwsaXmXA68VrBjedUXNj23KVtqH27ckSttCkY8HuSPmQbg0VrhyiL/kX6Ij45B3
nXGqvvNGLgtdeukU3dV/z73pUwfbRwYX5NsXaK5j3uYRNE8C+bNjwlFm6lKQeNUxAlzq0bZcfQk1
BAWNKGinaLuLPXroWBuMUzTxXY8vAoosrhpwznBuCY9bIvjKTjO8F8BRZTZKJGHoeZKzDGA/Myfi
ZnLQYW+6ZSfWcbrIfxknwh7sHG3Hkb+Qg4Xk0ihinZ9zeJZYOEzIJrUvwJuII06q5iJv49qwtaFT
gaQkNYXGyLI/YaODl3RbnsV57WA4jOxtjAhxHtAiOjuNmT5Yl0RazVBpxDF2A00+Kugxk6tBh6R+
SsNW1j1XIgKPkfy21RknXK6mKwXlZ1yTs6GvjKiMyLGi7tGphS0zQnOuEuE7VPln6liqA+zybKKD
2hrxniGRguGm4WE0BzjiKO9zQpWf4OJF31nf4nA5kjRZk896xRZaTl69b12jYLq3P4hdi1QKafRT
AR2DCGO87Uu3fCk8cNAZBnzSbttVBhnk4s/vJZKQvzV6TOGvaHlCyBn/wKOIEi7N0mUD8ZP6lIXa
b2Qqz07Ei4FLW2h9V/WEYzutM46Xrb18hrOgHz4X8/D67m3BH/rLQLwmzsIoHihaNEcgP+TB7LB6
SzdMkfxyGoZcX15JRv4WkGiVX5tUnaDKxG6Dzv+Pxev2LUiQCrObFXGqMcsYY+vLgAMBOnPkvXBc
WtRhob2EU4kXYIC0fB85oAKxIPjADm3ZCY+5DrWanVJWVEh7Xg0fjFlfIv0WuweM6h5cNHewbAil
uVnApK0/XWRraqGRU/6sZ1oC1RNxXxa4N4vP7crpfz3GFKF4dYIeyVKCqVfWnjZaTwVU3a24nN2p
GNZH5O386LvCXT5UwJzXPWLC711coGm9f/IyUxdd0/0GtN1rSLIAbn7XNTExAO3N0sZZNi/OZMGd
qV1yOf4xzCOe5eLyu/gzaspfOTZxCvB/dnzmunWz6KV+o3HevgY+/85YooeLquebNBQehjLCdE0o
OriX8zBhfS7c3xjkQHKJRgjJqR5j9w48+xNIwpkF6p3QZLzbONLGkmXp+JP9E/LVJ0UzDR4vKDiG
qMbCQ7ttLRR5Y5fWhIxQx3UT5sqEQXIQzpWSjm48ND1kIPy1MxGsBdp5zLBEYDcMALn1RyV07ifw
mTujOD0zzkV0yTdtATXePWg3+S26NTKSvscO+yUGa0KmW6k0lcZD91xfe5smswzXx8VZmPycsYY/
FxYE7HyN15wOZYAByr8kVPdfBRaLBjECD0J66kjzHH3A6CEY+FJ0reO5iMUYhmMgEyvrnUJCzmqz
9Ft24fj54IPedHvec/9nRHQExFbuM04j/Mxt/C1XjQZp9p6d5Yr2ZM4u9T+czKeqKk1+MNKavfBq
ja/XrvtpUCJc6BG3apLYqoaVfM0sPFsHNim8iTZ4K7/XqEI3eqMWjAoR6xfh/jMigdRZVNRbHKb1
VjxjVBYiNgYpKLIOCASZOkhNy/TdPxX/wLWQop4s1Q5I3H/5ULRYIq+9OAEbVOmEWdmrYnhMW+03
CaO2VU7BySAQuByMyrkoQhgVCwJaejLQYJ3fkDwy6kBS9UhbkZfvemGAcsu5c+Bz3N05sN0iaHcV
oA55ejgBqoU4LIQ3RoFeropDNtXcM+wPDk8WEOZrzSF1Bh2UhcvL5u6maT4ztjiamcqTzspGRDyd
ioqS66x9zYTBD7rS/iVqgJEe+hG23Phz5Yr4KPHrwPuorc0283d+tgUVvntw3bSWddTUToKDyrjx
95cg3KIGCulth0Bf5ImY6tvfIktuSvCbTgPasb7LeF402c5Qmru7YP1vGjayV4r2BSjzQmuOhLmL
xBZhKBUp3TR5wd92rkwKRPprAShy1g6aDQ84gnXg78XI+reCpsAR1KczCaWOKnE3zdprHbhLjg2F
riTTrgPr6t3YEovxio2Oeznfg2hS3q2lYF9mTygMd8+C59/4r3aCE1a6H7bolf1/nFwZIb1rjRYN
2uf6XcQCKpbNsKcC88qzt9YrmhvonQqH4SGL4vBBo1HfTUqv25aS9xV+uo68R48OykUuznh9l56U
eS2e4kz6sIMLREwd+peXvIiAbQK0A1dPHmTUeSmAR/WF+3Gdb5ykEJL4KHAYVzavqxf3DdMQNd06
xfk/9i4yuVk/7c0F5NvHReUoMbAaPXskBpHhi/F6JZZfOhTcb7g+WBmroT89GPVH7/FBUvHA4Dri
wJL3ujWvDvw4l8TkWOYAdAOXX8VJasC/vGBlYnbJG5ZhM4u4eh7XkjvsYvM0z1dBsbptey91Wg1k
QOSeo7otMHkgOUbo9yk0Q7U5v7H+H0MdK/aQXKo95QAu3GlhYX6pEsXK4w2AR2sLgKFqaxYbD4sE
VMfW79DZGX314vnQW3uCV9X8V8Q4+zYER5FV3U3U8uTx32+u6F74Tk2byw5zZ8234ojwsIHEGAYk
F6v3l7gB9v1sCveEamo0Sgpa4IcQumhfcfZrmvBSatZaSBUxagUdP6ZaXaLhxc13OjF5c1AX6nRy
ZjgWphBoO7y5hUGiB4NyCKLU5+MI1JMN12vPGwCLIkz4nv888FGthw6Q0Y+YSqZ32k7h8HxeMh0v
QOou2ktygzT9/gBn01PhP6aTQdoqSYNfXbhA4WaOH1r5b2ql/CI/Nwg4bFm4f1e/GUXBwvXLsxRS
QkQQJc0eTCb1HRhJ4LCmDtptFdZOUwpXynwOe4YDeW0pr4qxAOHo9U4HjBpP6zJEkdIEhCE7Yoqg
CFZKZ7qKZrIf7kSXJt+Nqwt2T7EAmKlTXszbiSAoFkonbAUKOALY6q83KByCtv6yQRmAYrV11iTV
9zv2ejoh20zpMTpDrNHlZXBvNQVWc2Z6U2sF4MvYXrObTNeIDhzXVConArvDGZCNHXwbLQXVOHy1
7Kd12vNvi1r3LJq+rcF9+xP7mlV/kQiOAGImv1JKeVLjqp6ERss63lfviMyWUxNRjQ1aXHlt6+qE
4+7fTqqD32vlM6X8xFRNiUtOsTXQCyYBL+Uqpdr/ELhkqV6hlRTaFAqCehX5+aLOH4T1waBU27FY
ToMDcjk2MYBevVx4Eb0ZhwkK1aIHW6Wp/iHsBqB5zz7OiMSxlNPOtlL3S7FTl+0zloB9hPiN9uh9
1ASA391N97WMh4hRaXgQdPVpHjgwJKYFubWRjZwJyGT2khO7MIzQC3+U1gaa0aAoiLlyP2DJXWfq
LuDR05Mi5gq9SU3kQ2QQN74J1Q284vZRe/i9eN3zyT8l6vv0P75rUcuZNGstGT8QDBq6Mhz51UZT
rJ50vN3NwkyQyUsQ4eGQLpp46DJ2df25d++J4BRI6yHxwYTWphQlR5i3j0ieO9Yabix2vVU7buLp
qtev8+jJy5SBEA0wvg423D0fZvRevSAWzK+kijQ82AAfx1fOVhrK6zvwEuZToSLlV8U26xUKxkHA
xG+ZfofxX7ia8OQ9RZVRlcyKR5jwA6kqsdqJdXe6bSLEgbY8QzHQPapwCmfnNSd/rW3F1EGyMu+B
xkSFHMar4dxtJGaF3BpQx8MUemRaPuKsQGtRh8BjLlDpvNmJ2dRuEpVkQP16nCj1ok8QnMi81LCT
mTrjycYn/bmtJ6jcYwsc/yCxROgME7rAXDyH0dSG+iDiGI8LTqEra3o2grs2j8azTN2pcpjR7GgO
LJzj4yFl+ytHsCrZ7b0LAS8dYAOB9DSi3Ky6mm4zeADLi8x76d+9vsRXmQsyfVbxgrtINYzXZIeb
+8tEU9CLmaK7RDVif6YxChewHF9kzie+e5SPsn2MGvvQlk3H4uTdkSOE+TyHpCbiiznSZQVGaPk0
kZYZeiq5bgK4EHYb3Eh2p+3//ZchIZBkLfOaNzQe8Vkv2KfRUncq2sxMrFKRtFoYimp9wF/Aa5Sb
g0Nv2l9h8sUJ6jK9GnX4B02SBJ39affk5f548fdS95yzuzN/pLayYu5QpvY1jQsni5XYtbbW03jd
3TssDS92jRDlb8ZOcIavs54Xpx0N3hdPhYJIE54aGtz3Rc4GAJ+2stymby0LAIURtGWwSos4Ry2t
5q20UAY8YVgb24r7f2KEDTFbgjGujJUbEGnrnRWUmIDcxUWk4IKAnZzpPj9hTNc0O6zREOhOM1tG
+hkzdtZ6YcPqSaX6QdNdeteqPKrjq5Uur11tehuDjf03fEaeYjoTQwiq69CiJK4PBJQtQuba8kkG
EDRhOMCY99snK0jZkTM6qBDyj5shfwuakmBY7LGIME15KXk7FR6Js90lZ9RwOE8I1tB5KulHfWOG
Q3bDc8b5oIwI+Sgw00GFseEB8LY7f8pdJ+8mwihI2Z74ih3ZZ89W9EgPgCQREmddpsnYEiR2/C0V
JHyvKH1wLaJJhwCMClQPLFl2cluvHRjZxs6OquZmyki08BIHk1+w3rWmzqBhnJiuuHrD26b6DVdJ
A7/WpZ/eF0LbE3sNKtwmxDYYXoQ3jkRp5HsKM+K8eEEK1VtNI4dQ6996y8by1jwh8Lc/xiGzUveK
PZDnS54AuNM+jAt4FXiaxH1IQUPCtyV2Msejc0+quEgLYWQIzieb+TcqLpXAwxKnlvZhxY31bwKb
3FEZXUQQbwnYp9LZPFaFtZ3lD+lzbIfY1ozUIc2EmXRVs0RisPoWuXWA3vv2oXGTwq1viXYiwi1W
rcCqJzESegxDbGhLp/Ktv5S7QhmA2RYbOI4dvqHZKaQAXxFgfEQCvJZ+l7WtAKxSPZzQ1K+Mpzsl
D8PAQ6+f/u/GXOv5OX+cGHb+N+o/o2gqiGIcAFX0mKAPFIAWl5U6eGXL87+aMo+hb6Mdm9APQ0yX
8wKhYmTuM1s2nOHw0dOs+A1vT9GPqubWNvgzLGVFijj5B3cPe7dEziMhZWHhWRizLXP58geyRdxN
sffmLfyVP6hdB8w/luvcTXgVlmZttrF7U/B+Gf0/MYmMsh9vLC1j8Y0fqXpo2bRY2CCfg8l+xTdB
n0lUb3nVPABosu/PJon3Nu0FjHhyeU0+DaKOo7pQoIePe0iI0/7am5DjIHC04NwqmvGv13sPDsgr
5z8Qm3J6zWJ4O4PwuP8cxB4VjECj5pPJmfPtNSrs4+MT0Ce75aRILn/VOE9ZJg0jse00Fo7xcV0l
KeL/rUiQjWwe9rCzvyUPdyrsPIWL1K9/8l51D7kH1Jbhp2QJTxDsMZMxPkvcn+mKdDtwIC7SbTbu
oZo9mch7ozo0j27LoIiexnRteW+6vF/YpfsZyP1S1tOF22Bdn3JbvhFFrFXqDM7dW+hYd9uascZR
0THCA3YiN3cZD6twUeYj8sovLYWYJ1VolPPIw0MlMUjjj5lVbhDgEsT2G6I2eNhvr5lfSnnKp5m1
NT4x9T9IPnQujUXVAPO6V1QsbHZMF5XROvfbOtRYdach0xyN9l9HbrzFaHxFj7QT7RmwYSGseMBG
jVY0dFGGdJ678c0Q+E1xM/PevgXdi9tBfhgNq48u3Tm9BWRimbgdCmKhwQNGuwd8a8iijYkiOlnE
z18Y9z1M4ftdEkiVGHqHmuSiKoJ4H/SdD8sJ0ERbt68EouvbcUgv05Ksa2PHYVI/mGGjkPZaHDDA
crjePhZd+5KjA1ymfV+LCLIih9XcKYMbj3XeThN5E/ECM5RlEM4avLiIEntci6aOo++q06OcXPJC
d3S3UV8hdKhXwczcHMwv/9s2dDjF7G226edPiQRs68vRQRnz32k18v9TMXOjx+qg1l9uRWBk6xit
XjfnnU5R/0JeTKbDIAGifa16rIx8DV7+hsFc4HXlPUIVe8I/o9PAIytYwpqUIAxNXucRsdSJBX2Q
0CeTTgiNLO2WIQn7xNZ7fF3Z4k5XbFS2N8vJ0qPJPGK2M3iIEI3b7BVZP+MsMEbUWBk4aXGLKmQH
0y6Rq6+Ew5qvKKXb1XG0NoAFKngB/OZJ1rOYeKkmXw4gBm/+uexfduceb5TMafLF6JhhDVUfvwLl
NyNkH7V5RNLSz7btJm8yN566VQW9ACKfS5SCk+k+UJowNMNwecPEy7FrGnuOQ8wXZPkjcNW/d0dE
RcLt26D2bNPdXcjTiykDbuAbBNgt7oUsoQh3/2BSRBnbg4021AajjSSkGkLqhSaH+gB+UGuCVrTE
hEfbkzzlxZNOPY3BsWKvU1CnY73jAJ4E2h67Zf5CwwncGz2v21kdGdA63KBcHZyT0tZZfBB2xXkS
PifAYUBCXJF/nEwXkrKpPcmE9B8jDmUcSNvghdDwcDJC1ignF8qc9bgLObUprmK6vNyrCZa+KAhl
YSmQx4Jk1ap5l8k9qvUhBT4fbHndFLlhj0fjmDFmwsyGDNFtOq//Say/zNH4/b2zMyMw2RpChKbO
YNc7GWhZVkWxfLT6l3DLyEVGqf8alHRUYriyoTxr9/HEBQrY7PD5iNNyTeoNveNyod1rBMYbHVtH
fY/iJ8Nmb+pOeWjacElNa3uAsDSOAmo5N8IScjrI7z/rB2UlgWs6naI25Mh5JAqLw8Vuu+fXJ22Z
QZAjDvHK5pQc8m6TH6PQeRL6DOWkfp0rK7mtnkWtA7XKPP6U9xrD46Ccp+LwUGzFTQn9t4wRsXNO
C8FXYR2tPsOvOFcDI2lBv8k9RSU6wdfrfUE0fBSLATetTWtO4YR7f/Rue0rpBqjESphOjdu+J2JN
1kFjdpAW7QgPmv/s5UaMiAwIShWwuYsocRDP5goXuavT/HFyVXArqVeaaht7xyxyyYitqb7PfTQP
ENfGcWbTGHtLAhjZ2556IRLMscO3T5ZPBngAjX9EyZrl8BbSBdIJd9dz7bSFgYlNsGQNJHo14RvE
Xfmru/Xj6KiHf8Wq0aBg4ph6UNo6NT13z3uy3zhHrXCxNEaTOVRseeX9KTLe37CKsrmez02z5whm
9qth9uM5M3PjLRyQiosUZoAKPDXXlJF4G1aNrj7hm8pPzKevJpqLy5Uca5WXUcMRtUfC0vlRPcxm
eWXbEE5Whj8o8axiSBogblaWNSKyIw4P7v3Q3EAJSd7o9pcEp2tWc+NiHHbXzTFQH310hwzi/19k
zIj1jR0Dz/54Za7LC2wgWUH0MlqYdda7ai8S0KbtcsSAqAvD3rtfYNuBpoQG2XUaz+6EmididlPF
8X9yuCqK7/hVWeR2Z6Pjw2f/7+MOfjincNvlreZLVftaJZpoGS4xWlgCPJ5GxjBTZgwGmhwveiWP
DpYJXd34S1w/LSJUaG7aJshxn2PEDgbHf+yajXRXqh+jr5/VC7oGHsOVDdtGsXnhPKRRAgBP+3qy
OSI5tZeGO65RaR1/JkFQIWI9sqMYHi21mjaF6ERWNjgk3Vub/LpsNA7jhLhN7ErpAjrTgzrw7Gr3
gio7ZPozJ+7a+s2UQ6/Lqh7FFsoFAkrTPnm6f+yADMLNBMb9VyOXKQqCfA0DJbp7fz+cugzWiIYV
ncfdTojpNuu6zhpwSFw1VgfG2xcJ1viiRUV2mI4HZu/UwwS3AnK+0B16KeOCQj3QSuW7jtSt8w5W
MnW2Anh4EpqcFVrfQHwurUr9fP7pbNB4WCXC/J3qZt5WtYIfciKV32pEJHwji3DRM5XwTdMDLTBC
RCwg5KAGEkfE7dn5Fgub/9mdNpXAh9ekWH7820iUUbHyoTXSnS+Ix3KZaKL2IwvFdQRRfX+pkmoJ
z4DWom/0RJQNTg63rUdIrW0l2CY7hydSJ/9phv4dj4I5uOgcEh6ii1qz+eT6G7qd3ri/TDvJ1fZC
cLvPiqltIl0sXshy56V/LyoXAUe3Z42UuPZGf7GKHbmUs5gKI2di1vnLvBayx3wG9IjZORX2jdhf
yOQkGBgsMOE4GcVI1pRspC5sBN3JKzEoEMM6FsUGuGiduagofh5+eAWpuedEN/QYjqVyZMh4gI1M
iIk0YIG/gFORvr1EtIhDgak3AEU1nPbJAWhQDkFjffyek/IAU6dx3zyK1n1fcRm10WeFzdsDjzuf
wEoUp38VZ11gTfIRN4KTI6cbK4j18IidG9Cv7c7QXnDIbRn/4SWcT1pJEgwITEOnDxJZ/JQq3xzg
bzrWZke8FIiRMVqg+AEbcAyFtkOqrt5HZpiLrsfY7k4Ox7q0A3GsdKghhKvYd89IID4tOKxnUdg/
nEH3SYkwCzOpGxV3DOgBpr5cXoDMUqFqUuZ25WiprTfzFloEtjmDsja/74fgAd+JYGpR4sDtsDTq
X71x6VTK+vWfbF28+nF86+tFCFxCOPf/XJABP2G8lyuMYQSEoOR6WH+z6dGFocKSSq+vqkQbmlOd
7T6xTaj16nYNhzVbM668tv4/MGT6u9iQ+DLJtphEB25qpku9KjsOhoUuoC8qNQjuJm45MvDrRj8h
6QZWXaEvWKrRR5BWB4oWdPC1dqb7quW6oyCwxCl649vQvSw9IP87n0LBpd31K7iOiA1RbbYJJtwt
LcB1mG8EpYbv4RXEivAUB+7m3ZEO19vh+Pt7sfZr+Q3prKmoW1esQ1ZkMMRmxWbYbo/MBIk+Zqd5
mrn2OpVlVRmmURs846juR6sX7vQySyRwOoR0235aA3wnbH2mL4ZeYA8hdyE4Lf0R4VrqnrTrxy1/
kBm8muJKIN1qs7/9GJ4YZeONGQ4Uzq4KeE/UxTrRPVkPHdHUBIjqFYsApiyNM5aXXRVNnoJxM4QP
y36GOtX5m789jr/4Wtwx+hQr+P95pI4MklXc7LEEZt1ql9fKg/r0f33gT8vs4q5vpjvcAvuwpcbD
fgRNKhAj19sCc+9t5UllEtiYXHlLWZxTOUL/ZAhtCJyoFVDFxnt/qrfKMLeWomm+m76SNN/zcdl3
S20zFmu4y0nGAQ12MJxF8fJuNZga/nRBfGsiYc7baX/tcXEOhT7eWW+ZclSa62GQvUymR9Vi4O4X
wk42HXLWKYKC6DgqXZe522sVuJPtzzTdUhcVVSoQM7OZTHw/3V7O+24shMCo31tH9LgvzTqgJ2I1
kQYnUTqGVFwe/3GLW32ipB2bY8PaMlGOVej1wEvxihrQYKy2ZM2EPWicmbIWclnRMdr03KB/92cC
lq+3CBKIgpjwTLRKfO7mFy15w2S7udENiprVs3u8W+dv1ZuZYHpzUNlTl8295A4FZ/oQAhv2OFFb
MlBMEVST/epDAG0/stq0JzoNUnJMSsnXsNIwNpS3jt8Sd8gMy56UGCkGgMbYSEOlzsu7buIyChLF
LKUekYmYUBPec0hNRhUp55fjw2s3yXUVWMquAljlSzd4w4XccgSrhQdkmCEvj387ZSuq0tlWAnCq
y0BTZQX+iuexPB6QFtRCq4z5HWB1LB7H/OeahpuNPp8X2u4nfTUIXa8aPARRQLqyZ0TGEBzvTCe1
ynJbRhsFCZNHIU/w9xDE4ENeig1qZPGcuhEE0vHxZ9pRuSuK3tjQWiqtgbyBcgFriGEeBTlWR1Ch
0YfzeT9jfqVd5x3kMZlHpw/62xVglFRJwSVSv/oFnNTWTyE0k0fEAGeNA8t1zsca1WW5SsYFr9tV
4z7mVglmshxijTm+rpbLq82PHSldLjjqsB8oGiPM+HQac979VwH+/qUagIQSrzllHqEt5bN1rGaH
pJNj74BK/HyFhS5acMwKZ1K48LqkniQEYtXcEztHOjLvYRzlA2jfsZ3kzy5VgsVcSqO4PCgfmx/T
gGHtyOTaHCTgpNaQdN0JSS+1zRpxL1ULOwHADREt98u5EqVIkE7XHDbNaie03U3XPqJBppZlN3SL
mBungwfYG7CPDisFK0whydN7HvCzs9RCCOt8+wddkccHP7NI/ARH0VXEr8Nz9lgeSb+g1gPavUxD
hWMrdj8NN42sTqCqbNbJtu6+jOyte/Y/dTWX3zy/WPrx5nPDiceye1Q2/Xz5vdxZ874ZnmtzwY2G
BBg17v+llTC4F4N0Oq9UzFAt/e8GNEvq7gM7jvBQNBFYiNjPu3ay8Ipjn+LioT5irCX446JiUF3l
ge0oUkMyFk8RzK4yVz7sA3g2sTZJb4RqcZgDeQBMsG89xi/XgDm4unvj0UT6wwB3OpPbwT6S6+mm
1B8NyHa3iclcDy+ZUlNbYm8N0J41CeuHb5/nKSf70BKu4FkhBGvmEPJ1VpE7AFNCiI2gQF1Lc6Rk
aOcsESajvickLquTbF7UMxehydyDeLvLYjaAqr5lY2kkPKyv441JpmyEGrLQxcOjqXbyy3tbV/ra
5aTh/yE9ecY0VSsT+TzHXBx1WjYoD36QJzOjriofPhciBnDbDlhfU84mgsndV59LgWJTCUdOMBhD
2wgTMCOu8JlEsINqvDGodX8McDNOXjNl/ah+A7yonSfZSGRSIWrb7qL4+BD4GRw00W3RchqerCWU
h+X7r6WguLPwELsoJvFH4NbsIDzK4ExC3kKg9U4UISqyKTvLWUbxzRPTfkGrHLpP/Vqr7cFj1mWo
rrQTnNIJMv1Z9i12+cO2ZJBk1WSAxgSJZFSHwCooASd2/PjsWVykkO4oONOmdpAiHJOw62BAF/d2
d/OFGB0RdKNzJ9ZEthQPIZCRY5Z1y4plZN9R5YZ3Vb1xNyByiTCuxO2RvYYyzUY/abNX+PKkSkTd
l2KhRhp51CaBCNauT+k552iIWnK9z/uS/yLYlVI1Kno+dF2laxVv+WotYAgLNgvVn5gFi/o07kGv
xPuuFoAXckvXlVALFftc6Oi6bAuJf4rPbQmN42IO05TTVAJuprR3oP+uDn2UmulxL50Rn45rmj5p
/nnWfHamzEnoFKqt6RG/Nk1jbxHDIYqzKX1gosxzwQCkHnpL5NqTWlXWtZkP53vNdSeKU4VGOul9
7o9inlU3q8uRCerRjZLCeSJ36C23BjX2PX6VKD8WydiRisi5MNpZuhtW2QiP1Rkv1NkOk+yprJn0
eEtx5UgkOl6jcSIsB98FX9D78TBlRgq9e4d09zUf/vro3TyFWjLanG6gtUOb0LLYH2G4HPFv8pDi
WoXoB519AKVkRm+jsfe8Mm3D624S5PonPaLFRA6NtqNIH7Ry4byrGRsEBcLIXvOPpGPB3XdgVNCd
Yi8cmOC+iA5uXOmAIqhl4p6A7WoMdvAxd8+x2tSO9a4NPVLSsoPucHGQ0cjMfM592XJBn1jcmEA6
cbvMYXp6stQtSathDL9XOK1ti3Ul7SGBKD01cXeoPQ39gn3T3jea1tml62DvwTkrxR1I5oGYTCjl
WU2equUyQbH8HFzkMncwXC8uo5h7yLnDFqviWLQM0xgcd9Q1M7x9xaN6HigEU9URvvvoJ97YMrJA
MW3vDOtSF9pHUAgei6V/pw+eG5xO+xGuZvpoqyICu0fMCZrfG/riiyx47PvYOac1Dj7EdB+g0ppF
fj9uGlnoEcT+akqMuFccmIQL6l2x2+Rsze7lX/gC4F57l3x0yKfwUJYDrPpfALcwjDOWR1wjvPiH
OTkxG055tjPB7G9/0NVSa2dKlOpUW2sK6ymTE+erwWq5v8c+1oyiSPNSrScQOPfj3ZZ84v3sfMbO
LRaagY4TBSVRpde7YE3W169z4E65TQmEXRlxMqObkYQMiAjgj+x4lDt2Wfz4d3Ml8uoGU/TqckdN
/5mMFraex18ab/od0ow8djqdyl9MTjCJkKkjf74fmPjZQPLvtgAe2t3t0IMUVVZAbW5PBfL6WVJy
Zo6n5n1LxXWeaqHmu49NVn019TRqui9W9o4fGsmHNTb/7nIgOZ/SpChCHyPYE4GIXZdc2VR1I/vA
PGJ+5DdFdgr9wRrqrtNjGIl6F8oyBB77YEvYvxDksp2o1Fm8wGZ2hRu9iceQx9Aa25OjldVFtmWB
IZHrDMB6ldwB2W3vG3HV/nDKYJFOSZS+aSME4++GMBC3ygur1jG/Kg/mXTR20YfNmq046dCvUL/Z
s3BxMsWtvt/EZShcK4GQ4CxBd8HjMHPBXjvC2HZZibap/n3+dTYop6/7ZCR/7/DM+kAypU7zYhyQ
1y6mUr+xcTF2cGkOwr5QZgSYHgiQXWbEK4jZPvJq59h1HsS9DpTngXys8uim4exxxRf9gjV3y9Tr
6XcVWk+gycyy1kj/b8W/vbNHVPV4u3QV9r+4dhFTFoOMc6u1qS+VGuXnXj3uYw8LFIe1KZSwKqk2
Av0/jRIckG3IHXO8knjPIJ+2M3QNkIq45bRzoykZdtTvpjmjLEVHqLlzglUrVjdDPyC6CYMcG7T4
6EKerFKcHZ7xk18VRXWgDtko0m0nmg+ncwIRqp3EHJe+BuKjjaMfTDOZ4a4MGRPcEyLq1BvBNSJ2
cka2OM+ZiyE65wPxa/n6rC/DSzm62UlcxTlCc0BBEIb41zjDfWLKu0hCDijgRywb4FAZxo8+WbjT
Esl7k7Q0q7TETu2IZH8DJBemjin3F385eFjeao+D+YyZ7ksyLbraSodSJ9+12k0esnOhB2/1FYTG
tKp2gTBIo+v9gcKSmu0GIiqKp1a3VmJnRDV9ZI9J3rA+63wzWu5FkmaG9BTMLDi9RTZc+9mXNBuy
zZBM0orDwrAXacMMgIVpP5OshO+nN9XSK1vWkyiwBGV0YBJTxUILnS8D3gHnvL0IEBNEx0GUOUe/
9cne1d0IR8RXJRCL9slHfoSgbIZae2uhwKDZH7j/FCPrlT0ETy/D8v56X9nfNhZ7KecVit4KB8MT
RPkDaedtrek/CzGcW6Yaix8TBVFrvCJz6+iZsUxJTmtTLw8czFOsYFBHz/H5yacajSWzGPcema/f
FdVM++YmCmkPVz6IH6Q2QEnhhR4TPMxhOoLlNQGcvNopFs5H4UQ2KdZNc7q+M4qwoAyuSJLswDyt
DXpqO58Pi5+jrO2dpaO0oL2PHJiUqvBh3l1KgUr/UlCO4Z6cn9jBs8kztbsmnIUyMIBVsq1lgnz+
KQh/Ds1/+AKxD/HmLx0dG58xDIL7HzLzeWqaEjQrSV1d1dSD4sKUxDamFC8ntCKSF9FmyLiENyaQ
vbnq/GVDqiNALlmN7SODHgj9WJPh8n1pPDO3Zd0B2AgnmZddqsyr/DFXbxO5rvOx9NBCx5CXN/V8
5xAy2lcOl3CrwRjh21mSsMhV+7jPFyuZcLXNqkanuOC5RwG25WqOa0oRaUPFTlpG7lxHPYK/b9wd
EoGa4oie40zzSQYLi+8Ct3zZ3s5NCgx8v21ahfTVF2hoSrGi49znyI2w01aBqWZqUjD6NwuUFpU6
QzqC7gz7qX7IH57F+n5Dz/eqINN+OJUmAxIHgVr5GZgKVKcLjOZAGu4b1ulqbZ9cjXVRDDhe06L9
dxh25Rz4igiWUIOxd4T7kWJK4hGDoZYii6SKmkXxzmga7agr0e/oEw72I2d7nQfcUUwThWRkXbg+
eUrgZ/Sump5mbVxHn+8CAqrH9crEX2uQGB7lZjyQS7xxe6uERXdOI161W+pqBpLDcLfbIMd8YklF
HkrXhPzHTqtso85dbGsR/kHCo/nV1LHnTtEy/URh+CTp+Y5uqphGb1bSgKGNKLkmV/exEaDdqQJR
PGfdXed4nGVZofqJKlT1ZPa3NftR0MdvdkTvRO44Le3vESVutCsK8pP6dQvRTm6b3mNxJtoeAqS/
WSYQNlPNv8L1Icos0sqgpsVIm1f16688y12CudQoVd/yBIfEzLfqJQJ8XH2T4gHLPghMcMcg9VNc
Q7y1meIb8Q7ozfLUIoxGIZht2PloH4FMNyH92VHtxmWrxa7WxC4DvtYhkz3c02wVLfmK0QMjDz8c
nu3KoR2wWAXRg7Dt9kKyURFKM7N5UjmeId6KEfcgYLVEJp1R88NKPghMfpv968WEyxBfDy8MwSmV
K3plxK6xdX5m3KPjahMfQZlcTgoyTOdxwqFBcJ1JIpE3q56DDHZMLeNsna2KaKGkDdpNpX1hnm3h
+8Irf+w/Kxp/Ubk2oGsEbjhIJxHiQhC8r7vNKiVOINX4sOwKNKAv9xELO+Th/DsI6F/R2xiVr87/
0pk3jTkrnt/CvCn2dibA4FpjnVHzzQaI8UovWADZe59OPgcEgczgLWcVjr7fA5cNqkQgJQRqxRIa
O8Lz91LdFvgVh+YFDTR0hsDU8juGSjYX31TxeYKf191eUh++kyTx0uuiBGWd5MwwMIwMZc/Xouv6
tNOmZ1+/Y3PPz+i5ZBrEnrni1Vacg61Dd2oya7jizz+TY66VnF48HAnaJw/9aUjrykWiX9Ek79Ng
SKC0vsbyMin3n7Vs0iBnJfvhgvIzTWeZuG7clP6lkugq1C8LEOGfdgYi0Xejjh+m/AEIqMl/WUoj
+SvQVi87P6VkZ/PjyENlQKtGFRt6xb9Ridpf0h2bMJtSOgEq6bfeYJNtwx7tKI53WbQ6Z3WGvX0Y
QrYB8I8lCOMoUYHTOEq+ttwt+ESvnNkYh09eiN7gwMe0+My1xbQucPhXWGl960fdPSu0dpHCsDly
KbtuKRkOMvOtiC+k3MfcBs6y9azcqOiyLAiKT7mK/WmSYtMmOqnmOdMxhCjWvlbGMqEmIKCZvIQN
gTPdW47PBgGjD7AWpjzbT1Qw36n953MZ+/6N78/NhKV2pEgN55SmXGMaRb6pLwfqsZUqCPEQ2bPC
LgXlLdgsZ7Lqu3SB093md2TxdZBD9vXAI5zMqqUpOGEO3kl4jEVyJrn3emqVc5bgdQwuZXCLvDYG
i2sgBc7v+CL3xdmVq9XWedATcgATeBTLcAzBsN61+o9FTMFstvy/8B3RTuzEdaj1etnXvftjlUWC
h0ueCN56Vun6/GPcMnHxh/55udFI4Xflh0Vbcn5XOdhmjFZuPaU5XmMH65WA97o0ITS7Y0ZdXXw0
p+Iz6GY19sxV2iL1OG+rm8aTrOL4WiQ0ZaMrwtwFvLkxT2yEtAX934XA1e3gO6CJL6v4jC48x5O9
NzfhDkYTJtnCPj9oNjFs8NsM1v6uvaE87642RCYKeUSyg4zCSu5CEv+vHC14Nhz44o83IAyR24IE
UUGscCyBNZdM6kPTFe4jq8OAZ8QPvirZi2On86mSW2W5D0v9cHtv1h/Z6ofN5d+DCOveOzgxJS79
/4OOPlK6kJafb0IBB4OT8UOLk6DjLYWz0iejDpjdOcoAR7pxUHLKAYHTUrwUNZScMq4VPodA9fNe
p+ecsFFLFD5yg2NnZzoEvva2dKBreeiZVJH8NR0FWkYTwSATtYY7gISGsQ2JHl1gX223hOj+iymU
0sKwMrXSMJDEkBuBPLiO2JKfd+NFBjmv2TLIe6oaR/a/CjJUAZOYykOypQRTS2J/IVpJEoTsi+lx
glYE5t8YTocelX1gss3zYi4bOtDDxJ5d9uIG06znYyGOXB3zfH18KXd/19Um+Rj9S9dUBQWOD1kP
XB+4o3gLLFZTbKCkkeAhCgxSl08OEJBDD81qQHsAdoJwea6xooXqPg2l/h8xOGVD0wrxf5goPEh3
V/qDW1L2PjiNO3llMfduNgM2XtPMqF6uoNAnVphNybXGddbFIA2+4vir9+LGp7f7n1waMp8DCWNx
dVrIKatd5kT5BH0YD7A2Vr2lDb6WpvFM8Hx3v/QJGgb3hcVz3G7U2YMzgiq8obPvaIyZ8/LkJFE7
4k38d7Zu5ka/TqMBWZr/vIefcPvYxGgvEEJYt4A4EXTXN22k3G0FJyIZ88RggEgGvxGzXYNrBtr6
1g+QWyyRF1zFwuHzoLY8d+nPZ6N50JE7TLkvwhFMWeXl1RBNZVn/pzzjSswZXmswU16A++f/2rF0
Jl+BZbAafeV36doq134jsCaLjOS393x5MPoJJwiczmgisGGyaKZYZdVdM6/ZpQ5k4dKzxXirZLRO
k3fqY+CGlNMeTGI3INLw2R5AMpZVGup9sTKASlo7qJznS8fhh9GqBtYz4MiCLrWDKeSBLH990QDs
/YeSMf+pmbuktD1cKNWgIqfKizPDptSGg1kPiwpOgN8z8pPSatASjvKV9i3XlZYhPmUqD4bZFGow
N/NfYDKHQqFdyaiPsbK0dhpdkr7Q1TkmkkKkLK4d+9UbTO+zqo3wU+t4D/MJadjJfLog7oxfG1cD
NjYdgc+NMHD+zJ3M/wllDHNveFV2bhsIXVp+No3axXlcRXkYzw4qwjte3KCws0K30/YG/yKqJtia
x2J/kKMOjxmIIAfl2kYsDoeyYjAC7AKpcq1zeoFuQL7D14d6R418QZFfJxs4ph+HrEsqVA0mxj0C
nfadYXEXTU7a9fuFNfD6mek4hJ7wCTjbEMWK5Il1ID54dD5LDqvtFVI4Jyca8vhNerAwIHRmP2dH
lhypabPSRQFy9sApC3LEIJEtm6w8R+bNgb2IYPU+zRPeWqlnZSaeoOKJ8LT7oyBAmoIMWO8ynLYK
HSEzw9vCvEVg5ih5RQ7my/ylVlg6hLFTUVMcpNalH8KeJOTkZcC03GjAC/ewLSf1XDV1EZDUenv+
ZnoBXQBNnBS8jo3JYByWe298iQ+l+yPBr0udrQioAgb9drmGUq2ZFdieFXfFtfJvPV9ijsNM6gOf
bFu1eOg/A4C29lrpU+9PkvdiRs67fdUjPtZzDCBqXIqkpuGws510bzcVP61n9Ceee5lAhYrQI7aW
pEgzcuJ7UGGXQ/Qf67U9u8xu6a2u6iGFtX0KT3LKrbgLflpM1o74KYSR8p4sEYDValsGMdzdQ/qV
ptGtIIGv4Ydm4vH+LRGMMoegivK+eN6kKWVCDlneY7y6qmMGxAUA8s+ZckMrXOBDvE9MQhFu4eAY
MsQ08ORuceX1fVANVzDshulB3+44Nz4cJZadBDacvPQ7gN7Co3V0fM6RD/P3hHXHqiaAeJjd6oyu
m0V09y6jxOlf5GAh96uuggUymfitawhkKCBjPKe31REUALEOvJfaV2i1ASCzXtLiDZLBMNwQqPwS
WoAaBjQFVVyyhwrP6OSE4WA7TpGM9bvrPJttr0FESxT8lc6DMFn4qbzuBfLDSxQK7+bJjHVyGXjw
PoumF3FlH45XQ7W+FS0rRMPUL/80ByTpukepJo0xSidW82z5DXaGrSfyEPGzGdFQdEcZMK7p/3VU
I4kAWaMwm1UlfSv1w7gvVZB9mVwez7gf9282f7eG72cNKuI2bWAwlkNXc+POAaGnMvPVSxBFR6NP
xLqMd2ZzoVyEyzrY6urBX7CO/RQRc9/45J1WL3WkFTtJOXV/n+OTCgDUwdfbbGDDp5KeOFGTJNtG
Qv4aAx6SixGd3GOxUl9ihzCEUn82O09JylhsIRvCOzE/jPsyemhPKFAlLV76Gq7/NR8lOwSiDQwQ
76628RZFQjqbza13c2euDREHJ3Til2Hu4q2cYA/b1jkLt48LKKpCT8vBycFwN9XCK9vXp0tw3jog
UoRShgS9G4zA9SPHs0qGuqYA/KTWrnTCc3dxE1Z/GDpJPmLnRE/Nyzn4hdSgMoWZjGZb1eCm/Jih
SBv6avGHVkmzmFPgWe2q1bSUOX2G3z9DxA0YE7sFYogfP7Y0HiM7X9X5oKcgh2J+U2wQX8SKO9SH
/u7YfP/Ba9mc7dOMuF6Xgii4Bd+hYlGpBHLmixIPb1XSKKSodfGfWvwFM7YlwJ9osxrEontxfHge
Wiz2BDW3dcqZ/1eIdSiDgwU85tI2ps7r3DRkKvkccS2pv2bGX+Xw1ZmSB233Chcybe1Z8WXDxbBq
TujJe97gKUWVy3HN3uwQqfSWCHytHsClhJ3GnSR5TPyLt6g6CoykZDUcMd3Rlg/l3cgcxe7cLnvQ
Jl5O0QA8YOljSfRzwXGnIbDEHxLgAXV4jMmChFNPXjDO0V5C9HUCOFvvRVmm2V4RBo1Z289xmxOs
dVoMsqYb8Sk1dujLIhyyuDA8ofPiXB2dNh2SCOknZDeXfJKtnnvUY8o2kxSnJt0zfGEGtFGcXC7F
nDmVc91pX4Abez+iM/NoZvFAki8rh5z9Qy7VO3fzhydgckbj9XnKoPX7QryQLYYp34BwEIKcsxqZ
sDv7Im1rUL1I320OFnwUbZwGNWp9xzIHH04os54ALMZQZMKg88IuuXV1Wg53oJIktojRsCXXDlzy
vZUBJ+eoxZ33LLpFnNoHgRdGThkz9VEW5zbMdW5EvXbQQwRBPvLfTHrnsNLySxCfBIQ1FMrBN/xA
lffsMG3L8sTDyz64XCB3HiWwGmAr8rnO1RsEuSz96HLX/QrEGKTDrP9BiyUAd08gX+lIZ8+E8mbA
MVMjdEN1YDkxWuckVVZAAdm3kcfFZfYO5ujwiPnpWD8LgkVj4iWKdD7k4jcNkCvmpkcCChiL36T5
qXdw9thBu+2G1FK5OWErR8wLXdCsKycbm/wQIuJO5fGKkcJyNK9h4octKURaC7fxai+w+LANhKfD
1qvxfm6L0uKgNwKuQsKQm8QnDTHcEjeluPt2ISCwCtt1cr3igbjDOFmFq8TtrjNbG15NRDBr8EU1
qlCOwON+dIHKUujoiTtAr7+0YVaEMXTt+zkrYLO9Ofkm8LODPyNwbNGu0Q24WWLOJwTUFx7P7n0U
R7dPyvc0UNbeX8Cyt4wv0F+e9RapBjYBNl6BZIJTXxr1dshViVJDPUuStZMD0xNL0BQFZF/ywEw0
Iv7amPq4dJo/yz9Po296Sgb2w/iCthkz68H4auM2A7Uyh9pLswFYmSzOoAQWcDMvL63dU0qFyU90
Kp1CWY2VWvwQ23xRB6nUrwoSv9yTF6f+UrfF5EIwsvbrzwBpwKyFp9THgRqq3H62w/z7Es40QJlR
oKG4k46JJ5Jv5HrfpnSCHrHylFA9enK2WS2wUKFtemMdaLAz7CZI5EM1aoTD/R9srwZGelg6t1Wj
ss15AeStSOEcEdXxZy4lzFGFZD5JFYezLHOC6u5qErvUKbemSrW65Y33TfQe3TZ+/LQld+xOylBd
6tkOfE0HZ2yk9ROeE2sv7yKG+eed4o8PQVbDm80VD9bffvtjIlpBIjcmosl6vOg5b3+DBZ8D1lH0
VdExRyyj2MuRFLsr1wUUFcYM/2mQLyqdi4a/rWlHnqKFhWMGZDm4CpUAQtMLsMRQkqUwnmGDXdSt
53Sn7BguVLjmFzh40aQzo/mpTIYKEkYn4sWri+jt+sHFdhRCkNtYvUJv3ueouzeLkDvjc2BXYzur
Zri7vSCnWTzdwf1gOSzEGDlKot2BplJx1ZQ1UnlwHIommonYWVfJb3PL6CJ8rh8cCHnpgp6FmKj8
wyh5igJ+hY45tIGdACCxbuXgZTaDEecRaX6YRzA3HflKiJA50BZPn+EdTfltf/xO9uZ+TrpfqhjT
FVgpVlv9zOLE472VLPfNXb2v8FT3sfTUN+i5eJ+uiw5ws4oq2MF0z2Ie4SQob9r119HL5urW7ZGC
2JA7KunPVtJZptlwtfwAOj7eppKCg9VlfEB/Eu4y0VRshGCDrFyggws2l5pNRycGi0DKxil5YDcJ
bJ4v8j7CFm1KXmcaouD7J8+bCqecac7T59STz2WOWu5Q6Zv8WACVASv9mnLia4mu3tPL98/bzi9v
fKAhgsV5NHHj4ASI2g3qpnZ7DsXautUpNhRBwyEKD4ovxoB0dCM15rdBRPPcawhDsJfgm97opjTH
za67qe5mPV3xse5U1TAsX7bli6MtO5sL0yx+DdGemUaNZvlkFjLL+Jqwz634x2ZSCoaKasGqiao4
T1Xx+xiTkmPwEc+zUBied9FUdpRWi3025DZlRKC2fS0cTKjJ2uoLz4J87Yyifaavdp0JAg/4t/VW
xf5FYDQuDspQE6VftS8H5GOXmE0uEzhbl4funWYd4LUUj6NDii94KKaMBeSC0DTsUvR7ujXSruh/
rZZfRx3Narg45n1jtL3zin1RkFN1V1e5QnjaEox7dVuIbBF/0ugqZDim7VzgUVjrwwXg9hULj76R
K6XddyM7Xs2IHsohMy8WS9TqkKQafz0xmd6pmDdR4NJh2U6KNNYkr+Y/+QhTW07vQi95ZiSWh3ZJ
mV2boJ5uUitnWMlib8M9bwlNTkqUazt71W9xL7deWnw8Id8Z9XjCJa9K5f4ulGfkTQWyAN+os6IN
V4s0OQh4QvdhTrp79wfUQEXBt4+PMs4J9aOI6AHZu+2u7ePXmshvdPKdqgurWpY9OI5G5Yl3fhTf
QOKoJDwaltZgtJoNuurJ9De94eR9vb+qtUBJGcIr7mwVQQE+tej2IcpLnDSnYqefJhIhFnyilc+t
b3X12wg2xsdsp3ZhcMuNi/eoLUIhaf3mHiYts56oF61AD5Cn2gzzhtPNWneqVNk5LWv59IBw2Ehn
QZv4tE68fan5MQczsA20cJf3byIkWMHGCTGBX9tZtnOI2pYlGYkuQbEBMMsYignoo7o8+foAda+t
EDNZYrMEC650uOCVb73A/xUk9uIXD4w+BS8F1UieBXxRBhuzbeVhHNdJv8ZEuxR8+GpAaVEniGi4
TLJS5/802CLjCJxXjxviKwomCpI720CRzKUXNUu6U4XYNT+E5wkhNGCaM0I6BQZ3hVGUE0RgNaxE
1KmiA9NJvC8y1T+nb1JCpMvAIXfWg3lN9CpU6Jh6tkUm7cRmHwvP7aaOKtJiMdyZmYntl9iQvOBE
a1qKioda7tY0I/YjBymBtzNYmWaLu5D7XqbKjIm0RkbZW5GCk/Nqd4vYDCeKVG1EJ2j0qo3D3r59
pt29VlhLGiGmEXFdzXHV0rwW7hiSXAB9cdp83PVvMbCyCKa1YHFYwtfJanHI0FyTSjEVEfcIWMr/
sX4U5LcfszZUt1DiwAU/viKMFmGr4TWYdQVxInaa5+loRQLfGrYt/Ie2OpG2EENF+egtSQqe1jax
0Tcz8ZPfL3AQqBEZjRZGWhpXRLhvGmu/yGSsUBxInMbLPJQyXlGf+r4+clxSuCXnozmP+boP2rPk
Cm9V6CTBOl8GG56MqxgPSiIQmk8KAbhZnAQlRBY6XLqbEXsq7G8+jNQBXV0rn7u24+EtZG5ZQ8Af
lKExiDDBCjPfolD4WMeN7MAITrsSnumBXQbpCkypjVCCS6X8dgiAcQ2aTgNllxZoRBuwue9M5N3+
XdwEAXPJ4akbPFNHucqVEClSNXAlTM1sYnPhYVhweGupyaktvGAW7m6ixx6E/OpIHCP497vLGBSy
6JZ+3RJxWHPHVfpMp6iBPyxVZNc7T+5uZpO2EFQuuXcnIod680zxHWdJKpnXUgIlphAgpOoXU+UQ
F5z87ysw+i+/F7Uq+AkOIH1kzGXe6+avWd19uF85cgr2nsG7HdxmeKkRmmjgTHGgaSB907eMdux7
NpVFi2Qr2L3ee/4YbXHFSPd0jWF82t0nMI30y7Nv9/WWLhpMzCigEYm7qGYiw6LrAWxThPIGYIvc
qyRE3UuIu1FNk8RDxtjZbsl3DAawkXzg3B9Pqi0NGRyHEtaTiwrdA2a7leaoZSYQ6G0EXqT8zlET
F68w56bcoJytl1xa5KVy/5mKcSAK/9hMttMm13UJqa2sr/zo9hLnW/1zVUH+dE8z8VE+SPhLRtO0
J2p576ib87CKKCTbckwEWzrpXqbAV3qzocesm0lz/BT5/O/M3uJmYWjBeGDEMbklOPMbITA3XcBK
40dmp45V2pc9SykxsyBFglBxqXkXYjbYcSooyN/KPoFQAc4fuEWHMfl3Vtm+eoVCOFxVW6MtDSdB
bI7uz9qKxNjl9ad8VzzUFjz0WrlPkDUgRfU8k4EQmTlxoVJeAtFQ+sNP3GSCd5KgEVNCqcCNqKRi
WuDWQmHOzB3C2BCT6yXCmWECi3ikth+Q9mQQFqDljChuSScX+htcwnWZ3o8HAFryHbMe0uTabgEJ
ONsNGWxdtesB/veIE/6c5L9SNDKZ+UlNpHjiC2sYNB5crHNz8WUlyNJKgGJPT7sEohIB9BjScOeu
bZti70Xo16A+zxyNH+/yAgYIBDG0kcNnRg9saB2hHAZGW6LWlnsiRIbfBhrvcOm64SLrY4LbKfZw
I+NIvPv+8g6KB3dfm7bi2X7P5/qTxlwSA4h7NC2Jf6woeJuns3pQq0kzNh34XB3e+l5kZvPx8o6h
mWSyah4DRp8QrZR4vMLIEO+ZNSM2idVlixbEZwVbbnDJhS0Dw0iBK44JPpkYxZNRjW+bONm1HexA
b0ywMvMUiAVnbX5AIyPWK/cGYQ3aRqFy07qypcpkfRonyLj5XH9DUHSSSMtLYHTO6G0SEhqmBOwC
xbR6+/fE23zBZOUxuwXG23q4iwTBlT8CejrZoUBaoWUJIf/6MHhzqDK0Y1LwGyNeWqwqFvn5QuyH
mQ/MeFUYhqFuSDd4MBS2GSpyr1rL8Be4GpcccWFxDoea2FDdX6q63LxlpZbjEH8SNaQ/YWhWA7VV
Lx/gL2IU4hpjGRIDX3GFlkrtYgql2CmCNYczanL3Ma3uIYoRurl7WT1UWeB6nYGiknueXLB3OJ99
Pudr1VbmtCRR49iKQeoy77q40gpmjJ/wewqY4kbNbOdMUREyL+IGm6SXx4MUzxrgMEUc37NZYMa6
5R4g3rMeB0OyGLsv6wo7ZjOQPsLVUdzJ3ssBqrPHQNGc2nP3D1KVOwzd8C9txs2V0uZ6X5z7iqJi
icIcW859EiBYvygH5LJBVgBQu0TBuRauiPGL4+ZZL/9JRsT0Tuk+rb2tIZODECXGs1krJvFnRBQX
op7KRgwGpyPveJ40qSoRqw+yJLY8RDXeFFrpNr/3U27Pddj4IzUmXDhYgwHAy/APyoXpnE+tjiQg
2ulAGatqhJmT1tvyYFzsgCgQdUztR6qJPrHtPUTuYbik65euWF61wOxibJ+cbBu5wpm4WoOeh5DM
gichHuHhFyYAOGnSoEf3C9lcBRInWScY38kdbT815qviBMJL+EZpckDwD+JXJFrUekkB9oro7idh
VCCcPHx9EjUS7S8u61O03xW2Gt1BsN6JzcAzTy6gM356VeUOJtiftCZ2IrMMcZZNZyvZUO2wN/h5
D5WfaFchaxKt6LmaKDCYSOwzQRarpiYniFyvMCxB71++C+ksUD7TxXAsCp2FeKyqs9Qc/2/wfKeo
d8ixUAmH/LU9fxXTjXBSFLWqY29YLTk3FIXGP9ZbtrTchmQvgj1jIjPK4yRgBELZsH4Uhm0wzI6E
vNHWfjEOFrF8erl/nMG8qbn+oJo907VquON4RiNMHITWGEDB76Ca2Y1r3/XPdp2zoQiv3RUvK2hw
CjJAB0wJhghV4dclWcgBZ+QSPPFHK91yx14mJ9ercjT55PrE96WEtS8r84FYklDD/C5O5UZcC1gu
fDFCuVI1dCrYb4EeNHLgfWZ2LeoV4vZ6B6dNULVb/zDun0LX5Xv1t8hSvmJkyIacgzq5IfBDlzvo
5KFH573EEv2yIdgOnZbeeL7G33FexnC+Smu/gUA2YdaNV4XbsXsneiHpyumb6bR3So2RvWv2hxes
r3UZuYpPkTwJUYS3RdjR3CCyaPO1Jpr5B8HkASGE/woz0RWpVN+GYfAMcaprY2mbTMoSEI08ZMHj
RhsOaLK1ZdoBjWZdpTavl3r3P74aHSp6wuLQZBFwoOANqLz5smxXNT8BE9BzGzTc5aVvv0w3gSuS
DXTGcKITFa2N7tbAN313lQr721Uz23duQ6RrbyDaN3tU9a+T9IHPchUz5QD84EQNP+tIi9czpA/B
t1LXSZQ7Edk60qYPzxKoQP02meHnjQluw2MPFZktpksso3EtwayskwVJ9b3Rp56aGNGtW+E5njsa
Kv1LyplVtDK4pAV3cfX/z/jWO3S6nlpoIND5wuncvpP5s4ObjA+Kcw0Ow8n/nvsMvDrmr4ZRNF8C
Fp+UgAIBlGA9eEmHgEX04ChM0nROPOkvhfhnRueizf4ichEb8ofE6s1wpE40oDoM1lswnF+/ULpI
3oOSBiAkz2BWco7+ALT2K7VHqWyKmQD9EsuIyuOFiV3hzGCGi2BmiGyCNPXnE4ZdD6TgkJumRrUe
AntvUCCvjyOqJhRcfsr5TYtMBJ9DHlAZc3fJXUdpCIEApNL+WC80W+wP5+0rHIaCP89/oOYM86Gi
iD71Utn0TdCkvWD8AsA7cIMB3K3ruy9A3BxZiOolpH4luTnMXW8gqdb8fx8O501smIZVb0UMwc1p
TREvU0S8zNypAf0XEofZloYMXxFYRb6li67GZoxduH9xfW4gZVnDOP3mLkV6iD23sdj6a1yy7WZf
DhyZ8S8L6nlUpKaj29ArPoqk098M1Z/sS5KOOsybBLJvsd+UaSbdlnDWcDRI921VOJZcueMuWim4
mFBRil+A2l2mjikPGQeSx+BC5RhZ9r4Qi6rYu73QjBJLqOLeYs/E5SNJhFc9Lc5fhrLH3y/d/8JW
Fej8R/EBlb4z0e13S4iCUy4f8BeBnMNFVmUTGFiP4inNSytAVd1b+rPZkn7yEv6cGpA5rW5BHZJZ
qVZOym2tqmZdOr5bkTQ4O1CGrdYkaPNRnB8yXYTDL2ClcNE5t/u7FW0vOdeQVHFMQvzrQ8m/yWvg
n3jqB+C5/r5AhstXACY08ruMQwamPi02iCVEu7537NFW4BcvowPZpQ30i4wJIbyknDR/cKl331+Y
iIg+WgrPNpkqSPcKw3zLAlLL5I2uGHdC5vOCcAJouJhyxHbLB6cc7L7v3dCJFQNHehSWxgCDRPE7
tpdJ0BTOfjTMtSmFCFvBOcQSRJvD7qbZ6Eqyv3iaubcx0X2dcbq+tIWjSFNNoT0Xl6epn8IcP85L
jHeQLzyUeulIlqYECDW4NoM8yvT54I0ju68aZFxZNXR0NH65+4Jb1pvGl77vhun6I5E9uvjg6cXE
prfRC+5aCXnb/uk+kM0KuemI27Zq0bVbNca9f/hFTyDRM1nId3DtlyApqAQ6VOHrMBfz616l5oPl
TrT6zEgSrW34LtAd4LO3+Zl8DXlaipDWXcqRMp1nF0RDmR9YfEBs3UMDWkNAR8HFhj05hs+uQktx
2TvSt26cv9wdCZqsbSZN53UsOlrcrHRaEHB7BREIHyuSNcI7LHWhVei2KD8F59bXhYgYSk4urxOV
udJtUrh+4otZNjx3xvlnFwT7TzMh11Gr0+kvHFIlqgotZg6kwTn1nJPKzGF81fKWGa2/EkZXlWpP
aeRM5cDqkw7QjN8i8fYTObLroV7E5O87STEdi0v1u2dLV4VhSbgl7r+BaOkcRJTRkfjLAj6VAZcr
bz9+JSkW3g+NUSo74ld1eGH1IYQQR9Qn7rwgOuJCDC7tyk3WoOidd3+vjQdhNVgjHTcP9zjofE/K
YTfBdaS5Do2qfxqMDvTci/2bl7p0Od/EgNlPlp9t61rh0MAq5JOlr2YbG9FDDALnTUZ4SzoD6oBm
q7TkVxeFMDNruhPZy0hQtpyN35+rDqtG6JkW9gnEdiwP4f8cqzAClVYkKQ5d3PIR6Z4JmQRdxHY8
ws0hSmLUqKsR4PPBIcD28T9rGPJGLDn82yqCvIOFCU/rtjgoeH6iezh/O/g++S/YelNFpWbscStm
faH22hxB5N8N29IXmZZ2f2scpxYRkPRr1EaUeKnOe+4eedNXNa6kvai8P82co9eCPfP5z6H7F4DP
BU3e1ywgeD7v7/mk8tCs1OFovnW0VSq6WcXVbiKo/hW3m6j3Fq9J12xVGdnabLyDcGzdNbi9wnVs
oXJqt9AHn3g8J2WYXbUl4+9cCy9z1flgoqDGctOAF3evbf1CEV477JcTxIL2XHb5bRkb4ZQJiZ4q
r6Z7G/cMyKTjcOF73b3iPun70q1sGe4HwkbJdjzwYy24oLe9GHwPFCBdiu24i/oaucfBsrzJO9XW
LuZSrUDOMy7u7fZJ1QFlglED2CKLKemjw+OgAzUSfURWFUo62zX5+Aa5hbgFBaRn98QZvqSGPIhN
QW5td5ECvsu0a77cmozHDOMS1419izZEPD+P2B5nwKqGQcTuzyYJsi4IVEveOdOcIHfhbyYK/VB4
49YpzItJGJY+v+JNLMsGJ9fDxt8MoD+c1BLUX5nezVEQCJcoNxhy+ae1Padr5x2GeFRlhpnloGU+
piN166lE9NminDqSsrysbK3V7rihQooG4CJMz3xEYnqT9kqYV5eQMi0NolEmuXZDHbCpAWB0RneJ
HpDqTPXx4nqDGwHAomQoQuHkLsoXb5f+G2LbSkL8us5bfvJ6MbU5NwccAManNwZsX/LX9CAISojF
uHjbrXUmbKd6c6nzsL1bRjDBOHcyaYkdF5LD+T/dSq1ifVDQj/g1yzDPcSdrxtobk9akyaGZGsvq
ZgziBNEY5zHovADvXkTid/LJk2X1QpcOnHHNEdAmp4rgKbVz3dm1pMFgq0uuH9t2FOsW3G05NWlU
LovX+EXh8FUEaiY68bggd+z7GIzWdLujwwd7Ujqli0t+pQpUtHBhT6Z2ln0MQu9rUzJV5/0/a4Vt
2qB0FcCRIczjQ20+W7uqPGrxVmlViLnBpf7H+3A/GGXq7H0BNfHJOZpyxzYFlHbzSVNDzwpv+y+c
qP9SFJSvmca9BkVEvZMCbFCHV8iBRY1KqkzwePYT6RCmqLDrnsg9jqZ0eRi+whYV1xiOsK/7UA06
QxYcRiBm4NQueTFgBSUyV6U734HmvYTstY7jw9iAMI77PJ/Ter7IxiGDN2X1EaUsuYYVz+t0+0UT
Dqsnvj0OhvIibPB+lUEdPVXP0hq3Url+X/+MnCbKJGx9QSZe2M1qcnPzk6CZuWLtpfgPR+MZQDGL
lGSyc6Mj/73N+7K30kExq43gLDUUmhbvQ5G14TZqtfO2A5ZlHb92nEjXvmCjEf3C+pSKWEr2OPoV
0oAXerjv36dF9vBJed35z26jIUe7NmuoKzQAszpo/GfPNGCrqVm4Nd6Mut3qJsNfmBWGTEpeNU6R
09jTWQSjlvymdmiFFisCZKZEtGNKfPe+guA4YF/0uyf3qJ3vUGEfhAXT23GVBNRZjMxa6ZVo7WIu
ufAFZ5KEGeYY0qG60xnrirDRrfq/8FTggiKEt5FToU44bbN2nCZvw/CttqHwxBgoRffqhwDF9x2V
w/SoFUMMekS0rRcbuRNf9/6UWGx0gkigqMSCa5b6WUMBgd+XZsmVNIFjk49TMZdD0Q34DpNs0GMP
p3UHIC8AlLouaxoDV+81pZqESfMWVThJ+0MCOXpbf2i/4n9RK8e+j9shJ3yB4soSDdVU+WfU1wMB
4AwRuo9QKQsIVrGs4WV4C6tKe2lpCzesjUwpCFDgoh0Ne9khFW552PBmdrKpQkszdWHC+5WUpOnB
OW6IL5sZAc7WwRuJrn0SfT7D9yk7qaz/LGdRX+J8lPl0x4G28TRwndiU1uV7p43sxRWYDWujug4p
Sb1xZRwMxEJf4+JGcBH1gjedyxGAnKKD8qwzekGjT7kRcpP0FZfiye5PiYB95LNt6p3H2nIMnEgF
02Mxi07/BVfSY+0O2DZweReHFE6mEXATW4y72iTfW42Yk7f/TJA1EqWZTsnM2BzD63fPNiC1L3vO
bY8GYOYsa3JM+f0woS3T83xJYIf3MKNkdpaoO+eUIvYUD96BlLlVvLERxAWh8BEfGfD3xQaqQhfy
D5C562SyR/r1oJT0opJx9i8kkuRdJPaAcP1q6IhdqhwOzDJKBs323/2fXaUN8FnvwCquxt2BEA57
rxcIAPNQ3qKmJgQDrxJqvFVn4w5C2ZNeowrntSLoGKYCE0XkWmZsfVkeYTZoIAtrlrbsMFny+PkF
uZJEGy3U42H0JhMTBBlSeRCQ5zogcNuOmF75Z0HERGoCHA7n7VkYuhL0vwgFKvSsY6U5/98D7Csf
fw0RauKHDhVROslvKGaViuBJwSm/6sElQKf+ffuG46XtMtogxYzbvj+MxMBjJwzreoIcSYbbKgsK
yAeHmd8bEnzp6eUd3x62uv8t1BF8oHqG94Cne4ueZYxgYkBcKKYay9nxX02IOUSf5qzzHyY7oWJS
jkwUSBPNfTwab8YFbqpNR6tj0CO0s6vURjgg8eg/dbfiwAXwSQwLtucHnUR5xvWxMFNvmPene7e2
F3sHFon6iypx5H1wqkc1yp9xJuxlwIbduj/Es01nUfhY3s6hykT+Udgd8bVkaUIiasnYpQ39t0DN
ngoKPqY2dSwTVtQRdTWsn8WjYuj1OegP8jQDbqQBFTeqfhB0mbjhI9ldIuGcly0WNS0NCCaN1Zkn
kRuy9qZGwyPVmK3vW3VWgxT6rU3Qd4MoPpwFsLdAw5yXsenoIT6PHT/ROnOdao4WbXHwH4EXYwM8
DXsEzaiZaJTjNEBzE6cmi5hU3xh/dcLQZ10k9n+gaEEMkA/UUzltTAUWmTsj/czehfHgjo7qKYeP
8WaneiuCyQOU0fQrz3V+GPv/S5GyQ5mJIbmSYLZH88pnD2ErSMGLXpUdQ5Zq5PM6/6NGA1Lw5Xht
ug6+430rlreVXIoTtbCwH72wXbQ8HAoyimzhNk1pKFwWmqwgGxukK4Ib1AOLnCy4lDNGg8SGV/2A
+3CvD7I7n5n9Nl6V4e9kWVy1bPT/4w+CobF8CTwN3jaAE/Jk19po6X3eTijFf09QvH1ufAOEplrJ
qfDNplwfO+WZPacWeN8x/1/fvLk1cl5CyXm5VQmM1ZrKmETdTzUk9C5TLAeMan89Q6EA5+oTPgU5
XPhq/IMBIR8JlgJYaDD6nKueJxk0BjxGQY/MgfBhL39a6ZCOjJ8b5f1M1myAsA/yZENZXuqk4GaR
vqm/IbWmlmuBwG0McysTth3MiT52XovRtbRxIciNPXQBvSsrJij/6WGJnRDbkX1ZXm0XRik50/wz
MYDUHE6bcmVZnUXV1S4ysyDstu51I0dFiUPDHba5VRoghBOQ7bPsL7gkl45YiKpAs/h5DGIcBtiK
9IdCUXsDZCNEIsrwjPOZNFQd33N3AE0NZIejX1ki2eaeVy4TI+jrjVYaLQPzzKXpenDsgawzAiLf
aik5IpleaJlScYM7nQCZqcDzAxXy46hXP34gOPRRK97Yho4HSsHG9QF7vyNlpr4ooclg7n+jpNn4
/zBiVafuJMKDR8TdW/IIhMMaOjS1GkfW3qR7StvC1bViLlIxYNuGp7SwC9BiOvRjrx+h5nS2xbvC
zDZk0O6IKw1s90Cq2p8uU32z3+V+qSgAs1p1NIzo8UpGTe7szmzYjwiICNTBoGbTUXszVN9a2XEx
Uhgrzs7to1lPrLwtqx2fIvvFxEqI4mxRQkV58UCw1KZ48ZoMMxwMR6Y+1T23Gv8p5hhW4ppk/FC/
DpBuqSzIw6JznkU0YeyQ2Q9xTW0v67N8NQJwmNj1imr2Oy1RmAwYsXFznky0QQKbkth+id6k+iey
mamrVD4DkSpRfPq3q2n9IOnl/yxXkNjuvJqPYhYolotyoZEzaitW+vgjKhlwOASui5G11QeSfwuq
DE/Zzk+gixe5MBUCG3LooCW5I78T57aI3jKPwbkcRIVuqINYaA9ebpd4DLGr8gN6peXee6mCOnDV
gnamVLhhGllIA57yvyPRCIiKFZs7t1AmPS7UVONuECF7UgtRndsh+8avC1BlMXeFw+2jXMwNsWGk
oOPdYAZQXXBJGq8w4iKVOJy8zQCvO37+T6H7EYnDhh9Zo2YD7s2I2G+bzsxzcoDe+xI8Nm+Eq3zQ
GSuGRIdlm4xlxUwvrDuTXSdbLpKP22p2n/UwwuItoM9lSit0lUWnUinAuIhhCQoGAaiSoBNKn21o
2ed5KIEXxzZlL6yRoxXbh2uwfWDLpIdfUqHW2BFcYkerlqpP66Mg2IFL55xjivgY8M2a9IYidWkH
4sUdkdc8m+DCpDoJm02Q3mJCHVqiIyNRhYoBjL4AMmneDaGTVwWVA/zlo6G2PEXQhkHj7YvBSuMA
sUN/s40qNfZ0IRO8Q0HmftGLM93r+wEqNeZu5xknmi9JVCpeHpuJgnwcWJ/T/qLDMmMTgpCdPLeX
YeDmKZBXuwUpNcT26su6l+iR7bgPm25nvE3b3lgTVTXH8Wieb71GJwm1djZ2JGRlhydop2AeoOrv
4mjgikbWWaTLDbmJzGxyERK8s1vwm9Z7j/hy9xha5AAP6I71R2ucba0YZivyT2k3i+iCIhBdLLvA
K2oHfi5o122cmek4bsRlfzdvw3ibWfzxSoVPPkjFKHVBMbU5KR6MooLrII+mv9dYx3sFbTg6NVn2
O+uQ9P1aXA7pROv0eb3KmiFyvJXH8vUGK2iPncWGFgiQ77OD6mccQaU3SR33uWYN9npWEEPNSGE+
5Q9ok1X4JAialtJGicBz2WFAB/InwYi4C9XEuAMTyGewTtEjygEHgzaQp1j9cNu2brurgL0arVaR
VgiKtIXe/VBWLHqGXS8r6/Mh+xkyq/n4sTqxs49aUHhK6wAjorWHvxlboxcgTq+Wi1qx904qdYAs
4YoHq9PjuC4lYvSz0KISCkpsJzBGx22rZP2AfUBhD9rUJ/En6j5aubZNNzBKy4WkAAebKoUz3d0x
Vi2a2UOHd5Tl+q6WvR1jV43XYNJc7pqeUNylyXRosGpsV4QNRYUEiZ0QYE+fiMuRWbDDdg7PJrKm
4Jpq85X39/wap73IMmj6fMZThOeMOTCHo9kEIH4xZKESukKfLXf/MEMama+AcDrHjZonBy4qhy8G
x33KTFu/kBf5knQ7/8rVx1Q1nHbmWMt25y+tu1FDdYZIa+t8hjsKPHieeGmWXkpAkPwZETXhvADk
w5DXO+bg1iEcTJUretlrhFq3zmFJ43hNj0YTtL5TJBpIYNT2z8TlqviJt5gesDds5rua/DxVXUwc
d+aqVODxYjQKi4aPelS56k9NyT3wx3rYCnkoeGzFKXFFGJaYbiAHLeUXpJEmtC1jOmmjplMmsH5b
632mvXy9m/sFuXkyXJsbqSuAjtbROiVDlVLo+FVFLSPf+J1fnFkdf8ByCdfpF1OJNbT+yOJ0brLQ
+Pt9DTj51DjC036Oop6YPiKrYRZv+oad89TLx/f+fcah0c63kHaAYLgXR9NhFGyprfwWsKIsDrWy
me3q9CwO9zl0K5/EOdWatT0p8YRUlyt4dWhIY19IOHjKlFrPcKCipDOnZ3MIg7It9BcTKbAV1p39
IFD9V4LUc6fR9lwzMR4YMeY8kQvqLP6vzTKSp+fPRFlmRXGAtDvF2BIGYWVCMoq4MBSXi6ciGQQF
/ykYgi4/QNG0LZMBRAHaj6cIz70OOQEC0dHgEEEsC3Q793pDdvlbCcajgwcUkUy76wKZlwedeikL
RpLLKiP8oA/lO9uCdvwdlSJ76c95IRB4/VJL6bDI16kNO/yC66Eb2xEMD4Nqa4QiTjxRhFMHmJHl
j6WJT23bqCWLcH+W14IYYAsxix1zU7iaelodirecxyApOE15BYbt0Nj/V1NhCsFjPWe3AXlMrDCL
INf6Qe0dDU+3J97cf8mtNR08BLVVTUjVzOB6n4iA5U+3nvRnHuqhm22nqKdY9vaWwDDQDt802DFA
yvzk/t0tifXarkTa2vhWtVc6G05xyh7ffINKMSCpIEL29b71Lwe7HxGJP68E3JRTkn2LVlcctC9q
5RXPy1+Wvc4WWbb7o0WdFLzn+mjROFeLpq/mr0V2DMTNNBWVYjCdTin7oBcwuXrjHVQY1XyoIi0P
GBlos/9n5RV9JWkqfErza6HUM2pRLUw19Sw10PPFc8GTNHB9ka8FpI8xQQI74VbWl0sXKfNijxjI
wh6vExdzzmo1Dmlvw4SyP6IkjoZU7am2sWnZiXAQDLmKd6VB4qY5O9h5egc3DOUSOQvJSmBZ5Oqu
noxe52m5aKFyK2AvKj5S2Snxfpxr0TbnZgbZ1cMBNMwl93pTjYMMca6w9O8MeLbCo7b6BZQqGSz5
B5xGD6xmQ1A9Pl8928RSfxmkvBcznTpqYyR2thK4NY5MveOgoCmD5SQ6abY4LGvyHpQJPEppFADB
VAMh2qRR/QgL+3omJfFpuYrX3hXy0DhWmMhStwJxaaiEvfKyZbppMdjOKwC32RGAjUe3S0gVJItU
ZEweKFpaW7ejY68dOQzktf13s9k4IdWiFeow4FbKxVu9U4n5D3sNnutc2j/4r3GaHjYVioO80H37
Kvl2XnlNmE92E3YpSwmV9H8ggrLSKWGyDjgJUlgvjxTpfGHQc9OdQYaWODzPGXwsjxYFGHDNuulh
iY4Ho4iKdBJ/xp6pAathurOvQpL1UsLNvfe7XBGw2KcNkat+NLdpk3NHBI8t39hHVs6X2KE2xofU
quTQFblxRMo+kiWrh9rHVbh9GNq6TNFbCRqoqWAzd4QYAV9uywhQE7/hqJw0oArAFQJU74UbrX08
KUkC938g/3c/2rflY2YcFY4GgErd1anDSgRtXfO0wk+r8GnmOp4sHSXoSCVCBhITIbw4qZ9jv+i+
0yFCT3B1RGmg9x4ToKW+EpuRE/QtT35yPEzX7pVzWylKSoi0CSyw+QRDUnj5B2qebqbfngd0WR+u
dSIUj53JeqF7b4pZ3/v5Tpq0537MrSPThm0ND4aKOEgnLPHoOpoSPxaOWXDzi/Y07t56BJ7mTTmB
eZWQpIYtF3ypQ3Qh0LJRLYKpq+8J5BjqkjUU9ka4i2moB/AC6LtcW5fR55Z1xa7Eb4BB3SjeFfln
lCeb8OFhtqfLnVRi9COD4j6Ba/hJzVpchkZCJzi95GY007VyPjpn1gxIXdfCVPaT7wOrpdAXcSuu
eG9Izk5qWN+So4OZwdNCuNMj7Rp5YHT9Pea2fFAlpijGn7SuagW6XObC8WZ0IQqC5p5bEM9x2/wk
sHFqTpAJAoudBThcwAQnUV7nT0LwZNZbrlu2Z6c1uA/1Qu2nxY05DYWRaXK8jDUW8XgGwFg8lM3s
5aQppzClQ1DJ3pWLSyP8r6MbZY0jKtkZo44TBJrp2Y/5ERgcWGhjoDGB/9PesdtlrTwcnd4EaYDH
yK316GfW/1aiIKnUJJoCebOOKbi+ZsbbdR2yLdDQiH22diUKdqJecmfL2EeX7eKI8tAd59sNBEmT
pgIwhA3QhJoCqDzyydwepYX7NJ2mu1w35Z6hGF0OFzJM8dQv2b5oUDZMMOnR4+8RNpdvF/MUWGTb
Q5ppOXy2fIt57Mt6jNkt3ZYJaYVqRxiye/vJcCVpgFQRiE3CnXoNQwWl0NH0WL17zHiU11yhNQUc
zs1vy5RM99A2jodSFqr/HvEZ/nde28dB2yB0BkgA878ZZ7VWgi1u5WRs57oyRdZJRowFWwzQozv6
K7P1KCtbOZTGbQkWuz25el/nSxLnDGPgKeUdH9JPvHJAWbwiJ3wgmQ/EZ0mMoEMMReFhmZCEsJMm
DVxYkXExfzoc2B1qlNt1UmgVOW4rIrD0fwmS85Xsro47so6+PtOz/qfGBatn0FcnNxsXiR/Q6x4m
WK+JiBr1V20MpLQnF3UOmKVtOcdV4k9Er2grDCQIZabEFgIxYhRRPitCc+tGEZsbFtIM3hHgbD8r
M0TDTzX8UdcqORsChK0MEgAXEj/2YupvFtRhNhK+Xn5YrhL0q781BdPEZm5LEjRHnkOLqqX/C4zR
9Pmjbp4w9krb5ih3nsDyq+e9mOGH45kN37GtB7ZqiAlPWeZoocD/DZfsZyQNmSKThstd5yZToOwW
snBgnbQwmQF5NP+OdffTFqb+Ie7843P1xFEO18vJFtV+uGUjAUYt35UwRXFnLiPt6XHLPs5i/fK5
LVSnZIWohNRcXnKTXsB27CISyfpN+ZX9nBvpFFT0u0WnH1k2OiHgMD+Q17DTBRhwfcP2lxj5klfZ
ArnVdMhTMctnOSqSLz7AF5s4IpgsmkhpYzqHdbwEr/bptZZkrBbppny+MpemXeQv4s7VF0xeGiFo
nAAeJV3vWMvkf+SMFeyNJe40Cluait72YIdxAiQkJfVGA7+DqtfMF/cyD4bcdkzjqnxqY0t8VOLM
MjWzNk5P06ZrgZZoxrT9QCejz3F7uqZ1P/liflfMTlMR5fA8PbHaExevg9dYeVIRbswdowGLpKyS
vjTeleaAVyIWM9gOuP2J1ctijePbMRjI2bgCnRzmcOTWKQRh6iNxufoycWtOyF3M4TKtDyTVF3KI
KxKPnbkU6/Qk1rl4bKxosv6bcfCTKYjdnAykOp2nZr3c/ZJ+Vhck0fjkSZZgGPL4P8WLDxMuLFaW
rgjD0MIUua4qgdaUsbB7LuxFYpKnA7j3IbR78shJQZWDCusDvVfZPJ74G+XxRqpgkv3gxsJh+uaR
M7335TsRvHD02xDHF42i/5mHNxCy+QnwKxrTyxCz88xy25uO3pO39QlzWmKi4ro8tLuGVDhDx8ZI
KaiBE6rySP/mb7/LvHivAH8flztLtujpbslQX1/JB5HCAjRawFa59L5ztLIGD+lImbdmRmLiuqIM
JkHUxjzfvS4MVeVqedG1x5nVQerUN0Q3k4n4oeIi4lU+05/08WfZKk1G5sHXLCH5Tv/ZD9THd+Sb
BVXTfA+JlwybYIjMpVrmtDZ4hQop7F2/qT5FOHVtO3eV4vIjTIegIINiePOCLy7NbQAm6sBk3nYU
VFfpVvA0sslWNQgURyc/A94x7ZcnEzlt1xWUkKx8VYMYS6x8oTsWjUWQpJjVVgKcTWEpOfBfRp/W
8MMVCKYcfAq7RRO2EGOvr18J0bPAlY/6Jm/TE3NSWDwL2BDVdHe/HNQXYu+JAVevXZbkvcFtea3I
kTsjjFJnTaFYiCPmv7babPE6byu1jy2I+3d5snM1ACuCwjDT+4NIBQw2B5z1Wy0Xuliqh07lxpkv
hpyXY+OaQRTKRIDpK5z7c5lomyjUCPGlyinp7egW1otPWMeyAWa3qfnx5greV0U1XG+D5tzG+iiW
5dsLn87QagBNL6wMx6AZcGK5cT3YJtyL2prIER63FncxQhOvZ+NKt9aA4ME/jziCM5/NcuFkeYlJ
Dwp9AMN8CoTnQmC0LmdDGh6BLpZt7QglMDLFK/1sLT2cGZ0HquZi40fdPzfHRr6jKJBpEXHYLSh2
yV9gkN3Xr0u1AJzN7j/rs7O47Jg2PCdKCv+XQQ+LReDdAKBB9c3tSTVoNubC57VAOBii5UWdHylF
+dXklZLiYCq0ovFWEq3mG+XCSgkFW1MhKNlGPircfhTM5CMTf7xatnJoGhzDz1+VTjGu2oDkMVcN
gSbAyUpg+LG9o3695W5CoyKUDh+OPhvCJREb8fMTv0kbzYQ1Gop2wxkZDbazghpXVuFxGN5ErgEK
Y0XDi48yhpYcTRAIUS+IQCQgE+mhJh7zeziv0o0jyADalMdYuW7DITuh8xQhsQr+PrnvKsZo5bWX
h+GCSyBDGsj1V8gY+YgrE0yPDVMmLtEx33JJQqMgFzmQnYDAEoMytEw1fdjnfnC3OzNJNv6JZK17
YWproKvllF2E8ybLnV7dbVgyXAoTSGMWMtFZDhPMs4zdq8E1FwJ6OIQ3iWscnG52fFwgOBChEx8c
Vxxcn60gupOtikzEXTRexefPQDiDd0CSkj17b/mG53SVoKZ2kH8gFHNJBHpI1Hh5lbKiotsq9GVr
9Mj9r3SO5yR4EeCC5IZ8p1dCCQrP9Zdzw3UJY6r2OrSDqm+2sYDd6PyEEAER2keJSWGwxiHOawT5
NN4BQ41XbikbdPjH+kt5ym9X8w4wX8QAzeVsUApIacyg7vlT6ciAxOYtDL2gHiuo5tSX3ZpiFyzQ
+zpmYWYd2Ccgzxlp6chtCuJn3yW0YRYKuoCYlo7sxjzqcnactpNrn54Fs13KOXFcL/h7tjQ5crfq
B+/CnhoM9Aq7PmD1ITu2usXzrNKht0NDErO3fd97033MLmc2SshusP8E4ygZOKxCSNy9DKh71LUr
4W180Qg6JaZ+MuLn+FP6PxSZDGljHVzhPM0vbKsHJKUii5LelukEvEGSvSiZKKbnjsZvCGCxRQL3
ct1XO24+QmeJ1tmNYAjh9O4Gd0X/PQf2pqqI1T9h4UtiiZd8DvcOiDhMlMfMG6aTLcQv1dAxkmis
e/Okkp5quXV709EZo/DwWUPNtAks4+nY9q6cOPiXEX6CbCvTZ0QBZf0kPZL+kqCKoj7iwHO7ICnp
iX4WN74pivlpBX7CZpXT1XWZWqHNUxR51oGXF8ieVefvo6E1O/jGHYfyVdUfETEOBlz4KiC+oQ5V
CC/c5roYXxoBBYoLMBioYTmCByysQJ5o46YZfuSvdvpXcvCDnwrKGCpHW0/2z2rXbvzgcEt1yMdc
odd+xaog/ZDHpIre2Bj1AY5fBGKK1izTwNDnBgUgMAK00u5Vj6CIxQQFzghI5VEaaHiDey+sGhG/
CJP0lLEFIwo+Dt7bwxj5epQZVSK3C5QkR7QxojFc6Ddhrkld820YNP3KWNIpwUrIRV4c4JBjId7u
tmUDrL4FYDe31y/+KK7hpdTZVSvmvLXCJONDRz8WkM+beKVXPV9hxzeZVd9LY9p9liZtBWBD1hRa
XlebCX2ykW1kHyL3v3jzg4bKczdfbx5oWhugwEaxEx7BcXNEiuHeaUqIByDg3/i+Bkwd++zFCXCU
QRJspqvqNl5VClu5iHQTJkPop7LkSl29n7F1LzRj82ecFJex2wPSzFmunXZCrHTfMIE4lVGh5awC
ndQPfQHf7VaXjTvL8mY1R0fJcSmRUjOv3ypn3d+7i7C0tdpE+54nLmX8F9ZCXoiWrGDnmaUyy1RK
2NEUgOnIhQ6BuC/db7b5khoCdckFQDtKuEqpQL42D6+fFMVtTviwmzjq+HXTMD3bUVgM4vik6/1t
dLzQet9qs4oSLx8RdHUnImiRnI/73KVtDl2l4hJ+tUVVTOlrvtsY4RSH3ZEB6RIN7bdaV1Yp7gDp
+qUU+u/YkV5ayj1hy1U7K1zZxbxrf1P1ruywr8JwJPwym1GoGNm6TZKSo67ZqeteN5JUzc+H9u6c
5+fXEhh+XCNc6KisgK/dNnGQoXFpeba6TU1CQEZSvHXLKKpRNv+Mzptmzmy1g7mK1RJEA2WYqW/3
a2lz3QDvlE/mv3mXsJUTyEA6nHzOgqR9Llox9Qauwz8oyxc4lhq9OYlcjOi2UHBBAGWDScQO+McG
k6XzkVQBXUJtjF6Q+9KhHEUegxZ281kAaXqRIh3P//Jv65AfpPoORas3EMtbTJd+pwVl5QrK9MNc
elcgQFP1CeZDuVZQqDrh7eDkCIBM6DTdNxvOK/AvgVnjzfk8V2FlBUh/1zRRGnut0PirgwS4L+Fh
MYX1DREvOCRIIaxYCFmt7PSGvfG9MBTKGbu0ohKaJTzZrglWChd3KEAoCM/JShABpr/uwe8rlUou
+/o9pDrnsvMk3J0R+Q4rnfKpRZoVe0xoqOj2Q6YhD974Kwj8qlrpxO5iEusr4a8Vp90CNUTePjba
YChX2jQPe+GWBbrugb0K9BmR+y0eAH7FrxQdkELWIDp6li5IcBCbgiZi1g3V9WViSbA/XS5HrNNI
W4zK5+o81kldEHn05eSx/p+u621Ez3MQx0fjrfxsiDfr8bWeDNNXeIbSP6N8pbByKkTHJcfYoFt3
/MmeA0mtqyI5/tu0FjOaffkKMrnsjlxGjV4IhH5m85wsORlHx6ijXK9ewbdHE8HMMNS7E4V7L/1V
inyF48E/UB3tittWNNKziN0Hh4EfmwWBpNIK3Nrpjsxlgb7sGgLjP9DQ6M/kxS9Jfak8FvG407KV
lmDkRk/bH9En7AE4RJKj1quM+eGTCi7/IpAhyVHm5o0Bu18rgXVqWVDTU4TqLfbEfUR5GYMd6ylq
Zm29ZnSfHdiT2vshbcBoxi7W8xF2FQHQlCRXL7STfCeNIB2dl7Niyj8XOB0Yqxnv1ZSoUz7UBz7P
vsmjD3L5zSFAoYrGVNxfxgVuboDT7pjREY/Uk+euGoVSo/GmWu2fwzmq/oBs5kRkj8BKCWWR7g8y
en4nz/ixBsNQYwkKbE0SufWn97xKy/9zHZMWf1w4h2K7wuuMtvn8h7HkvrPt6h45McI3gSEubn+W
Pbb+UC3zx0PormCEu4/rGEOIlQYK5VM+h6qMp0f9HbDSZEBnF/7UHFsX+t1h0NHfgy3+xROs8+df
ENbSCyM+A/KY+QtWR9iOTZnlpaOm3YGthEHRm5pEiYPqFQF2Su/BUQhMXn0MQDySu9sfIru4iF+3
9YdXTOzprDyulw6cF8wS4J2bvGS7ASnqofFGRL357TKHSnShCdu9j8JGYgT2ZnZQvktErpmGXmtu
/xRG5kz4kngHVz8IVRKF9rISQ8y8xMD14DVj+fMD7WRYm4DS1uN8axnOXq1hADClt9Zxed864atd
Ml/LMaQiyB+W3ehH/n6LpV3QGamSW5KaCWQr+FB3ijgmmilbrowFLdinZHJXQqVLYcd7KkhJonau
1pemJdC5vDw1Nw1b08DJncHSh7uTiEjQvJlNWJ2D7dqR7QOUupsebRi06WR5jRZwrhKduC6cimHc
ItZw8NPCpKHhBPZ97ZbJWJxsXiNWZXrdhxDKWnB2FS+gxUBqemzestSYvQGqDEIy0P7wEEECV4sX
IPIn6Og1imKQAdhRFs0e5Kk2b6mlXNRsTEdCnijBOXoSKl14j226Xm7Pa+V7RsZQ/QA/zzq1zKXQ
4o12lnXmMaWDbGFoznPBeQ+0UoGFRkJcm0EY6flK9WTTdt528v23tf8EfxH9tXdC0cz0WH5P5/vE
CeamRAzcErWrVt0qbK+zsSV5qzOQ63b9ne5yfIhgXEGLhCt5JNsrMwowCPDCAvJIjrbfEEVtKnvu
ydCbOQgp7h4UHgke3+H0ni0BnPSVmNZ2WC7I5/eCkDeEVz/2mTezV69BvkEggAXBufJH/HXymVyr
LbMnqWgk5vUVgd0ZiLGHxszjIXlKy91jUgvwQpXVQjDUtWennD6aDxa5x9qnRgrlY3KiwVMg+SpW
J4PqEG8p/in5UWPssF6R6RrWbnBXm60Xg8G/Ei2ujOU9YVblIVhnOmzXF58e4u5uJ3nvbtifgWvc
+oDAQaAx6eEgWsz0hUaOIwRt5Mnwn/Lx8oU6rCN8Y52RckYLLu1KB2/xWpIunrFCGhO2MyHV17sr
To6aRs8eMpPitIqkrsBBcEOpulfaqmCuvsHkW34Ze8pTwebzoEsU9Z2R46vKlo1RoNqiYyLlRtFu
AQkn20wSKb3fMKhu/qDjzPIdINWIOYWo4V9Iqtc2PGmWiBDAi3bG59LMpUi7XYPZE0mVmzV8Jnu7
jqHbDOA6ciyT7QPqdGB5taQXt8lfOu6+ffYMpEp0dRQACIxtF8xGy/sUyzG+7Rp6sn/CqixpI+9K
z/vuEs5XpX3CnNBvBhPz+tgTahh5ilxJaVPnbdRtmFxgtuO743DEelNYXQrL5TUH+O1uTgeYB7av
HqZm2FifuUhakIUNyI25wFvfNLG+A97LN2pZAoMfu3miqP/LEgA/+pGhf1uAs2kpmMCmraZZGS2J
2Sal1z2jlDZIQ6F9ovmVBAiNXKS7fq6d7Ge0OZZYryFHfIjtbwv6uiFjJj2EtQnmtYf2zew4efZR
JzQ6X6pUqw+XW3xtqkRemzSWKP+bVsw30vI+ASyBpnWUk8pQ2BxRmToEKIepquhf7SKNeG5Xmope
MiLWQu4IwJKXi8FgD2x/4fcs+EPRyq7vZFSygyJrwAcG1v9/fuyivg5qSg3ofcaPgRGNY7m4Vepj
tET1AkqaxgABJX5HOBlGIqms+7d0Qe7XyYRyeU64MFujNBUpHoxrY3mn3Wd2eMhuP8v73XmcHPB0
V8x6nzw+k1SLvPnMwuaOCE0kjq5QC6ekOivzSAcB3DMT9NSA4C+lnmwOOxy5XEKgiJojd0cExxlU
8sdjDhWxJzUdTunuAqjJnOBktCF6w7IVOgMr6pwBoOsc29hiSEr11Xic3Enzg4bSwfS4OEU4i7Qm
iWK5ksu0n24uF7cyY6vCc8qCjw4ZHvxyGx5c346E4M9cOZCF+0nh/E7JQgW9asqElyhol2cF59FV
vN8DbeO5+88smhQ9NkieRruKSty2wNl1gcAC3jHz14AyJXSpWypxbg6ktIwUcwUAYWRGdyVNFYqo
W0csIeyw3vJfb7dZ9WGItS4XUBF3jpoaIl6AphX3rFhrRIKhVx1hR0QJ3sVnZIgfizBJ4RZOIyGe
x7yLhRsUGAdxpkmIFWThp7me21WHmzboiL+gc5ai1S0YuttzX2DXipBQD2TsEgBQjPVPJMsiLMfj
MdrkudY8mId6iGkd5jrkGj7greFerC5wU+SVWuqBhWIy6bpPAQoDULRR2WhomtQZZFmzyf2ksbw0
C9jbQyqvjt9SzjHH+tRG/LGLxTaJYpNFG3bWC2ZW/ztZ8KGOgke7umRFqxbJogSF2wFQmJESrYw+
ZFhfoJ5faYUrKT6oGqduXRmCqhyI2M/62rxFARTExIMEgBiIGrDmOM9gJNJ8HLH2SM4Gi/Byi25Q
aG8ooAIxPNwPTDCiL4rTkr+6uGEO2W8htThj8rk2azPgkQjI41gpgqcViRwFWJPzIb4UA4E0Ap4A
Wyw/qtCX3TEEhlhDiTDjklML7Z6T5Zf6h85eis08WW5sZFR3Ar1Jpuj5I0CZoaHDqJ7VOTMorLhz
TCbeg7Ta3G78RSKFobzoTtLB/OajQWeSG4rnwYRWZFxWU2tpeaNy6fmsaUS3jRm0VDGMZLOSYhjT
uhJGFeu+WnHx+FmUMNIPjdgkJ61W281jUUdwOlmd4JI9+Fs4quqzZqiftwVvkPywZgy5n0+TB0/0
BjmWQ6KUE2mhVVQM9pEcjoeimscPf6Xvb3Ll78Y6KZDa03TKmcqaI5bHFn9+2rkAE0lTymOvzdH7
5sqmD66x0jFJVaJOWY9QHKh3wK2uaYc1LYgUflYf+D6QqGxEpEaoVEROq6u2bSztRgD0S+9jsgCL
PyIwjz40bjgOk3d9e7NFUr7eby7Ki2yGrKtQK5u2mRCGw7RY3W7RaMONIQMSvepAq2sLVDkKm2p8
A4jpFncubJmtyUDYozNUm/muXOX1BmYFOp8oqeu3NPcl5UW/S8J4oLXg9tNZWVTUoDc/yrTyZ3mG
nKY02x15NFfZTlMI/vUeBIARbd8I7Q4pPDM2UABaIc0uJN/fnzJf2qyIx6Ea8JGVG5xBiy4lOvvl
Lbp15b4MDUYP4rhO/HUrewMLl8/L/U195jdFnxNPArrQ3pfzM9XSU4hhv6g04r7CndGVMcxiU0JG
Zz0T89+90XH9EanWKz/B/UG6jBbFffipGm5k8DBzASIrh0LLU3xOfBP41fBG88W6hOBwYuFLrN4d
StCelgQCdfAPfG2A0IjV2epVclTLxmWgldbzLaCcJ5IIX39v/8mgI1WC0xuwED0XTeEj8kp9ZTnQ
uQdBVvfH1cpDXvKG+LUirjyNc+HRKmkFYnmUiEZzhjhC3QnRc3qpDZjVjdPGVS6J60puxu+iV/XQ
U9P6KKZhDHgNOLa5VoyFmCj7jKsTHAt+2AghVXsMLeS/f2IlFwi32vDXnpMU43CEea/M5pKZt72R
ryke3gdXSYFBfS/zK6NI7M7cfLk4h8eSejoTnjm+VIKXkY5HlI9mP5WCEK34px9twMhZfTyI7g37
EVDdbw/9JczmF8e6bdyGMdVYc6nQg77h4KZEyBIj0SKiEI3+vfAifS/gYmN3c6xQN0XSA5YR3549
Q9Wj0T8BfLCuJwtOB955OW0egMRr4so08eLu5/EgrswUfZKlR78lvPsccLUXI21KwfW7jsGkidFQ
yu/KlkhXswDfkFXJarKkt1NxQYyUJGZLc/JJaXHVC3oJ0aKEx5SRZW5u3Pp3hCZdYXE1Ot2zfnUN
2Vc+znLY7B49ALAb4dMzgFz2yMjKo+uh4kM3tZEdmEX6DcD6XhTPaJmBAiT4ZXSQRr9y1udE6jX9
1PlzxV8yd5iQnvt800mJRAy4DuzqXuxQmX1jKdeSsZeyrZnHqTAvYku0yainQmQjQOK2EN/xpLcT
Y/ShGpxZ770I74YoeD7Xv7cwHJjjsgdfbXvt5tX6qcq8D4zVUacthVQndiiS8wpPb9+h8M3DoLx9
cVObiLLvhfi7C3beA9PcJxdLQj3r73FL96tNEzTXJr+ikPkdOwXltUFC/20dOxnEOnen+mZNWYA2
I6Hlk0M2FkmD4KLUGDygleGvZyzSqlipa+x9sgiRZ6Q5UaOzhu11jPR0jZ1bUI7T3kR7Tae3gCWW
8acbBL7llLB0gdaiODg7X5NmdsEFoCsFv5xe/DmaRyAxiAF+YAEjIlUw418ziNM1C2+dD22OGWsp
4+zVaft9Og71iq5LZPIvgCDtgQOO79Ro27llez6wh7D04uU4bwlsAPVsa8obWQgN6CjwJmNU5z7d
nPYJgrTXLukpG9Hp9C4sCcJxRy1HONjuRWdOYZXnqvkL4Ib6K33uTMwePufCIU4Ho24J1+TiXhyt
FdYJiZkGAgXQbEDGejdiCBZn16gqBfEXsnQ1qYMWVrInYFTjhTbRdymvSxGxidvmJzwJVGEqleBH
c6HQybg5gHAIqtwDVF/IA+zMxANi2U/2OqCSef1dL2EgRkU6tYwPITRKSFgaHiuV1/FIGbJ6bKb0
tRTY55vJSsTJoz+GPb9MpnHc22wzMHcHCGQ6L0XwQ+V2hSHynpGEu+eGxzD8bx+hCmGK9BdnwVlc
4vzrOwFpSjRWPG8177ff1GwswvjjyfkvggbDhiPlq3QSFUN6YbqpXv76N2btallU5DsEw3tCPmiK
UW3uvOTl5OpW4/m6ag2O5sLShyjV+PSrmRyv4/53Cau9A7kdIMHOcjvKEfYcQIbCtL5bh6eErL28
tyHoO9JyQyeE8OPSRrRKn/wQfArJA/XercVsSZsWcSbkoWnP7kTMA+4FA6FSLYflRHEsrTYUuP1x
jzfKRKjp1Iw8L+b1LgGn+X3DFoqdaE6cHf6YeWleUhzRBMRShB/8cW62vmBSOabKz7WZ8hCcWU1y
uFOwx0LRyrIr4UbeGppM9rEij7Zu9DzOIWzjdwXUKvtbofLaFHZUyHW/IXy1+4deuz08RAsfRfua
1sZA3OfvWgzUOc9mncgjw26CmDDthQQO2If8/vf+a4oxRi5TDfhWuuhMVxljlLjmnXQPr41S+lSc
qqUfvvsntZH5cOCRjsR6L2cYxUZ5nIEcu8IeMw1HcMtAKGx0Rcy3pPcu0yldTU0voix1L1Y3e11P
4i3Ijk6mR1YCoMh0DngR6XKYz9oKJo8tbKRWOdKoVuaf2csgzJK/2SOueijD/rdtBLYDanYubrue
OZ2XPEukpDDlrQGveLd1A025crb6zlNgeu6upiJGFvjhuL9rDOm3DFl5FkLayCTxlasSlNPO+VNf
iDxM8cMmPowawPYtiWHIkHQC3mMUGWfZHXhFvu2yjNZZc5FH5DMx+FxYWimRp3X7MZi4Xcw1s66S
z9wZzMZ/VSu6ArJ6zWLSmO3TgD7fwrMGjQhOx3AcByU7Q7+QKvM3gF2qHwaIzJAN5GA1d7H7An/Q
t9nbMrl8oU4XhlqpPl10j5YhGeuFpvPTE/ViFjEJYyx8FhaqyAqSmbPwMAHcalhNsii+vdbrz8K7
7X8EUCKJJdR5EIPSkrdt9wK+Af8OhUKd5gkrCSCYhJKGU5mkJWJ12t81LtzmOuEVXH1gpCaI2rHm
nYc/TUZVONeLECHMX8qx1l6HKZKMv/FD9PqajdFJSsPFI0kkHumtS3JKwIfbqPX0NQWr+Rbm15Ae
mYf/umjqQHhY21P0dIUPsmlTeLz+TLeS5SoxD7xevs2YqOwjPBGJQoihHJmRSvDXg5kc91NerY7K
h6ILdMHdxhDApY2voKOI+J32OY4tKNGAzgwL959Nig0eZlWDRe5/EQzZ53/q+Ri0m0NbYfeFpy3M
cGydpE5ZkQ74bwpRYm4OLnsel54brScwVA+XIps7E1VUzScOvcNfIRO/JUcn/wCDNUJAg2Rcc2BI
/0BvOOcnd5J1teHmXR55rW6/9Xv8qhP5eY1K/nQ/wgEpgZUyClW1T8jyrJ+ciNxysZGg/5iwThSy
eWNJS7vTrC4aHb6827dcY6Tvsk3Jiq4wjrKdy3wJi1s3+EVb3DvcOJQ2ybF4ihkccy8lgHdebkAf
HPYBXKoHsPKLzkqAUNpUIcZc0FV5ByyG4JyTMLczk8gMFMYrbz53f9Ywyj/dFNkXukXKh5bt7xKc
YeYbbCBgh10/tIru24GifUP5VfJ4+kvsNMkHSldUtqivXx4n/FAJ+eeIKkuwcM/ciyImqc43YYVO
KvixFne99CNN+RDHSjBESGaKXKA2uD4g+sK4up5lLIt8D6ejHnogPNTGZLFGl0SOTaWqNzICpd82
USImYzekBuH76KgsK+M+OWMml3nCN8FsYNk/DnF8e8DDXkhBXnLjq9FLXf4CqXwhhaRu2/fpuNuu
26QBUEwaRAMz3MYrltM1GkEKv1a6vZia1cT1lwdQFOCv+8CTOjZyQxY/tQ8MY/5O3LVxX+1XUel9
eJLvr2c+nWQEYl8cMa8vMevKWp+aPSpQVLPPbzJhKlfvvZfXg6GlZwBtSw1fSH7fVuSV1MiE7eTg
8jSd6W0nUn5F3gMktIuXkRA4lFVgQkhKu2+Ozh0xJLsc1b7HFhTyYwx+szHisyBq5edVoXxbrC96
58k9jqYqFkuS7vBhGxHvK3Ps2uJ/2qjneMFhFghBiErSeJBoXS577fXwuw4tu5j16xlE0oYR13JD
6TV6fX3kBUhRD6AFtsYkt8NL1PLP4ehJw/F3DzjHlEHSl0s6Y4XGhYeH7QXUz4KUrOxgmajVaFB5
HtEpgHQtIvUjq+/B2tTcrnWAJ1Vl52dJMv5ERx9E+wq0zGTbTyzmY/jeJF+d0qqGRWhOJ8hWF+x1
nRmzvhzEw+NygL/RHRut/nE3fMlHM5dQ++dnSn7j7n0d08FB4vUzGkzawl8GlPxcchCC8FvqZrM0
qjwpfDk7x4/28wHstofA2gBohHa/mbnNq2dr0EQ7ogo008pZB7Do7u5V3e19TMKTyoNpra5nhH9J
vdTNihB1Z3OwhsgP+02xGtlkz8hq9mJ5Fb3DgzA6rtApRjJ1UgasS+UEWcdgfHVwyJzweye9rhx2
S8ImIqILLWn9RocxjOFBYgi1aGiyGPfB7hmaqfgBiQeSHYQ4uSQBb0q6NPCalZDVQslQ6V5CQ6Gs
lYtlEbdjX648JQxacA8VFUv+X/B/48P1v0UD0dCrTf5iFOewJsbm22BFV+nCJXzBOi5RPIoaVP2U
u/MbGqw8ep/18roLwyOeQ+NntpLPzXG7eHVHjYoEifJhTRCkTyvLJfMSssZ6PeBUs9dSLYf+jxAW
CpE5yqZjLNMynFfdTlf3bSsmiGNb0wwEueCUjjYzfeBw3mSPQa1A3+rFyDWViOiFSKJJA06/BOjT
XyGI7joecfjdhwcU8eS3u1rLbNhXyZu4/8lWsEHsJ0cPCUxD9adUuiXiUMP3VEnW+k3VD5R3ZHA2
Zn3tGw4ccZ3F98WothOnCIfU0Ho/n+X7N6JZlK835dON4oLCDnB3Q260pZn+CA/ZyXGwnzXH/MIM
3SpvmfO+I1/UIyROJD9bzESx9ynx5gkV/3QOxw5juw1VuK1i6F7G4ajQquWk1sbTZb3SM2/ObvLr
w3OK45RNX1S7D23/K74WrJjUVo7jWjRAoNrkCMJHPWtEdj1mSwPYMFWs15nEVPV4jgi4x97on5ke
Us3+K+nzUBG+Rk1yBUAMC32ZVRIXF6rh7AXSudmNDEH6nyyQtgQH72GLoqMTrktePULvqFdl5DO2
+ii/9g/VoAmvm9iKiLpPT5T+wtuMy96GLFw/eKQmazR+ZlhFNXKmD2QH7e08odunFL/3+wOKi8Mp
8ufalV7LVk6iTmMEJ2PeVW5uA1jxi5SO+3iayyFtYO8a/9foyD/EAyvdN5NPuY0Hnvay4FV/Nu2I
QE5XXuREX8bDsXSdJYFOmwDtw4jimyHo6quMbT2MSJ//TSD590dODPm+UF4pO47tSQcjQGcz5R19
3cKCsUsQj8Ys+SE2oBiJZHe+3UJNuVyyq3Jcv+yF+H6wk9u0M0zDvnq7jW5VWq81vlNwtWfOUKS2
cLxkYQnFMi223hFAaJs+OHP0zRm/sQJtL7Eo6/+w4ML0zh2y24dO0NJa+Et/0DXkn5mmBuLxnih3
B7LjLxjNDlWXrgRPJhbaZN6b5hPeLJ3tqWokNLhahM6i847p1uCG34VHNqSYn2pl4qWklxhPulVJ
j3bJg8/DKYsvhIBw8qAsncbBsLWWSbvg5tr4TH+6i2NhrBf15E/p5tr2QqXd/wOLyGaAfzxO+Prm
cQsKJ/OdtiZsHZQhniD6mTBXXgpmP2cqul9Flx/EXTFHT/RGV7AdArgmHzhsnGIp8CjPxG1o/hh3
LoqOWhF7rAoJAvZhCxcoscgU2pbw7267ONYkzv/Rjr6MOEsNX+wZBFuBdYl6gE9H2M5+SF557q+w
8S3oc0I/IETc2G3b1rz9fuI1Gbb2DrIty/6T31knaye/s+boy09plD2QVrkAUVLFQPvblwE+QuJ7
UXw4r8U1OUAQaUpWNK/gvl58IvS+zAZPqrj2g7EVcuh+o8F6XIWJsz5yrrOTnLEFgigIuYBXzQsH
tq7YaKmf+mMlX2XpTIkSVBhPWRFuUgRfuzPcKKOFEoygG0Y05ul5WtAFXhOsDAIhKwIYSRc7lxLL
tRSxP9UqzPtoYntZKQbBB7arU/yuM5+jI94+J/bUsDP36hTV6Kar2xJQsBKW+EWuhyWJb/daTI1U
pHmZbRwXGDiWDZP8ViagZc72urg3nbtj8jvWToQRU3PMhaas6dWCbeEWJKN0sl3nkIH5PH8W0NlW
rSrejKHMsWcRpZl60MIjVWdo/Jr3bUxe8MXatQoiUAx5DCnxe193XwdWkN6sxtvSOlpj/ObVxrQY
RhkAqEnL6L+JV+Z+VQswvF+LEjG7/QUfFDRkvLf7OutLNrUz9jLEmbrEipHvgLwA+4RrKh0JRD3L
PAe8UmLIUxtwaTQy/EmbQFSYPyUQTwSHCmPxC0tvpYz288q7vK4MQz5FtgYXtJrSE17pcHPOCM9t
ksX26TVV2ut/Nxy4M4245JNRbDsJBpLis5y+cIeQeXxte0Ei0ULz3xJPx9IP6ldqNjLv4M4YV5zj
yJYbGaetr2hnR735HBg/avkB9B4aQIpcWdJI/HqK/zFKe3bhb5o2ZzufuFp8mxoLJiQ9G40yk3Pu
BU7TPRXD0DwVRLiZFjCER5qXQaSmGLz8cSOk0V+IGvo0qYv3OZFH4UDz762x1d91q5/AdgcdH8OS
qoP8haXW16UKpv4BNnEU5atZHqiPg3GGGcjdrQa5oQ3bXgFQ1W6iOS1Gq2EIfM8pLsFc93VUQf/S
f9xR01rj8M7XWEVgci60W1MWpt6qFfmg11ZENlxLfwI9JImDXEHpkGv1FkL7gkSjQkJj/9LykORV
JJbATaBSMCp+uDD8DJyGFeTDWvGMZYFRI3VKSAHAgyN9EZxb5bvCw50bItMeNSKqqwE9Q+jvxJoi
qHquuxIHIlR8WPHvfX1Djc6lQ60z4TxeMJVVxw0awCdEq+/tEFaSFRnt9cXgk0VgC8FvA0mrIN2I
Ex1WBWGCIEOs7YSa2LKqrpnMxIW2dIaKVhpDNNGTp26qVFvMv2P7irETCn4k3TMGZNw6h6VQW+UH
zYOgNr+cweEyDn7HY9cjEE1hkEYOSxh+kz/F9BwZ8vsSdanLk4xdYw6B7jPIeHKn0InIZP/GuuJ8
KUX0j4EhOrYM2SM4xQ6VKfvmZAc1Z3DHh4CNItGnt4xuel4NEcici6ABXKPeNeBcUoh/7zCwhpqC
1ZJ0eZzj4NiGAMCvrS1ZVV5stKx1Jzjn5IMpar+OCwDlzA9IOV7LJLvxjM37PtSvFmhHn92ZwDdj
VQTt3d3lfWXOx/IMx/KOZDCXOCeCPvyQuOLeRgaPvg8rkIz/ecp2aKucgwR5AeIxhH6WvceQS3yo
wGD41lleiuvjjPcEX/6gGRJmP4/WM0ngL3HKpcVWeh36t+QjCF/uX86+yyTYVwpFfrbbtYlqe76G
fki3OzpCjANwa6zODcMNPPYeUn36JmPIPOhVLn09ZEXnBuk6mlcbcGJruPn4td6WhY0EzwBQBS0x
n1itfmIpzmRGp8UPVnKNBzFyf6DTzFgW14FD++P+aVHhMWCOHFRZ/RYfSHxQ69QVn+7HS9sPq3yc
Uf4TFkI6VHE8AqEtbJEhEy8ILQme6Jk/GeJnk/bzUFeCioXVPpgnvqNAmtzgBTnU8WftbCgg8PoE
63e6Z2vzf72GtZpEhe/wAqCbYHtitM3cqc2s4ixRDmFqXICOj9Ycgv+pLgpCrUABDg/15DCpT/4b
iGCU1Yyq1IrtQ1ELuORZ5H+J7nqjR5au2ZsYE/5YQo2L13TC2c9L4TrawVYeD1OISCm5BiGHnZbs
bmsdObLrh4wjLQV8P67qJZtS+GTp4z4dDDqTxDGaVyNTwhsrn3d2YmAgRkzGh0hv0PqbiI3ilrWs
opgi3lvTv274W5FLcQPrZRBw2fFsCEwvSTmj7H+fZs7pxzDtFOTIJWHS/l6yuLsAehtCqM8KHKsi
ZKm9g1S5tnaSNQHP+7/Ai836ahJvmnHv3Bqt/yxXjf/AN7k9UNy5sg/DZJCdF7mKC4Qa7keq1Qoq
gCFq++gv8I940W/75Tz7zKUpflWjPoWl0ZwF7pX+LLBPggADYDmTRr6HqUlJaTNwN2p3fqjTuLO0
eCTW6v6ZmrL0WJFlMCZF68oiAzSRKyVMnRNHxXG4J58LmnYaSYxtnLmhm10+AFFCZAmlcwsihcWY
Ds57dczTNoBHdwDWSV/Qic4jkd2u3j1jMLsJXXY5NLjeUq+GAxYaEvJZlyOngewG4pYOAUc/FGin
SgHP5hj9dQBG/zjjZEF+qkRxlVgJyFiGMEYVlxQmHIjoYaoLNLnY5JHziQnued8aEgvHt5rfGqwp
1XTlS0apz2ajzNFOLGLQTtBrjmy0goV8C8mF32Gyq+h844mbWy/R+Q+x3J0aFSkIg/cdB6Ju0tgr
dBRCg+CwdtDF5gfjuu8lk5tcGDaM7xfdF8Nk2N4lYuffb33I+As+n4616LWqa8i98m9Jr1BU/meV
vwoVxhvzlA5l+ILdnLiBsXPTFj0cfZGCDrsb8Avq6BoPEdS7qY5mrPCUsZfsLYRo3kqIkJP7X9oi
v6MTv19Gj6UnWIbdyMO0REUfaWnJEwv/O3tfphEenyZKwm6XZNvxfo7xyxzpajwsO/UYMkSSxIRx
tWY1NohIHjL+IfnIRcnxP5P/66U3AhdqLGwgx8GyeNYu//P9eAohjp3rrszs1ahcqE2OJAbLJl4+
vfNKnkjsVhAFEqKsHLMZVrlXeed+MFpFqnGmrRGGtXlrh1UU8dzDB0GgbA4S7h8LO6kifweEl1bq
VemYz5e0LFNKGz+JieSxgncRLA1vvEvo1FWVJxK6BWAaQiq080S2NRfWmRlpx3rzM9kdHH8eAypN
OwmHCJarg0c5lr/vnmaEBcZ5XnOy8Brn5J0LcjtZO177mx4QJt0gW4H7PP2lsxa39OgRNrUXkNF+
Hc5xd7k5aRx83Vi/3MKM8w7Mb1FnUSvk7pPSfsxZNufcXBRLaovwWt4sZuLChFlG2f1Rlqj1YpyE
bkdmYfuAvA7Q6qiPXWwkrk/N4/wtiTmGvg+q5+Vb+TlY1pGKZ/fME0C6m+4f+flhxWIYjQEPuv5x
LzgT1pJzYejZsBMuPxpOX1K14xDkz2Jzw7JtqBPaS5BADbz2UY+E8SYW4Z5U7InzWPFXPTTOJb+r
JegVYwCoKaX6ymsDZOdC5plSl0o7if91wx74X7yZZ44ILC3khxo1I0AKudAdt6Er3dg6J5QP9kay
9bOpGFtM/tyvxPZu8pKA/NkKTsr5YRTrRDtmZxhKm63BB4MXJ19sl+jnjanWWabXND8JnIhpU3u2
RjylguxN68MiXsjX+h4OQXrKq0qPhVhVROmacUlwt3bVc9YjjoKbq3nRj85Hn1i06VCxL2BR1zN4
IJtAEQypxGc9rhu4NMqdyujiXMqurP00BiFIFAHZPVG2GeUr2legyHx1gyz0H6p469Ecwb9rm/Re
xNY9eUHhmuMbm21pnDsQy9sMg8NfP6Xwg+ivO+KT1h2N0z+sc8Sh8Fqof3aSvkmL8xvxAKS+vxh2
FQmXmSeAX3DEVDfomUUqX6It5zFArNrbGb/eEf0+QUpAgY8AJalWBTZoFNM6ohe7ofGrA42ClSDq
GoB+ymMxvujEwSW8psS2KZZVkGZbmDCbt6hqUGbvlW2gAtl6NgtjO5GBZ1tue/abgb78hPhLkpwj
hJjAqLJsUlKr7K8WfXGgIpYAbO6/x9SzrW96iplHQ715Jf6DPHuHOW95HeSCWZ9mcb4i9W2zOuqW
5ylL6LsG+dTJB7G003Bh03uo8SbS/MCmBpLE1f66VekiuVux+wtvrWXldO5San3/fnmGQuMpa2wa
NFqN80mVAVSo/w4jTtuFgwkuWl+IhvPyW216VIoIKVHOaICFY8k2EXbVYbNToO1CuNzUYMH+5Bxi
8qoc7mYk+enqDwcRbez+K7uHEY/UtqPgtZAP6zRgu2YC+/VKz20DZBrpnJwiQFklSHnq5EbvpBPW
+Ggd2eUo6B/LWtBOqg5zNcs7ki9Y4L+HxBRACe17OydtcohGzQwUb88y2j1acDWwQ3r2TbSEUtlU
u77icCsS0FazppUHfFtz3IMOpbMVaV7fJa0oMAFMjnjYb9JCttnZzBTjhKenkyZWoZqEew+KeLfL
mz2PIURBNtF+auY/cA6q7EHf0x76qovnRM2jyRY5ZS2Ie6NSx89Fy/94PKiHJYQ/6yX1h0nND4SZ
+oqkY943pBo/nYPrJs9dWankkXAlzFQd90gRQzoYqiKPo+R9JYgaGPjtPLF99ZUknqD/SGufJN3D
YTetnqbbf9Mda+NMyAXrunpfxrhc0xM4c7NFV+79OT1+LidK3gAcabeGH3MIWFdrRgCyuGXd8Mjp
XkhQ+h8HO2x3mX33c5v8sHNZFc2YxLm8QWHkiO3TLIuTRlHCtqauWuVyyrsjpgTm4Vk2soqz+eu2
os6iQppvvwKrRc34Ux3SDYa4CRTykmssg7SYQStVeXLxAS0WlJsTPp/3EuEKZ6sqM+R+r5LJYP8R
CFN8z2MgKNqayLvxswWXaTShX8pvOOUHMQB5QBheGsB9jONuStlNI3X87JLcNkAgS98wENBmLys2
VmitoEXG5uGFrOCBQSR+e1Ww7bbctpcdVkrtTb331dsePNc5AmvsPLBfBZyZi8yMPWf4TWnuvTPz
fdXNvW8nZ/Ddf0Jp9gOfb8OAwoQR84QVYkAKprRuXx/39Gh3QaIGIDWcSoWYJTBKfWzj/9BOfOpG
sdby67jCfWHobZKmkLTjd3QAXpukMRT+a3Q9P4D55eCoBbB1fpU3o8LIqkCSgfEtOwgEpv6THp+2
tyiOhptvuwyimeGGktHsWo5qmVd9OJ86u5jZUotpWR2ywlJx9pjzj1KaOi4/hYWJouwIyriW/ZOv
0ThrKmXAMHvcFIM2cB0QN+clXIJrpTEN2gXFrMZV7FOk2w2XhUBiKCRQ7miFCriVVUCtwC5FS0BI
ZGxMoFYNjeWgX/znirhDsfpIYsGXRk5/6VdsWBAG9mSZqnEVHrQMEN0HTOHI7ZZwVw75HL1yfIBf
CB4TNzX3fvnsmvdBoxmz8i53SWm4cJ/+QeCU7Yra3BEHub7JH57gljjhdUPqLpmqhSMv1IhW4PHU
vpjgF10vAmtjY1iwMuQFtzcMBLTCBwbk+Q1MOpIe/38BBlOV2CoiOTfiMeAFDkKsfD6fC6u9lQ81
eEx/QKqlFr42p8ehAVLOxF6RLQOFYjV6BcWRMb7ez68fijlGulst5MIFIYsIa/tP0j5z6RQrwCT+
6mfW7RzhqnRcb6FZ0LO/2UFrJybAeLp3zihMq+/IBcbR+pwgD+lih6efZNcXNETS3VHfRsJlA1sc
/ToQyGtcTf9VrEg3Nkv2cy81QyLBilroxK/xG7Jc1iCUEFqpVU/b0ktYh6zzDFhZpoJ0Q7eoN9H9
XkC71MjrjXU4kEQfTyO9nVNib4FqpCnFjAS4v2XV+yCWFT7wvJF6oRCDy1YdON2Mm1ALDeVPvbZi
YKz/En87DcqemtsNSbi00PC/y6CcURGurRdIFt8SZU56YuoZ9OA/H7Mkr5tgNWVePvHbkBURwDyG
RtlzfvCx+C7QbI2PaR+Tj+bLvaz/rsrGYoSG3AuMIG3iKAQN1TNtJQoY5c+7wo2k/BoqXSh/7Xq1
mYlStVzMiJCgDUBX3CkRIwK6vGwIoGCO1qv8e2BGN213hQtWfDmZfFd92AuZCm6kevJ/sjre2nE7
b50MMwxKj5cUus0IeIHoAd/hlNMeq3xbmceV+RJce5/H/Sxk6KDIWtzN2R+KBayXj42BNAgXw7BD
v7DhH5i9XnP9q5Do44HucSPgZ8Nt+dfljWVc+3Kg5Yfw0YSPpKCaXLRvBJbARZqeY26lWkiyr68E
DQQ3/ukBMtmVuqjR8W2aGM/szyS/w5B08V/80z28933oIgJ2aTFLJbtDgZXX2XJ+2n9O04mBHPCd
Y36LjNfKtbSOurESkBkBQ3mD7veVJ1r0o+KNlQWiBDIRFKVs5ObCGFQxcQ43h1t1P37BcK5Ju3wk
Sju88ErkfOdw+lZ9R8mArMhwqh1OKIHieUoLCXBU+hxS/GoNn9fEsVjhQYzejNMUo8EKozsb+Gpi
RCpEtpNMt786s6Os/OOxJ0Au6pR4CCMmnB+lP2YzYM6pwAF87UelkYl1zBg8rUccF8+yOqF9827i
xRPl/1L5yWAU8KYO+eOMC5prnpd4c6WhBzWNjdO1CwjWEq/fRU3F0IIQXl5g11BmfLxXcmTdrIqV
omc6060l2ikYKaKGOkl6Y1ZmglvdJ0ylo3npn+J45d8lsGXKDNMkExYKekhHslhAfSWrijXwqZlL
q/Vn72NDNIud5YzxGy/rJMipGhPIJMzSuxrnxslPF2PIZ4ayTyqjarzGntH4Zh9hty0D4GqCPTYg
Gh/OnB4tyKlK8nbxRAnfXGaT9HQD1fJv8A1MEAzR2V+Dou4angCTJZwl4rb/dvUwdCXvb0Efb+ZI
A7Ap6lildGu9kMGrdcMBnTPDg6wecB7D23fPWKm2zVfHvg3iqUlaDb5iiTNhRX15aqIMAAXX1v1O
j2JRVnGCCTBMigoIonyW69gPJy09HVudH1RmdivOOHQaBhe+zS5Ex4HGeVflb+snHim+mMlvZuKG
FrWFolWqimOdVbdq08VZvyFlppt601WGZLSe5p4eaUOjecgbHYZNEVKC1WOrAaIUkt/zSFhos/7D
wR1Egnohg2EWrJtcZHr7Yyjq+A87xTkDHd1I/ax/PQW1dlfje6IvzFrAC0yjh3lVNrMyPVBBOZGF
A5X/U9kE8IVBnUUbD20GPIJIQ+mpuoGRMYhtoJQ5daq0y5SpKFG9R6OkXMjT+iLNlILHMdjdUcmp
U/07Sa+r0hpB5xgH6MnaIHKxdUgILKgdCDF+tnz8HoxVDoauS4iPVPF2vFfJYhCdCw09LgtrxI3l
1rpNfrVfm5mSomFsca5YrlE1g+T3v0d9UKKFuFmw6NdWAlwu0rj5NDqtbSzcwoLvc32WSBCrhHva
z+jEd0EL0iyV/DGNEwfmNhHPLC+bH+a3Xrj0AChcVG+jU2wScSqa0j1HVyi68QHDUMjPKAuHiaGa
KTVcc+N1+xp6xOLJLADDfXno0QsR5NBkjYjRI0bXNtO/ofvXECgDCVCJoARl2t5+HSWL7pTWKg/p
khF/uIk1RtWAsl/DeuMYvK6lUoMRW0srLrBG5D1QMQw2rWVrXdiIS9AiYqsxcTlyukO8rD3y0l0h
/taWY429wT63gBdpzrRGt8du10JJccXCzINTdnZOAUWNMynBdcKoZ4IsZ0ev2UvCQ7B0lEPqVeVT
fUjx0gBKBftKUSO/uKehkwMo3AWkTLoin2c35yrgBrcErolma2op1P+Q4t8cXQ7U/6xAKMZZhXLi
m4vIKla2RSnqSP0nYDuKpar/msSjA0PQPgJw4V1USQm5doUkuEUXCDXLIQ51Y90J3O36l1lT+PYA
vrWXgiPWOv4MTPWT/S/Dz3XwLkLRq8M+js7YKNQsHNfhRjzFV+5RSTLtAr5C9xH0DhSGZFR7BbiB
JeASYzwugreZftFEXS/5sDBQI+pyY/YXo7puWvGokx7qC47uF4S+KsxZV5rOo+I7D3lu00zbXzAq
/Z8qpB+MjJFUQT+MoG99/oVH1t8PI3Le+tPrifGozFmdJoBuFVwNhAqCSo152reJQ/0/W51QU6Y8
MSWpMkgfqr9Z+UiIjWPSCwpUi7MZVvDu0GFAIbHcZi3NWQDeOYP6AuUEb3BgpBheIkcuHqv5SQuR
kOgtya9gbCkACrjhTM48V230pfvSJ3Mzv/pvs0imP9MonwwL/zyHRTBbl8LcQhGM19PgVFjtqoX/
ksXChq3EvrpUCjZiuWT6ykCHUQkQEPpFefEijDLeyfvnMF8mnn0Tn5jQNKu+nEAe5oklzLs0BGha
OffGBMAFuoTCk9UBrDWdzncNO0OBM6px9f3sTffudJJo+HgC7YcFUrC+sO0bUCZJYFL2bxm3UVAO
6uvDj3zU+Jzvv+mCcICOw5DWyoJiPFnAAg4eHpc59GKyokLpc7tyPQBH2ecLWdme0wycdffLAjrp
JrlYPti8HkAt56gL/Xu2dM+fKQQkqTiLHniDc0Z0mTk+m5tuAaoapXyRAfgq60hxtSEZDifiyJVr
IEi5R69hTSkEWO3J689hf/6Jzdp/U97dif0eeJ08fa2bBTrOWwsc0jO0I5txh11YfAvJk96S2i8j
sAFjYnsbeETdSX5F3sRekinlqckKzcEAe9/mMiDDmsLZD6bHAEFnxP7SzgQKidY5DudyZaBCsCyl
biSFnaY9bk8U+mGbBFeX0//0ibzE8UDR5liuS1SwLXQBwosmEm0sW/eD1+pmGDTT6R4a5IXq1080
ec9yPtDvbKGTl9UCwZOtElKj/5HeL9x5b3NswksdkIMNHAb1Ou5g3dSjq5TKkgqPpeIGk8FZgYZe
PVJH04fG2WiyNkCueOO89IAFOKUDnrAU1+Iy8hsvNwSxY2Y+EY9yF71FlkG2egh4aoyFMjYom31B
ubYOwQiPov2wNCY5e9P6H82A/vbXFX3/R6h+uB+DXf7VSSTN7sSwqoDc+iO9XLcbCGBTs9Y4mAiv
oEfzTpWG3Oe/Uxvv/XM6f1peAb563NDMbFhtxrqiVgilXegeAXBLyciRDZbJt+3pnR8cdsMG7/Cu
kpBEKqdQgs6tf6spyEY6NHBBHlhwgaj+IBxM3JdRjnu2Bemzk0qle7C1C0GlN2qVP9FmorGobH7j
oW869tyHng4KedeSAc0wWrM24LWpZHFf6wbzi3pHBjPDfUZeYFbocTlzaINcceEYJnmb54TfKTm1
DLRqmMpVH7V+3iXaKmTa/buiG1Ye4yUE0YhiTEqnSE0G8e5XdzbWYz2YPyaNSxO2RvApJ9B42iLi
flfWXSuFhtLZJ5e5cabApLQ2scN6I4QuKr5VW4blOBK2mKbIL/0IEXzGGIzezRHfa0iRFBIyoU3k
1zSr//eSjwl1mOOzqnpXY5gFZPAN0hBN/IU4QcBy/bg+3rILNsdXdr4R5sUtsrbuN219DX/2ZbK+
jaUjBJYVJhZN4LRi7ohTvWyHzjtHSgWyS8aOj4Pbv70FMJEAgpi+qnRZt6+Uv07epwkVUf2GZVX3
J9lHMgL4l9iR2Edr/Hee2mXnQlHDJXYy6Cw/EikZkXCAZ8g3iFbcZ0Qr+K+8pud0BRn2bNbl/MoL
REswyrS+cdA0xNxQiPz2xMQNXD02rV3PADyn2RkZcgi8XyOJq9XRblYC44LaM6jrmnQcMCcBLTWp
EUKQfSPP8fl0wyebNk5iTorJQOXJDhQczoyFlPUDq7NbwHP8w3WfB99OQRGsZTws+HmvKg0g42On
zNrnLg9U2ecyTL3B7DmZD5a0elxFoJNQXi/q8bCgCtIIc5tel3MJMHpcs3RqgJSeSJOyE9T+zRfe
aiJ7yJs7/+Yias2cELQpW9mnhSwE89uZepcdMNhte34deIPYNk5OJvD5lZwiwMHEjRm6q3etUhbm
0JHpKeLTdMLp+rlg+hJ7XHXrUrrRv6z5+XYmeNx9vTTUJ/DCH9kRPX1XK8ZjphIfLjqPzAN02isu
q+X6mP/ht2CTJEcxC3LRTuANeFk8na3J6wRGXSG2lFOL8Y0xWosapEWWokWl+pczeqO1+yA0/u4B
HFkxjM5qgTNTQrPNaB3RUkGPgmxD4GxqRJZut53UZ/u+iLO7ChB2AkPu7RF5Ma95wtBdxjz2Jv4V
Ct5nPFm2GKheXw+sFVNmBmtveMjQnAHsJlvdh0fVZfEzno9VUPyrC4YQbkOMGOk+0frlmCO+3S1l
Kqvy7Lgbso5GYo4dCBKTlCdvQUCKok/xoAq6wBVAV72Pz1dc4hQ+FhLlchel+xwcNgBYeqEUw4Ct
N0hCil9Gn4o14ZuwWBuj+thkc1ABpmaorqbiuNTZJO5q2nhrtpFdKOclM+INNetsKim3Tz7p0uF/
of/EIfsZVtfdbhwFWOmpnn9B9gyaVmI+ckZOVjgiASO5HV2I95XfLERccBjOO3VTSqrXfhdbOmPH
jpr0eAv0wNuwGfUCjLv13g85e1EnpMUZtVs9xT+hVPE2C9OaU+W0I5XRSJtC+rcN30LsX0PVeFhs
Pry6ctWVCVcdOWLQw37D162F7AKy3TOYCDKBUMiv+zoGvARj2oDxijDFoBOBM2y5b1OP80Nn+aA+
ftepSZ18GbmPhFOitTw0A6It7PZEoyavSdKf9vySeqGBLjy7pXglkTuaWPAJHi7LEY+EIvci3EPe
hjRJ0A7a+SXXyhqwuSviKuD1NCyGi60n6dw7PqSHsZvyrgHJ/ASdFJsZgkAMa2I3K82AafxialOi
Jc2BgiHWee7VHWFs/f54Wsv1+EVGGqP9D4joYVLGanHRtt3acMUYyOYVfJA4hGky9SstsPdkEClx
YMEPNcUOPR27NLC3wqLD+rRent5LY/jaLydUEwLqbe068KNMnL7/wj/8wLcTr9/dxjD79DBk9pk3
NxxtC/rsfTB8nGdwXcYvnf/p1ii4/27u7X/AO7zmw7xI2haPSxQhgJfIZL9YykMPlrK192GEQ6vQ
INEIWvj69o5vAeuwgT+0cqJ7W8i/zOy6BYO5KVOfuTFChdVcmTqp1uk9AlSZe0lKgBjXx5ZWX087
uN4AMSABhLe69TPsahY+f7s6HtTPj8GxbgSlgiCkP916R52kwkycZkfukgWjkhmHdUePgL7kYcoK
zszK1UAUOPlJ6CfOa89VX45ILgM9aP7iciLTYL/tQzMirqhQOnhZ4P0jUKMTgl4TR7cW1tO/gh/F
mXqE5MjkV76137+qwfoI4OFImAhSjDG7ozrXELkRXCTSU/Z128bHoscUW5iWOYkcf5O5IZ7wrRjg
OzxJBuly4dgWb4i6TmKU6bxAHt8/1S5GTXhxAwmtq5GvEiaWyvhXNrEAzomwm5RvTIlZNwIv//ZR
DHCcb0wFKSuYN1ebo73kXyJ3Tq6WFugKUi60eiVxQa9k6IgVnH+JvjIXVErUVEcD8JdGNYCy8+Vo
eR4S8NPEDfgOm7D3ewu+UnLhf+C6GFs5DvdNZxYTcQwADBLu37TAvlIG1ZC7iuGS2cYouBt3cM3E
w3yQ3efljBVXa1i7LGtKibxOGanlGNXeC0g0DRB695mK4TxvPLw07BvIb6t7NeKJaU+3GJvs+s7b
ppy8qhojhiW7myfBfYrWI6swXpFWLUxnj8lSKGbJdMQTo9gQoQZFeaKMWPptvAfpnn7b78YFcMVu
RvEMqDZBWvMuvgx5Fv3jRVemGYbCQuDUzwRREhXdXgpDlINmJ7Cl6qyA4BupsAEJfdSqlPoSBStM
QQchAwLqvf5Q2WH30x7G0QyPFpT/9og5m95zdB0cByAIB04nD46cGGET0StRyL0OVauNRNI6bcHY
P6ACDGbhwBR6WGzY2REWr5IqkKNgChWmyWSVVJGFtvF4vJ7SIA9nk9sTESvcUOAy6MeMWPdNU5I+
gsYI2gYy/m42elYV5Xo8k8JecO/9Y9g4Y3VoJdCwMlRO3nb3lmV5jACs6R9+iofxgvrb2ReEyZ9C
9QGIFmZ8onH4vQadJKn7WSFX2V46sowecsIjbh43Pp/0UvLuYzzQ2O4U9w+fx6wPALXpY2aiv3Fi
dd1mU/DlnGR8bYLVFXZuyckQFWNsyengJEDnczxdoqhZBFA6x5DLxp6tKi3RzUPOUoqSnIKWt7f7
Yc/D2GSXvrzvnUCVFKtGNCEHQ0HnZNLjEZzLCMROA7ooTYrDhxhmZ1AUI596in9+O8C9xvlGDXQ5
FgVVAQp94smiNMc4ahFEVtcAAc/4rJrgbH0jtcnbcmrOjhWJMcHDEKhDvb2FQM/OGZhwmvyt+O65
f9sqgiu2YVA35LYAhiz3AQJLwFLwm8mxQFajEh20yvCL4hh9e3rSgU8PN/JxEM7kkI474LLWzBbv
oLw7v4heQqPI5dDiipuLFy5OjMJS07O8d+hrVwZzTJ6BUlcdO2pT64FjAHRExz2Olwt2plyjBLGP
BoHPOS2wpLeGQ82tcsnRwHZE/w3P6X++qTs68f6PnOVDRcfFs14ZcDHcjJmd7l5SFYW8iaMN8Cwo
Ucdk95Peh7rdjtl65j0R4L7IEmtxHqijiVfeibqJCkegBVnKB65V4ff6RaZR6jWG6/d41awN3tKx
tjw7g7PVYF1SctwzHJ2HuMcai0YjpNUbabqmEHiBa3JrPJYE/2DYfcLIAyX95ZPoM9WaVCzd2UYQ
yABXWwnRNSucD0Ubl9B4ZOzEUrk729SCacIpgtBjxnZITI9yqQJJoRiyjja70oWATaQelOfu8Mx0
Sn58sXJl0Nobnkrctt0qZaVOr5B79soveE8JXtGFOV9JkKxFU8PYzTPyOdxwEGiB2mJYmuKPijIp
6H/l3mZz0zyhDaoB4r+r8UPN7X+kQvkUlowZgcOQlWjGQFQ0QiQt5fLRB1eiJCP0d+zOH/npzov4
oDb9G/W1bfJHV7dWb0kh3k0VIQBUVK2IhXrem0b6Ux8hgHHTT8H9iWnA6ZyZNHOtXOxlTr1TymHq
c8pa6/ue5EBrSWs/xiNlOfuUEYxmNSjmjWtJ859finMuDTf22AW8kwfyAE8p4ZDwLKBXOMVwCy6p
yyUtQ6FHuQXC2Ls0gAc7td7mi8u6JCOaemSe4J+amVJKi0QjAO8+IXZNpAWm1d+V7q+wawpiGdx3
J4BY8JQlwrpjKtwom+bxjaFRIEyltodzyrrL91URINDrHF5CaxNF+4jbnk7PIIjgf7Qm89pSHI8n
R1AH75mffJqZfBCTTv/Rt5FFNg+hSAmgnNOtPW4AsI90QMQHHburlbPowHAHNFLaNSx1zqR/noZQ
kgupRCcfpt7It7ooR5rIMQLq51FIZQumwj3oZfDHTdSG26UpVNHUdtn+NtI1h/OlqsNX3mERgCXT
EhwzG0ztQJIpXNXYqZsZcnWwNvb6+wKthQJGG4k40Hv4jJYCiHHo5a/Ko5dW/4PzcMqnYb6vY5CB
3VKWyzD+bG+rovdJsaOFcisgGA4UOuJcoK8uo2QYdLWVXicEB1Hbmrz8Y6w2NQh+66YylwhDjmkH
QNglQv1SYlrSo3XyA+SKAlDPI5Ph2U+dRUKsIF+pAl7DYFpZWoC13/wY7lQUDVenb1bmb5MzEll2
9rH2CHDtjtfLX1tJkStOFAIuYhEOeTPf05YKmCkoBrIHNJLngVoTRgbfHoYwEsmWugl3Sv+1eCt7
hXlZ3ut29A8jPg3ybYi7lPLsuYm7gIRW49s+B1B2IOeIvDFWFIdc0MLqKhM7h8klyWdT6WGtA44C
jpaAd0rfoFuhyLxGikwRnzGSUnYpZG+XeuNjkmSW0iVBKFMBUTEvLKpos7uq87y2cV8rGeRpWTTr
BAwxmCSR+nzfu4ALFZB4bUknrudMO6Iud7N1khjrFf+X7F4870/W6weXis6+nVxeHDIKkMpJ0he2
D67q3aYKBoSpbeE8l/8MYdWe32HnwWGo3T/wajeQ5e7sID27gU/1eDyYrLKwrqUF6Fzsj2ErYciU
xDTORTR/iWnfuMiC2si7r9ehkg+x5ygD9x0haWr94TTAZO4PcKZLmdMqBG1mo8fogkJ72ZIsgmqf
rsgekxNGhhhp+KJFJzt/r1iq5CkZQiQtC9eQTplRdlNO5TEjmWhHzAa0wMaY/L071tqy8pB9BWsk
yw/bZQKzzQdA+u+vvWtifVOvISRPfQWpYg4G+4VJEfqieDTplTfVbA9enHQUgSSrpZEUkY4aqlDq
b1/y/PKp6uoMS8R7BjdsNgTD5QqtZMrVaSvab0pG6xeXDLcYhviiUFWJg5xnteys9O+/l70YNsrH
oz3gGw/F+bwp48P2Rn7pm95W+E7eT+t9dfUWPuulAIhvSnZ113w9QTEVstakQm2OwZG3vqhvA/8D
fVG7HXwGEoyUf85adCzC8iK8IXBOtK5XY+Ev9xsmXPt3No2a8y9FL0OEu7tNm6sLxDZcIb9d8MAi
efEaoY1B2Tm+Y2z2JuPCTdtZ8MRiSjeNmqVjxFg1kpoK8pk/1PyJVU2YWVawdHEtkjqEJJqSLlNB
EGoDqlg5dgKTLz8OgqHsahx2sYtum6eRxAZ08PDYGx8QlPJ8I571Meup8cKXumbvfbneAJ69/0J5
DV0ovWTIe5sGgsONbUH/qrTIIzOcjuZSx7IU4hmC5T1x5LTpADDuFwGnGJpKzn1b8YaBSm194p6r
NslMpBhcUlvREfu1NMtXybR1R8EE+BAfJvMHbMF40BnMezQLTVyWwuYRMxOhZ7iuo458FzLLAdYe
O30zrxrcajBJcpvk07B7+kvpBHlC9Pv7t1P0FKgwM5Fp9jL5gclOVdG5Je+XCnN0V5ONO+U0AQ16
bUzRm5wONlAqymdy3Lo7XZq6+C99cdQvRaPj3xcgIjKvtOh4tpXKV2iVN4lkmD2E4RqtRrBEmrA6
yM1vg/8dIbl+bWnVBiaWGxUHaaFpNZzyD38puNjw4xgv/eP6yo0KwwiwXle4FjSTBCChoYEEpvVy
MwFnUWhxf16VvAPvX5/jllcM1Vusrv3k7GiI3cHjGz6dbXVHkdyvy4+4nufgTBoXHlVEepkBhgQn
mH2cAyUSxr2qfY8rUkT5gC2n0uaaVhDHlaQKFQcMTX7K2evBSnGZLCZLqirlIuA/I8s0JpzI/Kyw
uE85hZE7kNhRCqBA6fO0HA3swKACu+LzzpTno7Sw5wKhDON+BFzdJWd4RWgmkMx2/0NdaKjzF6JI
SDEfNxdyB9vjCMfuCAUE1Ks+TXb1e6gbKJvCCxDkjCU6CJ/0DyjSPzNkWHomif+/+RQiSedPJpEG
H2aYIUvdegM5s7axMF1kgAmhEraiMd7pqYhy9SLEP87Q/LqaQ6Jp1J4B/2lPsO+B0hZK9nFv/Xvf
ZNwOh2MNaz2Qe8hSDxhCgtXiSWU5Km4G4kk6MOluXnA9fli1P2DXV0/d3nzRs/Qlj9kUglh5Ol24
cycOzzoDPoljzcydIwKhzmBQQs/xUvPczUsaNtKu0Ff9f6cKH6QT+hs7+KareFWNQHJ8iUMB0A/F
RY2J5U0WvJUjQmvSJovyMPiiNxoeEi9yhG7AOcSAw1mu+A6OTrsSYYzWF+16rO2DOn6p5kmlMn4x
5DsThEHEuZeMGUMUrJEFpp8KwfsBkLqmNrw7OedaYXgEW+T05w6pyzCX7c6IfHMJVYl97ZiEGkTg
X7+t9I4tVx7HKOYkFSFXRzVviCz1mi+vzbJvriYFcSEtAgqlcN4sC/KBB7xXrHrdv/jEIXr2Vh44
DffcYjg3juBA8FmDsyWThNMUrIoEIUyPAhJAaigoStzbr0f02kjJg9MviB9hvHy6wMXzHDUsUEFK
Vq1iBb9aLapSlsGLvXFxkjsHOW3S7QcEUFKKn33S7f7gK4sWMGPBa3Vh6xuqbZETsjNS2VZ1hu3H
/Kk7SCGr8JO7WpUhBTUbFCA+KLBmIB23bouoCm8kV/QcZ/trdaVaOn/zsruq3y31tBKKDy/6iycF
KOMStffj85ICOP6Zz8RtUhh+jVWXiXuib2zX24MMaD4+8Hdo0tKigoGMTwqVD/pRpsWyiZHxv9UP
zfJslGzmjRsVCzQMJFREREIAwbz3VQXH4h4vm6jkwQhbJPqnQkXaGuuYEU0bNF+R3zfC9OwtCdLq
prXItEfr8PkU8mIFlxqEGvWB64Bub5oeo0dk5yUP3neF8qP+FxA/wavDUVuMhgvkrPeaLwZHdP7i
CcnTvjUBXABo/3dR4oVzaAw5YZeFDMDAObUr4eu/Gtyk83qPihjd1Fosz+EewMIKq1vCbREfd0HC
dB75ZoctGXQtbpm1ld3sxnprlL8/LuokB7+mXXKi1nAO1RbG+v3x2YLyaFB0ze2fd8BQs4XvV5a7
rE/Chab8Sx0xWtbWgeSEN/5U32RiPxX/vg93R9gKd5rbef4KIIld42UH/LGWtJe5F7SZKUZXCtJA
mNYv6wN3zFE56XYlEzpCPjbLt8mnjqWrUX692WyGtlwJYtWIxYt1H7Cxyk/gm984C8WTnM3SiSoE
yVZlVunL1hA8zKohSB8sdnER0JLik73n55bkEQZ8VrG3cpv9PWG4ZxMEI72PduPh7WjeBj66CsXv
Lvw5lSF/wEVozClcvc4GxtBgMmhte68A8UedMT4G11PoyIg0/WuKj+7vgUSIycF9bnXmp7G2Vyhm
AwTUPMBokhZhM/08sCHV9xge6ZN+zCMPmYy5jiZsGgmjfOQPd2iAVgGXAzmWB/JnDJs5bzO2aCM3
m54Ren85eWXbUvcq6BI4YU6jTNlpsx57VsJuJqp6/wOb4C4gmfct79vBijlyqvDfWX45PNwaR67G
jHst6VKZJS05app63klzE+DaNoA18O5sJp34zNSjm90O6Dbfd1PS8MWfWIQDsGiMLM5xkmwxS9UL
V30Hg11FcMUvr+xeBohh6STWxt3HRm57/Bez5VnweV+rpcAbtsiYEBFCwH2uR23dWOUqS+gOCHUx
lVFVg/wy/T8lb3YMjLc/xIZ0+4YMQx3jdLkrAoL/ouw355/vtF21dtiX5NKauNh05zPRT9kEvcix
OER1xG5WYu1ZXPYZ1hKnBQm9EjM2rw9QDXV6HaS+SrnJTAbt+vh0HyicKclHVwFhwwFYIc9+SF+w
WH++my/Rqi0PV+tZxJsaj+UJJpNFHRleaCp+0+ejNfIRojmOp0unEs/u1c/cBG3TOEdUee7SmvO8
7c6WzL6Ch7R1rp4OUPCgAUDm5PI8x7fx4PKNI58NF4gUeFvMzaQD/GkMoNyHC2svOCmoqG95T5tr
GZ51QShOlsK61cv8R0zW1c3Y3GkxRTIYENU+Ka4WecuoMKdghpkKZqI6AoWvf8CPTjWPgNocxR0F
OzAUmSUF7WCkmGWco5rLkhlMLFfL4y94pOY0roh4ApPl4mPzb3pxncViGcovgDb9kq4M4yQfEzke
8mvy3/LeYt1/j8/WwreplzV2M2SQ84HG7vjvf2w23C9+HNKSQbhIfrQQt+zp0qd0uJ0m/wQFtpnr
TZrNo8l6aEJuU2HjI3G2OqiHw6vjjyIoxvGLh4swfR0jDKEf+/bbAzt4cDQR6e8SIDftkhEgdhz3
e7b8iqi+Xb3TaX0rlvACaPpuo9T4duPOJY6pg8G9lfeRWP92wGOK0Hxt6PpYWtSWWk94bGfnNuya
LPceyJklf2qnClSd8PedkNYC7N9nhDwDqVoJ7EQYQOGn/HKVWWWzibrvRJhjhbU+NaqzaSpKKPD5
nisU5Wq7B0+JJ//xR6QrmIGWn0jwePbUPr2jvzIYXGkWCSMEbh1hoHCVSOwvRKevdgIs9E6krqWq
SOQccA5rnGXQ94aNl8PVKiKGLPpY6VCxGNUR7FB6EgV/fU8EtY98YcZKEsOJgKiqpTtKeT//A4jh
G9cc4lVNmCWFxBwUDgdT8H1w/zbBNY7T7H0SpmQtL6Ijii8DL3WfB1dJK8xa5yGG4pL0xQbmWjlj
ibTs/nndv26v4RUKaQAr7aU1mOcMqe53Si8My6nqLRUkGmCWFMCle9PX7XPxL5trKvfSCfzfS0sG
reNBOxqpspSXTuzeGhAeig1GNdoWZIQCyR62VIsmv6zMxjBU2QvXjxaevgUhay3GY69EXlJxktUS
6JYqR5+BXKcHyjFoxkPncMq6kaOf2/XoDgFCBkRWZyeBJPO458l/DtNkcXS5bGhyTtwxJkpQXDC3
3uSB/e3qUJUEvV1xT1L8Bw9yzc7vHJjqkwkMzTHQtWo+D0bEnhckptMVLE42Urj4dn8IUBA1ZA6P
WEOamHGBJZgVRm+qJ0/kdsDT+tsMj3WP4yGwT72PJuw+vQXhdd20xrVr9bWl8hippbgc0xrkhmfa
f3VPDiDVhOVla/GcGJ3Cm/qX+bYHAn9OMoevRwP18bT5IqC6dK2dqHbpVLUsX2Wf/tO9pDVRID8r
sU9zfLCJPw2PeaI3dr+4GPej4d1crfcLMzP6w6+uZ2MEbTSpRTfXgOHddjQg+lEAfpaLvozNgz+U
U293l7iFS1wgUdCSLU0b1LNOg9/dFX8OEbO7nOIBPGIcrSkNuQR0O/UCPR+SZHZS+1f5UI8lLqh8
s32CUdc9WfVm9SUKoTU/YkdVckTLP7+g0FnlfCV8ip+5Qb6XOIcUuc8aCkucF2LyhnP4YVZ8Qvjq
7uhRgXMzzceXt49smQfA1fbwwgj93NvTj9uWrH61nVIvBQSgX6QArW8NRBRiSrw1ehNbxUrrx6O/
2vQJr0N5yX8iSOV4bHVAhCc89y3FrJL+AR1DyeTK6oKatyvgoZCbTcBsAb8tzbYBP2vI9mZGFZUp
mdDC93EW1mikeZqbyRL41zQ9FsQbCFMLbvN7AJzhG5G1/a/2ZozOczjh3gWWRhDT0tfEYxsy7DuT
fxSW6AbrKuxfCcK++R4CwG69/5vOyQRlXrSikMHC+OuDBALMYPHbrVKU2Hp+6dpff4xMi8BRM45s
3w8uhwYr5bH4KAcqx+EMEztf+/tTQ18bdmTk05NSW7U0kZqwHQp4eppbjxkHY43QZtBhxNdrh02a
+lk3/IWMUCLX8OfY0FOiqTtdy67iHwqd2YBoi4AxGmCN4yevWb1LvUDCM/IEhS5EUwUJVMd/zc1/
zVcoCjHwt6+AZ4XWRt9ZowFQ3n0y7MXBQdwoaRimp6eBQLVcVCIPuCdZlSoS0yDlGc/F95mOpfuH
/cCh7lEmpxymjP81YR33VFHLJH5c1SkVEtPwLGGatB6o+wfCyQY6WF8QDN47H8xYO/C8vUpTH6QI
dbLwe7K3dhbqZM/mT/4l6BFwy8RpsI0CETl1ZDiNGBdN/ReZqUorCygwXwuWf2AG9z3qcn3pjako
lhFge3MLwlG9Cbj/Q4hh0rnTGp9lbNz/LvRMwQaLIQbi9mP376mI+ymwYnBRkjK5YGEsSa0c4isg
qp2hGbaNX59Hfr157yt8hn0zh3QUsHJOODaS0iYVzeLaGkpcir8d9L+VgJHFX95e0FU24UaBXqe2
iTWNdMLFdmwolQ8Zg2Px6YaQPBTJJBzEi4n1nB6nffP9VdmOVzCQbW57wKbvuzuM8lp7vPzyLLhx
Q7Qalm5svJIfXxVvXvYhulJ1M66tyo63R0PZWX9lGiKFjYX31pL+fVdJXV5S3QGNyCkNg7IOilp/
ZoCm+D2Vhuih8jP5YtZjLPoFORt+srasOuEF/dA+8KLz58GbNyg7QwkHAleLGnhyalDAdWF/kvP8
B2QvGY+QBBf1UqvdeC6uhtWluwCJSRmYaBVkzWjfDSwFExN62wu/Emn/2oSeVDDV60eUR3x7itQ7
ilIuW0EzovjA4F+u6TarqOZrbkCFkb06/zY8t1V1KHqxWZ88m6mdu8fPNOrbhWbHtgFSFhZ4/Bq1
yKKomvbBEjGE8vRc+WpT5NvGafYq6mlPbG4GCxfJK1h72eenxjXEE2SaiqQhRiydY6JtxrvUW91T
fmANeWIQtEZGrM0kMYxvmM+Hrxd7ThJBw3IfGAoqAgndZGEgAUqK9YS8yL0fbU6R1sdyR/t8XAB9
RM61jCdvC75AV+s7LLSivTTCgikFCsgbMqAPoURrEoQm6MIpzc/pd9MDMixzfI3W50tprY/3BX7T
RHSqjTL5Ouc3T5IpVmlBXaQa1gaV0659iwd4lkCjirzSHksXNKpDdx4s6TikfHQiWmIFTeIkO2y3
oKSl0CBzSy71yUvaZ3YI3xa0wQOFfIfqq9LA9jOSFI16Tfvx9CoS5c/4eGdoUU2gt4Z0puUZayQg
mHhgKTVlChe1LKO5c8w0vA1eXGSwNOdhWJFLBGwINfcGGBWwZKkIvb59Xm1pGf2TEgb5mdgkCf5Q
eDMr6j6lchrMIjSj3X5RQbwCnoxnPaCNOMtwmRoXZHoLVGIyK6wo2S/YDv6KclqWAw/22H7m/ubk
9mIylINb4AvB/rmsFX6/wkIll+Lg1E2iYLqgpO0ZIyr5/GuhbnvnGvvKYAIK8itaCWO4jg05KXTz
+W7qv9Amb9DcbdlVuYhqMhLqY0VnZLxBeofZcJ7x9RIL5+oPZgg4zC9/DYymTJ77GqeUxUBURHLD
tlAT1z/oNSofGqB2Lz2I7KvljtIBEx90BlrSSetNC6/8K/dQjjqclZXTXz6Lb1OBexl4NNhnCHpw
qRspLoSYwcnAKlGSeJV6hvu/tN7/LG2K8WIisGun0R42eWqkRIXg3cSzjrzOArUcJtV8Cklkv/DS
eAZvR76yIfLcMg4AQjIGzsSpG2OBVJYpE1Kwck8xme2uIH4D4fTgcRRsoMbOZmiyxb536N709bTu
y7oj9tjLpa02BbjpPlMMBTKQZaYyvDBn1HYPpmnQAhaYbX1mQ1SO/IA9OVEfeJSo6e6pBGpbdCWs
P2oR0z/YF/sPXQxy4W6leaWs2B6sOpfKg1Agbs0iBXvJOMVNGpLCgD9HKTdWmjPi/zYs9ndEyjwO
cOHA3Prgq2Z/Apmf5fAFtnzXxL/8AbNHp21t1L0TckBilH3R49tiMbJbND/3xI/yLWkE/VsM+gSH
wWbkwp+uE9vwFm4RBWa21oQymB8Ot5Tl4M76/x2tKxSvf9ivQa3xmFvm3fJhoVfndp03556Lgkgx
sAOBarBBsPEs8cCiZ3iQrk2X2X+Yy2i+J7hOBicIwc1OJ/er9YY2TFLrs0KuWCI15UrxRGVISzGw
w9NqCOVYrQ8M2+qNz1XW/Wz1j0eeD+t/2z1agvq9dKGRZXWqOd/ELRsBxvmjxLvqn4VsuU6qIlE1
FuFczMWmnBOM3SdEC0rdbPoW9bXSbNe0BmNqXICA8OD1CKGeYzoEz4EiTftMzhnnjlECG+S/Au/g
iTIBGT+28/F4fyLsJBGVK+z6zyJcTIqtCLqtdR1FQdkUYOlLOUY04gbpwjnbc1YqNRX087mxAAYU
vZJBIMwPMLHAE25OXs1pktCkOpuiQDtzwfEGN50Cs+6xJqnSPLT6ZxY/8cCyQrfYmKRHuUpxkh5L
QC635yERbXUO7+VX+6/BnSdkQSMLalVEuFtAR8vrtazUgNpimzdpAfi4Z7WibKl/FAHtRv9HSFrF
h3mjEnGZg5TqfJVrBNVzz/qSiwKDqbvjG9y9zcwW/QfZn8y/NXRXY4wAvDWaVhfb7gYoMROCwN+x
xR2GhsR4ftTAe37u2nszEl6csClohmleu6ioxeGEv2dbZ4ELnISqZuePy2xh6yRsUqL9W8XNBdqB
pXz0WPlBGQ3SMZyq8UtMTM2L9bPmH7pYHaEa5atzulRyyCaYlTkElu5Cl3N/dpjocbvUfgR8F7+E
W3n9LX1aMhkLXRBceOr6eoO6h1epaSlb2sMOdcd/VeishXstFc81dmCx0oWJ52DhTbnGcTDK+MNU
fvtfhsydHPOqa6MOls/bwaseDMhNdprbhXFgYfQY1GCT6151qrmLG+GhaKmm/E2vRMEp7Hq4LYk8
zG5yGdFTLs+42OsWzzANdYdvK8oO4q7zE6j42VxoeajxpAITr2Jv7XOE0lcMST2PkV5B7N/vIpLF
k12gk9IXi7zFeOAn/V4/9AeulsEW6ri+WCOZ9xKCrzENObgf/nTJgPVtoHQ6FWtqILLMQs8Abtor
rzDKIJuRWaKYwPSka6uiLVsMcghK3dJ9qSxGMZVNetLf/BAlLs7Nm7Fa0f8u6R079tEko3RdfwHt
LtobD3UJ43livaeGsPYQPRIlGivHUCjfL6Cw9mIhLaXEadKlhSbPB+gPc2gwFirO7WVsloDWRzM1
lKAlIHt7AVo3/4zCNJeW6L3T6W9ZGTBbSNfBsYhQPRgb3R4Onh5+gs1fa2azK3QxiWeMW6+KdvKv
9aJkfuJ9MwLKa/U4IbKzWgXPlf7Uuva5AKHmvwCDcfRjBcdbZk8Di5t4DMeucxd4hllh+2025asV
8AUmHKDg84edTdKOUam//CYIQO+huTSupdat61MHIkAAPh3a1jbPbm4KdOvqfs5QjrQn+M5w0ojd
bp/pC1c/A6GI9N4KJs87jbcZuwC9dbUlIqf44nauDVw2vpZUaQhJg1cwq1Z0Re/twRDqfyMUrqln
M8k2AZ4VnPmCcG7E0YkUhU0BUwZc2flNDWGD0yVsreSPOZlmMtsbrnlgG8URNgBYJgTP1yDn4/Dq
wuw6ZQO8ulTVfPjprD+nymUPnAOOLJAo9rQ9uYvO4VUZvGkiR0AJy1NvfXMi5xhxzcfcVcn64ndc
QqVGFPqULXVV1S1Dx8TYrY3vF9WOopagoJ4CQRYiTUsY9a41bIDj1FKx5LuzUAPM3az0NuYcG/6K
2hgCHCCl/nT5StkSxVUI+iYuu/05eI3e0yBrN8v7zuSqTNmt+4Mx1XKOcAIOK0+1gkCFX/jA41Q5
oTuo/yOVnVDtV02o0fs78LmwT979/IzombBPfclr759WXiJFELkASkpiWDnm5JUHSp05s3bRbejk
bsm2IcN+dFtvqHmXH8v3DfLyq02RtuEECfcK8fHjEJMa8Mn/iwRgVGTy6xXt8EYLmzs9JH/pqOum
LNTjXvpftLHYBbfxi7OV1l2Y7OEG3PLDKzpXy/voiRQ8YbFuOE0JVnhrB7Ll0Irs8K1gnoJeH2jx
a0ToSgZfE3To9/j4NHNmlLugMcwElkyGpNeDM+JLgqazj7nCvClnGkEt7Ib4W9jwqsu/EL98hPJw
F3ah97o01BAiEw59A6TeWPvcRI8liptZB9VTOIKuhwi6p8TxdfClmv208p40Yr8PGPjQfX2dVmou
MoX5vjF4+1nUgdNk/VObLusJa1d+0HCEYIUt6rTHiHZc0zSoITJ4gj/gBh4iQDxgk8c7Sc2HOVBY
Es5LlCdrJeOSWTPFKHV2j0R6QcoLcKjOVBaom2UWWhLar4/l+akKDreacoLuftL3oBwhhNUJU4oM
Oft1fmIHK1gTJ/caMYw+eUkYf6B/j8bc3DTEF5HpgaC4UburnYLBzeesnMdkBHmNtqTtckKntQ1V
9eCyW/2UbJ/8Pse7h8qCE/eBUbq6raMzwYXYktR0rib70ZIHwa6hdBq+gzuAA713mlakFBfn1f6I
RwVDWI13Op9x3tN5kpK5uwsjx3ATZqfCQK2DIZY6r9RfH4Z5fybNtVdAJDTCbJvNNISYnVoTpdvJ
StdmPi79ga9IFBg5lz8IG3w93Bm3dCgVFKtCPHlzJqhqdvURz5HihtQs3lOGvXJs8RwJdYiNtjoM
AsnXL+d3p07pBva9FvY8lesJV0jXFNNabIRbR5S5CzW6GaUh2C69xf05I9IfECcmkSgurh4hZAqZ
xh5LI16WVJN5glTalpQnjNxp1rn0N49LdxRj5FzmgVaScc96+nNNO5fjlNDg7xoFBlPJ+jNV5OuA
bV4hf5ajUkCOUL1zV+knmGxFB/TCZB1XoGQeGoFqUniCkQk7Osr/4idk8Nd6vm1MT0Yory6K1s1X
azl7j6oM+GAdKq6oaLYIWZxV9BrEmuBrz4+e6lg3KRoQUv4sBccpbSZSO2RfuLKVA2Ap5F2Vi28C
L1GNuDPbIOjOf1zVwae0ONCNBaZpkwmOQxCInH8/EtoZsCTXPNxuDrtivUJST1kBkrJerjzar+JF
m2HFYFRWM+eNtNehwnrW1cZqXZwTrleu3dw7BZizPSmDSFIYfC70M7UFloMYuzQ75/k0cjTDjeVp
npp6WpYwvCsFLDbUVTmHysdRL91p4LXUHKikq+/xk+Zm2YDj299nzoEuQFQMy65Zwjc9aileyZlF
y4gvsN/y81U9jzN4fP7hvGRFTLbR7vXH3Hv6Tt/SfKQ2zSAXm6H8GnQsEUF7JSXEniSQ9gqupbbb
gUllWzA/pcRWr62RiFvjM0AzS8Fnsg94xbNDYGpAIkMCV40gRqtPWBGGeFUBXIoBwLCDqTDgL7Pn
VGIkji3ghLxz6XDFZGMQkKzCScfH8rMi2afKYKr48nAPDJTcN9U4Mu5IBHtMA9yz8ZHgdls36qO8
uPmAT9ZbP8TIVUswYWN0MI4YvuYtXc6rq5f7w1mGId6FDQjRN9jmqv+rHxZNDVU0s12+v1cFoFq2
cW3kjgDo2YXhCVeKyZYCMPpjK/xBn1U5ler3ambnp51NROqBti4q79vGbaUN0IHvUBbEAbULVEOY
sTrDa9F0uktcXkoqnOsnfKx0k7WiYkFoD6k422ZvN9e8iH0B4jr5iaqx867IyA0dj9bsAet1w4+L
X5Zz02BUSjj5YuaQ2fgwvqanCxs4YlIktyqkYCDZhQ8D2czi+sgsFtiFNFrvIcECQrdBG6G9N+uR
4ugTlUkHkGjfHudjbnG2USxqm2JuxKjJjcN3SfasCGVZ7Qexf8t41vAnPMg9zlTkOvpX9uF77+KD
nE+ugP+vLJ333OYkFQMjNc1tL8+ADUK4/PgLP+YVqkNGbdWLOitLI4Nx6tNALo9U4p2lvc8jvrwt
jvtjOSBg8kd71qdkXMxlM46JMuJAUU/6SCJI+t8ewWdqxa+1X0sotgdu8zLJ3YY2tHb9MngUuMfE
OuF5ZWjEVDLJqbW9aNlt5EBT2cll4jw/5esN49I25mZcnqgIwuyG+6t3sFk+fVj2kv8AFybC9pPW
HqvqxgDgO+KcdJAv9Wsi6XLobIEkIkliDg07yqpRSZXOjgvpmYeIyYMyh9HYgDsrKc6J6XtzqOga
4WjNgdbnScbL8n8l6sL9xGXu6SG/LNDQT+qLoUDIWhkzPfVOMn2FoGbfWn/a9f76w5BS0f551Fvf
G3vTydhmVwFcoXMJVvjR9KqyRLKq5mQvQlfbZXgEyBTauRICuzEZGnBYNLL4USpNgDKbAR+EAwkJ
ftfSGko+MtY/DqrQNZk/B0VU11nEoYrxm9bLQd2ueOLn8CxuWStGid8vLwA2ghLLWcE76Ka5rDzU
pJ48UNtaf66Zz2jGmShipStVQ2TXY9ZtKgolvAn8h+OTDw10uraBgoY0a6fYn+NZNXer8YFHpQC4
+dG4Po832UBbSPnT79gwtR9CCem6hfgCCAm38aVsYVZXUzyZ3qNXyYqCGRZf/Vi2qx7L0lr0kApX
Nm155NtDQ3I5vuq+3luWPUiC8I+U22EKz3EfQk9DFEXuEvMl54i/2VvYYAwzFmiErH8EO5MNbjN8
z8N3oYgGmX5gbpmVdhIwY/BW/evAUdxAakV644mTpDxY3SNLob3+HA/UTMdjN3oba+Uz9QrYz25U
pNF94OUHJ6CLdEAw69zyYkejbZ1WyfQE5MnSEK52l1wRzHItvrwBsjv7NhEJHaO3bJiwyiN+sebq
98+fD574LD2FT+JB1OVoqfITqlqAwtaELH82SqP3JpXD44z+ELsXLptbIao8FXQtW+tOZcdjHb3L
Il85u8Zqcrz7xe970tvM7OZD74HW4NQcI1G8LigfSst9vf4733pAe6lBJ676RTtSj9fHimf5SJcC
jaZeq28QaeyysX1cDEArGfRxuXZoRjxDQfC2S0ugjRggUXIbK3TwQ3NcdHwE49qB6wqCIqVEu5jR
0gI10MzdTeI1SCCr5SIttbD8EV4lGCoONjMm4bk44tPfNESiDCAnPWwllGWzQVSiuA21N/Dz82d1
BWbbBGFWDt3QzWeLWp10sIxMq/1iVjDYJY3VvS5alIPRvbG3u8tR8GKUvm7hUKz8JSJxZTPn+Cit
kQlh7jTuLDroBNGYFw+RTlqAqkBUY/5FEKCm6CNUp+gj0NnLw8Fh8yKNYsSrev48wW1apRtSgMiF
vp7VM6OEgBBi0k5zxgEuBnFJ8DwN1lbhO1qzI+atusY86X4aoM+ErhWMT1T9PDse/6SF6+Gm7ZR4
2I6/XgnlH7KTAkPDvAqkWD2WqwwgU8XswzyCria5adwctNVU7x8e2HGjEw4X9iHTCXVZUOeM1vu/
4UXL2Ziui3WDwuEGPDqWhM4jJ621//3dPaze8g1ub6f7HPyodofOXfW/YpQjHWpoiG+6p2GJwcqQ
g7Ly+8NdJYk8Cxt0XSx4QmIPSqoxfeRpvF1juWDbDy7CwZvLcz8eXCsLgEwMICiEpjhiYGp8PLbF
ZAjpKnS0uE8q+4omI5xv4qDLjxLupiNShQYfCoSNv7fQFXESQ7rVmfPFVLwOC2E0Z19lQtB6sC6a
UUYAjb5sqTTnsVy4UXwaU1Co7msuN+9g6iPUFWnkF7WJHc6Hqu8yXcjhRUNl+Payzxyru55jGr9u
NFhqgyyoIskKMOoPgM+VVAV+sr54u9HAXhRD0AoFiT5OBeQwivadnV+mmf2dHQkSpjMJY8oLMJjC
fOFdrRqHRiC3jiz/f2DbF1ZflVR2h8x14nqtUir6uZRo9PJaQiLgMs39s0xcAh9nkckjSo9Tm1xF
mWY9oVY0w7dsO8MXpUoauk6bs1l5VqVjnyH7mWbyJAx+ntva4320kvUd2HUscAicE7PRhXMXUQR3
4QOiFV77U1H5AqatZ21gJKjMsmv7uy2WRIJCET0JzP35k/IZTlExj/qYJp6Gjfvo9E6G6NThqWfo
q+Rzezoc9XA76c1efc819AtCsRqfy5CPUwrJRsGqzwJjqbzyk1Ai1BTA0ucXiyIU4reJNTzyx31v
IY5e9GNlQ1g8OoTrf6ImujvBU+j3eTGDuzyAlJzDU69elLZZWVhGaR+HcPXlmu14frXjHGmFIsk5
WbfktNkmR7/lpw58z2YCobwsFQdJuhnFRziflvRfxX0wXDTdJNKSFbIh0w+Uf1lk+i+phVFeSLAr
2k7BC8aC3Yox44X4W+nzTgulrvtU3R0G+9vxJF/z1xUwlDWHxNSmqcQKBt1bY0dQshBJ2g7w7Ns4
R4i7m+l7xiHAWy0MtPPJtn/F1/p4ftdbRragAezpbPn7fRtsLS53OTzuJAKZs4rc+52xuVAYKM0K
Hxh2pqYB4SlXFOtYBzBxR/kzlsqWVUGkLK8TuxLmB3/lP3u+h6qN6UE8cw9YrAnVu6suWxoQHI63
vxXCwSK81/TIls75Oz+4wk8OPxsKHXO38J3N1RD8Pz7+62ydq4jARtu69PiQue3QH1Ees2AgZ7RH
0luzwQjHk0HzVOBS1DK6o++1mVmKCVAC3/7DEJq8h3hOPshJstAPKA6+UB+VYjf+50CO3decw9hA
sVb2hwbOXWfVxlSPf8/+Ar3zaXsAStYiYJ2FQ4DOFkL3w3IQ4/76AUBYoJYNvGR1qYj2Wu7AmqYM
THG9WJVc4BpgtFSsDUGwRrQcjwi4Qs1Aj5nl93o9T4V4TYn1YFvg8XJeiTfm7e8o2cyj24Kchr9Q
GLgE74ku5SRHeTgwPeMCspK0/zk5de/52gHZUWQXNg7sPW3aLG4X9+tgcigE4Ap3UkdrSorl0XJB
r8zroqZjFbn/QkT9ivMQqLgrdAUVew8qKfzcENdAcgmVEhunI33XCe3VdxrqmUOdrnb4HsJh/j5u
s3D6xyCs6FiNDyxBsQbptV10crSJ9ZR9Yl+vB7/eptgfhzJhGB0rzCx0Vngrtv++f+IwiuX1BI8/
35AAXQsjoWZbwAquIxC8jNRGYG/AbvmAlFC07zGkjU2gFqqyLzn3aRSO00QTqDZ+/uIQ8cQljB0M
/a9njbw2oqmR8sB4hbvhuXi155pLcGE3smuzRXN+pU9mVtWD9hGOgTcZQoUeuYaGowerbDPrUQ1L
ITKX7Ft9aBgmr1l10j0ddbPzPcjhSaNwiowZVCkB4vPTrTPflBDfycQ6xSDpxMpdJLSO9tT8aMoA
GYi1GrAIhCZi8jQJb03DJMmL+Ac2NVeyPLeisKo0OerezXiIwniG0P4qPPVHoMpWpDwzix8gCzjm
PUf7u/G6DrFSId7F2nuiCYxAvfEp9jmCsHZHySyR7jCwoEj9+xBpFAFkq3udIOz56P1g5/sHN4us
+mxmZESiMyxCITgqOIKw5Pgo+bXREQ4TIesZFip5gYYrX2Rk/CwZIAUgcmzVk5IkTefggUi2gHxe
+DCz7c8MFbXA/gcaAAlfoBMjn7VwO7pclPsSI0+Go/QqhfLTXLJuxOt8E88GnQJAueDReQoCz3HP
3iCYIEX15kL4jHbL1LVnSNN7pboD+k5qNNssUDCESyF+uvtAQTwMBfxjfUlvXWaSjp1NiVYRxC8f
DCS+ensiv/5UILD563Q9Hs1ls2pHxUf/UN1fLUgqzbw5GBO5b+VYK241sX8HRTKr14EFRoCNGcXh
c7V7ebj6WSOHWenH37A2hpvELE9zgU3sAHuRiF0rR8W63qPBEcWVc+aoZUh6k9nF4zXU63HTvg5c
119ZptPpDfFg7+1uhehdhq/l6XmJRNLWBnpP4j5wsMYSGIqwSdsRI4NSPW7CMw+I9oZJ2Qnq2yNF
iG2qhQplf0/MTIfBiCJt0GEm4lD3CLSqDYGIbJyV5cHsWWxLVn0pxXZbJTldL0zvbM57mQkMsHAP
lJXCjAYhKxfF+9cEDtWwPtnDMsl3LAhIyeN1BR/niqgGhOibYjKapDcQt3yT63KY7KRjtl5cQlOW
EkjlEpdY1olHhFEBEZrBOHmAdSdmOK7F+rIMBFDLmpo/o4lwGBJ4ugVcsLjTr6ifCvJ9acmgZBc1
GSuClSjsWTjCytVj5OwjTH/zDYg1CPbkGmyJX0oU+ilSATQjoWzZStKqAKS+DkdBy/NMgW97fycu
tbpmeikxgafq2eQGWNdeZGBs/ySp19vqImi4HA6V4O4DevB26JSMTBbI5ZOmc9kbpFrhcQMYsdns
wOerx1bGAnhJ9OMnTbgnoW/Rh0rXZpBO8I5dp2YLG1jNx8XE2IhTW88FMQyfakwFeYeuT8gtveKg
2bgo1Oj5d/4fwcbRi4Ohkhiz4g8wLOglQ9uNvrPRc+3qY2FikgBUYRulmBmJ8EBm31iT1ce1jVHz
pux9mXCoe9C0qRiqg1jkdBjx+Whg2K334kJt8vbtvH2hnjjzZmswqHjcWnuZ5euxHS6c6jLkR+Hq
PEylzG4BchQ0+DCiCC6mkliXKjmKxfFQkzRNAgRj4ElNVFQL0p7fZvGH1Z30AxcvrTunDJImOq88
FhOIwF4F1GeN61NF1RpD2NA+eB0E0a4kbXsXs/WAA/6RuFit6IdVDeyxZQIlnQukXpTUzwPl6/hH
nsIT+h+VBNUyhyt5wP/K+YyTpLbf+6EdI2S7abq6lZ4+tuNxHilvMujZ44bdfU6bLBK11rSrjP0j
SB7STXWxoLDeWyxAoCDJC5rxT2xt1StZzln1H0HmWj4rzk38qiNDbNGLtb6F5Dkpmm3t4e1Tosw5
vm52VCkeYLZoNAr4X8mZ8iZODLsF1ZCHFmiIdvzCoDJHNoaq7THvwyxbSezmMw5zWBWpXWYa+JSd
MKMGuiSt20HtU7tYpy/hERkc8J5Qma2r31cq07dCNC/lnr9duX0DLx8aouFIASzwY8mR3cNHlYwb
zSuddl81Tf9fDXS/26VF4LZuOh9u0KFoQPBwIcCRwTK0rCHbBEDJkCQi4m39xpBjW2JKfmJcx9fN
RjmJrGuwuzJ8hOFBedLs9ezctEIhrwW+3rBts/nR2jFG5JQM2EgjQSJh55in4OysCDmYtNtE9mHC
qVmzddl22b0Nj5YKZEDA5byOpJ8sO2V8JlTeTuqNG7P7LgI68Wg6I7j8kRie0kWjLDJ8sZPragkc
eNuC2/vUzi9LYvb65yXiKyGl7+YD3yYUe0vBOMxYFNjCKFSCyO3gwiVozEeYDp4d1Mj/pxc09F4b
VCQkvA3X/QlVVkg+xVSTMORp0aiWJvMO8OxUoIE7e2wWv8W3toJZkxxTnaPGnMBsUV/iaBQ9tfZl
rYtr2cKTUxV4V38cd/V1GijFey7raP0MoKV+4DqkM5DkT4jHop5dSNeytGWkFgI9g63AqKcU37ct
MMs9bBJ+O/UrNoy3zb6xbNMRfUIi3mnHiQ6/s/7NHrP/Qz8NQcgGbd7AdhPwU4nAjnovDNPWPP1n
RwTxTZR2CYvSYEGNtGRlwHROo06QQgDw9WgljbYVX6j9ox0YuSlzt4kvgHAQ2jUNUdLCVoFbiwtS
d6DVRmI7kBlzOhC3JZdOOmRgFsd0ROQrxR05mtdVUni0XQQ0u2waAVnTB0ao3mqLwirMJ6wfMwnS
lM2dAIzqygRl14fE/0Y7bYN9LMtw30Q3YqHnWMnWnOs9oBpK/XVygXBDkvzLtIMu72/BA5aacyUV
2k0e9AmNedokCbtu53nran9WGXnJmXDamK0sht9im3fQ+6hH7KvxdTcMGvdQqqsx98cPItki+vY8
4WDiV13+05jlZJi01zdC8n+A0m2hjsUOvuUAGc008Hot8kCwRGVaOJgvLNKLVlN1yFnGeXToZX3Z
vBnYlt8Xr9ErcjPLUdbRePtYb04APlnquwp7pI9aH9/jSQ0fBMsfuah/wAj07RbYcNmKTnJrX/WB
GGN4cTsz4fMvFcm6R78f3PR1LvJyiCSQwc89ChB5/BrXZgJ/x4ta2r26mnaEUHSAcJOqJvbkb0XX
vjNFKsWO7BsKwdpu3O3/FDFxU6mEBbhPwu4RTd7MSbcIK4TBc9dxwSfUQ1xsLxHb/ZBJkvNITv3D
VOOYzIdiv9nxv8yhrqZu0qHSsy1AG0QyE3NjERzXIhoray54G8xiAQv6Tg90u2qYk2FfcF1AW/bm
KuTVxxqN8XE70c1GabFBUOWdzxDpXyEWqVeQY/i5bAwQ2F246nbID17FJteDkbeZp9TO4eZDFzc9
gt0IlyMnLw97U1fETOgvTpLT9g9ivI9+dfaZQ0lgkHtRZioLRQVcr2Hp8RMbUJPr3ZL+25MTvGjz
a1cua28+s0SvToGrVSKIAqqyI+vqEQuLRUSb0DRuOgw8uohRmXtaJFDqqoLpfVM4fBX10i4KITZA
e5VjJZnzKpkmgBEwyFU/3JkbFycsEpsWGU731RzuJ0iwy4afO/7s9qw5LQoxFxFg4V+fszEabTm5
F99EtVUw0FvuocjdjewjWamE07aj7xWHatEesaHu773exHFXW2u2jHntdLndZ4MYAWySsOC9gznG
wjpEWLJFIRxxsfie4c/kzOvSaMjA/JhyS/EEsvpFGnk1/Bd5KNGmozdzTXVKxR747iVfk/7QPCYP
PTnvqw1+WDsygw7i72k/8vislYTmCjarqLVPaWGwKQe+sZiqv8GLiLcs8BrcPtFH7Zfo7T6hgBVK
zWVDRQSqLRmYV24V/Y0j0Ksnj0UjUujywy6qjRYZ2msI6DUOy9TdlkxQ+SM79mjjNcyN5pJkylMR
U1AkSGG0pTfQOzdNZlPdvVRp6xkZkHtyVWx86a6f5oRdv9PBGlAUeuttohdmTBaXPYx5nYIZfmsT
d98FfHq5Rvaxv2//rnB/bgEK9ayCnqXKW1msmkx52oawQAuZIV0dfrzMnGRpisnbj+bpu0jcpU0f
qMLdLf4kHbJmuySl1TloV4NZtmPdhAnUy8ZteLde5LaEkIzJ04X9IwROpGMyoNhX7syBGPr7CY3O
Wfk50EMMvrt7A/PHozyyhNj+WddRNZv7mURqzOeIIS4x4CrL8loci5ufTxEJyWyjhj0l2AsGQw5+
4CbaggcAn8FFu7MF+QtI78X5298f78t3oo6qMRK4rVGhVe21bmjtqwtbZJtzCiDLPsOeGPQbLBX9
T2COswrD/U7MLto3mkBVcZNhjPEs6DUdLd1tWOUCtoOZ8qlpT4zkeOdxEz5n5Z2Rg/wOojNPakpE
/fUmDPueONRPjQDZJe7dmQhLzJQ0JEBbkg0nhR8oeCzRchyArWgacYl3jR1uVahiRXiDOMsSJQpp
cCApAuSJ3gypUJQ0OA94L4YqigWzEEz1bes6wr7xhus1uz8LcPkXnz6jlkOnm2mnwgXHEJrfqp5f
DdmnaEK2p6IEAfkx4a13wwgXZcBPPaGCiIbS9TYema2ciJJPrflWZbVd1fcerezai3yilKEWTUid
GJY4H0yXojZgd6ZXz+nKgetxUsKreSQg6bY4zfFxYO+yMaO0r4u4/AZzv8Ye+Yzj7FjCpjYqk10K
5D8JCBvbpnh+ZA92L+SXa0I7F5vHRfLBVcwpbwx129kLz1HHhZJo48ijiVBHVQ+ArJPMQgO0FTPg
1LFA1dqq6kgIS0PB6ogWDhOqKNobAVUS9RBFsyR10a+VtLjjput5sk8wcvOYOW9TJth0c3FF02av
gl1k9k/bdMsVR5i0YnNDVWlK8ur4u2sB6gRjfeYi5eE7NkozueECkuKaX2lrwtW7TugYyLvbPRON
rMs3N9OoAy6vqOnG/NDfu6sotdSNKS/AErZbtTHCxd48sfJj2xeqeDbUD9ZBRdeiXk04MXWr0a1n
4+4WGKBHwFl3PXc6EbpX7vURBqdia5Vu+LznsnjOCA2508KvCk/jcdZiowJttyWkDh/HA7jKZkfz
qw/19WywZXGEzjrJsp23hGyIET704KuSeRwdgYwZWg+HbjWGI8RjTYtIfKSqfnaZJONrL1voxtQv
29OpXnnEcCXWQY98FvrQAh0c/bfJAlwoZIzz/BOKFFTeUzOAwM5dKS5tJucHBaEg1978rgyj1Kd9
mOfyCCUUaVCJhiCLG6voc9NwpxUieueJxOqvDoUBeF2Paiuhl+jwc4JgxsDYp+r9l5aVRZYE9uVL
r+gDZ8gO0jxgrChH1HzP5RMaotCG8gnVBAorAln+VS6Y0fR1g1KjJRCUUlInlU7hfmJIA5gKgZEJ
0Lo4CbQOvFTW6/ee+ac0T3vGuaau068jh50VcqKV5ulncOsNT2+WBoxo91SP+GhYyMSJiPHm8inI
eCoOYWnZVRCsUscaM6RbQJ7yaQxH3glEllt4otDzWgGKWH2l2wKARieD0g/pNrQehXT5AJ0EuDGp
WDJR5TMcvD0zuL+I6wa8AiC7OGWI4cTSgQ8ab1FhNyO7T3Oaxuc4wTrgIqXH3c9p0QjOXdIPqBHX
98/cQaUC/pBUYtb0450aqSvzLoR4lCruKytKg8ooVoxwix+JhX/l0TPbAu99GpibsyZHQKqSF3+x
UMvuT6M/olsgBOfWBYl18rioBLjaAGWa+H9/DH2Q5DRsxaeXbMStxFgZ4iZbjH9nxbpYUIO6ZJW3
hPqXPX0PqWR//bkraOKjOchQBxfmGV73dsN8LbH27vvj5iPK7LIBnQTFKapSA7KDi4Wuv8S7lkOT
REfZR8F03UL2aEEUohKdA94lwwBrU2cA7g5kKp5kvX8TBQBrIBuzRshdOJHZlR707yDnCfnMyGGq
kEVVtyEOsx4nvw7nTn4+d0JaUkZaaZv4ILLGMP9ZquNOD9AMmxIctFOwIX+y8PMX4ZiZtSiHJ7jk
CIylyg/h8awrgeReFZyFMr1cbGM0TgcYf4sd0u9IraLAbsfDptZUq/5Z5J+B7Vfea2PVgAaDhOSC
LuRQaPX1CopYJw8P9VHp8V3iNqMSqt+qYINHl5VoU6tmyY3Q0mk5BGWE9MhCxdJwDzSr7QivKWXF
dQMOy+h+flBr8ZuAk1QKNjtSqctwgNLRhfKUMFligHuj0xqPs/HGZa8UptBn4eeICvHibMUPV0LU
4+ZSzZxOk2Do7sOlyShxX3oNlXr97g+M+MKwLOHLmxc2E4GmdaMaRz5TkvvD+1Y0FKp5eJzPAHF6
aXdNU/Jj3Z240csMHLzEw8srCBIl3XkXrhWoOwru9CbdC3daJjmIG1sE345FIcpHefxn2bwWx2Pe
OtGXPy3ohxAoUjf8ZA9qYHAy2uvK3QM2pdyXpvH41oe0luk3t/A4vpUz7lK6yvDXdzBkAjlFedOb
n1F9jFWFOrA3401yxRPxRf9Rgze/iS1kbVXMFlgL2cV3Ed7XVUbgYTSHVvofZZOvfm2CLA9SlYjc
iSll1j4eLDluFhJDw861NxtVkEFTT53g/SM2hyVDRIEMvlJ2bxZQe5s43pg34w84q5xoYienoEqp
EGrN1t4k2HgMYbRIBvsqMt+hKTLySrv8psMI/HeRUblfvlenbAki3D8Bw9E9nx4GklefYNHQQUmx
D8TFRe7Kortdio6zrZQaYsx/fj4Irm5iKoSwdOQSTH2EwLYCWd0mEE0aIxL/yMa/bAj4uz4EI1IU
RuOVpux5QuO2rkO8YyZQ951BGQY5v+fYPL3SgRlRuZqB1p9AXROWidGj4ShTsxxBmC2/hh/syF2+
/RPVxp3n4PJTFMmzklK/91xaMEGRq0crMS5THHqPh9a0FvxBoXvQ22/U6f1bXZCBM7hZtGY1q3aB
yZiTHLCEcwTvOy3midrdx90fub/tufx6tnQXp7COAjY4pLsZgTHQTmyp2LvgzipqhZThoYWd8TIf
5R8WtJ0vwHiy7Li5W+MdrVa3/RV9jtzJJkRGgHjcaI4pdbVaRAXVkGfEmqiMjiA1gpv8kZJtGgoW
nwAQhtMt/MoPpVfZ1DJ8epZT5EGbh1U9VQDehgoC7dhp3vMB/xjqXKZ2KukAAeT6nApAOiSJHSmv
J70kOxHLAXRjrKBjhCcUuG2ha4ppf6LA7Nn8nWi0tA52hc8I1V/4+46IYRAT9/0Egp4FLx2bKDLn
kZmrtpAKFHecMcs1QiswtSxnqAeIkA6omlTZiYaeU8pbZrjh3WqgPz9rkKmplcnu+JW6s+uUUYPa
3tO99fjMgcWtKPQ4UAmwZcYaktsWyOrEbQfn0+hNxPjeRZjPvYnu4tq88PinLFmyjQrGI6FqhZyX
yGi55aR7T7a7j7sFl+RcjfaMzpHPOIrKyv5J1fEScUAsgVGzC+3eYygUnRDoNBMKva3etq4LnM2X
OGz6rImDmZv0YoeA7x108wEpQWdz27IaME9I62Wgay1D9SVb1ibf5fFZIVDu/58E57mdgN+jC2zd
WIS2XqJoM1nNuHKToMggsbojZIO5Tf6hSqb+WXY7a6w8OBapBRc78MlRYierRaBmGfYs0sdnlEet
U0EiAKBsNim0IL7LVkj9xTdyCN4zX5a7Vfh1AFLEkmgG4ZE/aCNLn1pV/2ywmGYyy7zsntx64GsX
sFeEHS7g6mYfEMIvhs2Upc2gHCZ7bR+wPum2bVR31dhBePjreHy+wl3HMqIS/qXj8utYYzfv1KE3
jg48Xex/n1qSi6sJKvKk/2OJmfQUKBjKnu6UAKNewCw3Dn4xU+CN93DycltuO9XOu9ZoEAtUEF9L
fT+v6MsSRoufsm3/A+XNGaQrzZ/jL8cpNeaSx7WFMbhQTqFeTacrUQYVer0eAkuvwZNlPQg3wXuK
/KUWiLKnqCHVQVlyBn4xSUxRHsCtuGCs8s9uPODsH0AUnHNN5rpNk2RjEha9qqNlFUAnVDJtqiBM
SSH1QSr6LhUSlU38bBOReTqgccX9uJ881WmlXKfHDKGz33fxGUcYUdsH1ig1LxuiwF5+HRPt9DR7
jaE33vb9LwZfHAQNmdv+t5GpZ3QJ2TV7TQyG1xnOHiHdamUoG51aPHsxxfvAQQ5yg05LY6hVF2H8
cenXzYuSvQ08ZpROp3nRSaO2maSS2Tqv1fxw9IRpNombxQF4ZIPT9+7L3/lNPy9FF5HxNpVhestb
ZMQl3w8cGzYiBe5JCfjFpXmczq6n0BCRJ8RvdknBvYxiujh9fakj8z1XQinLtAAVUtt0Wms4qbv6
EzlX7usghxrvLHgY2sKW/L0nVgbqXUchc0NpkRtEFXHLW6mfBpOps3NZAEzuqXPZGO5/djysrpeo
kOOnpeDi/mW+mnnjU8Mwo4hYmhbQ3/luggUgzzM/7q8y3MYhdUM7dLqL27G5szwh7hN1ztlFe9Si
FdRVO6Smm7z8JpqO13mnyUPLRiauDbz5IIu2J+AXin3M1dbH9X6fKlEw8SPQ1UaxhPbD7IxytnoM
9ettqlrzsPg5UC6veuBsepO96+O4J0/31MQopmYnf4ACyluWNIXANvfVbpnLtIUJyPO0OiHAmTq+
nSNaDTqcGRhtvPwHq4DKGkQ44/bv9Sx2s4wvWk/jPzXXilavhmRdFZpKYb0EHapmtU9O7Z+aX7p5
umsodEiHzsyrHxT1lOhg0yA2And8lff7CUqm11AxNNsQuN+OxmA09YZMEYLwpTOnoT/mzPqQM72T
9x+RTE4jXuegosTUYVa/RgCvRE0P9NLodJXvWdiNZVzDTXo/XKyF8+b5V61v2Z8BjyYOLXNMFaMr
N+OuVc6pC6RT8rXLQsD6vuBwCJPAEnPwecIZgREKjfbs1iGXlIjXOUyDXR1BdCiSwLLwDWgQqwoW
14uYH2rHxuQ2TszkOHqYNUdFye2D6TOoKqC0i0RYJR2mF83Us/pBB+ihp71eij6GoyUX8da43aMa
3oTd2/XIjhrBNZuE0lxjMC8ysM763My3GumDd3m6NbGzM6JQ+D8pGC2KdBYLWwuQfajyqUzXdb3R
9p58A5Px2JK3FeT/Thy2mrib1VgjqIHbdNTfZCNLhT4JBzqFp6psyd6NOTDu+tSNUlMQtXGd0pG+
FFMp/IISgJy5Q65pQCETs8kfV1aFh6VPkYZmwL7fko9bZ8JUjr9iHuwOGi7sNNW4ORnnp6SgGt4Y
bR8meuIiPFWNlUqrHO6NZJ/wu+7WO3ujikWladWRbdQwHFhxs7decvC35F9Tnl9lSKwi7HmeUjXr
d9rjIJrTeyhgwXQZ6+VxjHEy0y8blzdaDC7iB4SWdEDPJDIvaxR/xnXhBFHA3B6YtZMEyiULZE+z
CukitR6WLlFxaz94wvqV/vUyIbGVGkiXBSdLLAMtRTlYPmQ7RE5kk2sKiSuEveXEw+ybPBFYKxZD
Ck3jdKjsaRdXfnZCVkU2hT88g4ws1IwaxILwOpG8yvx53CKQq16TurPcfHvj0NwoftNeVrJR6XwJ
7S3N4TV605olYGmVouwixDQnSzs4Qsxz/KiiQKJCT74G5qw6Yxg+dvhPVWIGVu/ojRLbEIRt6qlf
AQg2G9ksxkms3Pl6J2q3MzLLQej4xkQJyaPEbHUPU9eI82n3bispRAQYjRtW3cAHLczxzlP6IWRR
vxdfzYY0uUE7oHC1It4ktxReWCjNA1Ue0yv0NwswXu2M0kBGGm5CZL6qBwLC6Ei8KkKVno8KJedf
g+f0msGFnt73Vo7xDNuywywx4e1Szx8nH4pDSP2Wpr7VCeDF1UeFaZkAnyab0jJUkvPwLygO2on5
ewWWzFjRv5cowIeQr0NBGFIGo0MXx0EY+m4YRu47MBbs2G6fQKBbqBVmzmnlP/SN+UvBEh6H60ri
dDT582oqSH/aJ4ejc+hmL0v0iQIXZPdTCx+Gjcx2W4eM1VKkVdiXzOe0LWDEzppWL/dJjwg3wyTW
JLIpOGkvGFM2ZHJ93ZowhRG8zIk1rs7tAn481gCFMCdezxY0cWYi1M0upGcFGZQ/X9qCDlgznEug
ww8e+MeAgSApJFrlix+bOH78H/pcl6JvZS9IF08k4pZtDqUKi7Hg9UaPsr065onoQfNxTEfPDmEP
3aP9JWyr6a0r816NpPPFiXVYMFVLCHBOGEejIqvVX/6XppstlU30jdlP9fzJOtgo1W/4SUc4XebB
i3bqIccmUmgzph5ITywWg/dsBmwMQ0hAqeq6rhdcJ1EQePP+w4vXuNOeOmoMpF/EAMAGN+v9guSr
ZuXaDxS+BZNPjgN9rEY3MjjEEpsrYvGdIAOKWoRI6Cvo+hjIiB0m7eyT/3Cf5efMgzi2uSY4Rr5F
lZOdSvOq+w7ldiyiuQK8SECa9+mzINAG2CHZm4p+2GH7N5MROHi5ZeHyegCw2LYAkgYfoq6RDAuZ
l1w/K3ZVm8LeJTnEiy3AjRDOrxLKozoER0R3UXYbHly1PUVPunzD0Y2WWukLFIFh6ru0V+Bi39tj
gBd6cw/a4/4LOzu0+cfIoKC1bxjx9MwSEZftMTGoHNXdQky8x5H+R1jUlCV4nY1mVeh02mpiysGT
o947X3M0GQejXl8Wfir4KKOSveQCsg8Vsj/DACOnsr+omnJ/O5GiYBQFD1nIfQh9n6snQKRZ1CLC
KUjP1Ip3o6mXHCjYTiIavt1mMj23MQizmk7R7i+Hqfwz9rVeJPG3MtBXTp4ha+6Q+7oPIP8x5KNg
2bg9ZllXecMoCfsZynWM60x0i7DdkWEZJ9ankPZnukcWRz9kDkFuH8l3WyxF41H8q3PjrG0F3/Tl
U3A62x7s8mDlmJJuD3lpXkZm1DddYVWrRj4A+nJtWOVYev9OxTgX83CkMsi4GfYCuBFqkdUsFia9
HHRF4XX62yZ527AhGP9g33/jIOFMZ1iElQ2Ies+/o77oB2X8UtnIhUMicLLHSmM3+dsIO51DIKmH
mBVXPB3i8CyB2olkJj30CDyjAhW/t2V0PQpkvssrzFkJcacFm2WAc5TQHY5J2vBVGGuiJOeNfYoI
XEuOsNAvOrqKoVp/w91kuWF/Ss2uiBt7wYLUiLHj6HICi9h/Fks8HxODjZnNxv8YZC5uA3SAZmsL
LsiMM5yWD3o5WL+0cXENJbDeAuESssWjHBj1zasHqZN3kHP3A6/5azFlJ6kFWS/6PIuPlMEQ/1oT
0/Sa1u7X8A20FR0Is3qi/Et1kdCdHYzwzW+8fyWU8VC2eJB+g4zooHAQCL7tZmdAcu1oLAzr2ZRe
Oab1Xi/lUXtBIixh+nDEInuvokeLPCOhOvqPHrBCvN/TOy40sSC7lQJEvo7+Myr1fuWq7jsUcOGC
E4wQLNwvChafw2XWQFxLXv+YpCw9gJfNKLO3J+A2VaDEQHpkHGpyS3PcvttnkRDMpRQVg3XROrd/
JadNCdgDmQO0DOLyUtO+c8zlyXY8MW8bfGhH1mD4sHbLpiCuNkH8XyVl43OyOVYbuWGu5kVS996K
25ckbxSYlzBHzq39Wrif7KXccYEWKG8q+88I+KbvditboGTBaxOXlYc9iyVHAJqz3R8PCuMDahtr
OJnElDkhuxo4UwfqdhnnSJfd87cq4XU8wT6yFPk1JlImhuff+lAFEpGYIY3Cd++6X36GCopkmb3U
vC1mMuoUoTnKNWflEevpRoQ+Mt/j0Iyvufv8yC0kzoV/ECJqfTMefrHj66I10Wxv8ypjkkMwUV8+
djwNQSRQHBzXsxHKruwmnfOnUN4wotX402g20EUaimUz5BLlbEtN9CL3edX2SmY0XmLXIof/Gg0f
qjFUpiYYZj36/xMkQcIbSNkP3yImyzdJmFeci1Xyw0gdiQrbpxMChuBP0PT+2r3Y3JI0AShvMvzf
hnvY+RNeI2r6ztP9mymHDKnitOsorqf9UJGswNpYLmlSWD5iQgU+xM2DOq0i8cjWR5Kc1ucR6Dk0
ureQHMDcDXxSYZ/CuOEDlZphCcKHFnmb6aLr6443NGxiA4PKB1iSDPKoNjbKc76491jzFxzG3Tu2
wLfysq2c/iVoAl/JNxwQQbVUaCvgKd0pzOQDQ5hXxPrzYkHPTDKTpHKtCx7R3aI9p47GApRtTP5Y
w107rUATNW9ZlB3xF+B5LufH9pl3bpvMhovlGIjY24pGWjvVjq+w2S3iLcIXUU8N/gA5OE/VSyLp
DKX94PaYjmd7l2ckNLVstGFl6vAUD87sINNoWL7NWvAvFME3PHX1TjTHkjt8Bz/JD/85c/a26KUx
fBxJqVg+WzuDm8PBgb5nk17ns/6/v7mp8UAdurtWrvBiG7znyTkySBFhtDhAR5HOge0lCLsCrDdH
LO5Ejlxb8rVB5sunKjjctiUEv4DvBP/ftL9tSjld8FsqHHsIC8NIztkBHL8esqu90JyIWfYRdXnF
B+kaGdthRkq7fImluTlq1T72rTjF1AwwItqLhzNmkvfBC2Hehsb+v8D+L2cR8ieVcO6rit8c/cHw
JFU+V8BwKlmBlUZzjK8ARFjJKf4RIIAlRM9XjH/rXPwmAuG5+HLynk4hlB/vvGO/7stutlxCVubw
qq4/dgUaaHtoGTbbLcqIQXZ3I5OAg0a9hzK9UULqlcVAKdeOSZkQDqjaxydD6t76r3qoWhoNCUXJ
nj9v+pTUiKAK5YmTf45yoG13vH5HQcrJ1LP2q02CK9AQrWApnNL2eK4/NDEzcEtU6U2jdu9xjhmD
hqa+RYkhkL/Vbk+tu5x1ZD+7qBuUlKfirHRrkWkXXMMr/dRMLF77c5TOoYZL9Qr8jIZD8rK31TzO
e8JdbzsesD9cGeSwNP35FxMkS5KrH4bj8dSvP9c6IW+ITmauyZpfUhwDZ4uOZ1XVW5HxMY9a0v0O
5FIGHMZoPg7yLhK5jUtVXjNBcsqhYTVogzx44qiZbkAc4EzBBF5ie2AS7mgZ0B63vJD7FhbzAQeg
EAM7iz72w3Ys1xAtaW7GSH3TdIfl70/pVJLWackKQtd+CHNg2/lwg1m99/t7KKNoCLXnNSTxrgw0
sny3tzX+CYMamGs5eXHjduc5JO5uD6Hk7+1XzMAPCfQrsjxWgen1/XQE2kHr26I+6LyqvKvtYQGu
0Lo42IhvzDKEP8Cz/Fk9pK52Ds8/mFhXQuBjjdrrHyginH0DsBRsGjyvy31aChLjf14crVSc18d+
mMiC60Wp/NzWnXLWgIxWtNeKn7y+VX0IE73b9sXJqtcta534p0zSRyCIAY9MST6DqbzmMbNBbXbj
s+dsR8vzKqsomQvt4/jZrYhqudpSSI1SanGHcFlGIwXoqPiF6cZ23SdTG2I7we30UjieFASoiIGC
4bkUAMlU7lpMgDK+Z5zH9HlhL10kFXjMKsctNkmnGLqlC5k9N6Djn/fY4J8UKzCaClvvtBK6kmvL
JjMzBIRlnF4L5/H6AMi/QBf+RJFKZryx+/j4AFsJBLBIXiQWXKXVY73It+juQ6lO1M+djeGi83+E
VNyik6ksxjL75SJ+Mo3A2XVMWi2xMrerTE4nGTRC0jRDLgJeZeMiq9+R+4V4TTlwWFhIBVyP18JO
OzXDfc4kF9Sjt2ZuCPsgFOEOWoohYfUoEdFG7yhA449qn6B/M4AnRENkztxJDgjgaptm5KRcVSUm
tqu5X2zBI5+aQsdcVpGy9lYr6HHvkm+zBvhEJX6K6MU+AYS4c3AVeGKa/Kd18pEJ208FL0cN8nUA
d0lsHR4rBZ147EZLfWb4dn8p+V3Go51lSTi9gA931ZsqbqMkGrCRhlz6oRjb0WFCZUQVlp9Pdy2n
WnB1OpkAWmoKkilPXdrcsmV9fRBhZ4VlroPwpvYRHyxYolpdrEis7TOmPvMJNXM539OanLwBK8f/
t0zdbq8LaxQAp3PnEOo/eP+Y9v5LXpYUcrXW95rWDSkoonq7GjIRKmZRJ3foEncLzgeyY9ITgyf8
rCFFqZ622z8WEU5lhd8aDgWLMXcaCGnTMNQccsZEw1A5rN3KmNi66UXMiXu/JAwFA6RxXN50ekB/
1AK0pDB0feb8AvQR6ths2e96NwPWTSEhF0ikJwPA3Vg9oBMBof/mYSFHYOq1mwQ3JyE8IrVoTUy3
OmlPAe+AINEBCpNGD2Z/XnY0DtCJNP46276UoVy8cK4s7/zndVItafEJ91b6z011oxbOayBpF6G7
llArUBrC25uN4yLXETxKMC8dW4dOaR5n0HdpkmKUCWRjlEKVDunJQ1hJsvrkU00XEkVKLwGCWu93
IryxeWJLlw3sF0HQlq1luvWtHiloIWLAQPvQkU6TLRKIDte/UeVdcpca6jYUWkJg1CU1nki48Wev
WoHIgmnEXV4DPgH2BJinV1C4GOvK3eEzpWjNp0h/mIT5Kmx2up6paMKYXUk8trlIHrVqtSg/M8Nn
xBu/2sBse6lu2HI0s0X9KJqf2dtWVTSyDPX6ihl1+BM1oOYbkxI7FFOYNaA53xWmU+Nus6XSzREt
I6/ngvRC/Yhe6WSva8hf5rILfQCC5ZaSZvXkfC2p5JKU+uRGW30vh8M37yVgEHXIfxej54AhcrfQ
/yFLiMGBKNT+NYevsotAWIgrM74J9//KQHxd6fkYT1aZaMqOHZsSEaK/Zyr+eeKezYW0fGueaCIX
ZVz+H9h4FzvRoEkbIrhDNRLoMOosFDfrCFNZpDJfKunbm2zaIxgfcX7wZnB6Rx5kfNwr4D0R5Oxx
kgdLBJ0qAXtX2UB9oaoP3cadv0S1hw4cyRpj5RmH4Iu9HA4nPFSokcdiGpIR64g/q83DCwifB+u6
GeasKg/1vWy1llS7VkARL1OVEbhMoqsJvREQTK/Lb7YIM2y+qGx44v1Oob8BblcmAMoWNRewQLKY
oKU4t66EBfgoAhQ8CMkxfOrrKytlVla5BaLDkD0csLBfJWld7c/okaD6v6er/ZmpU7PDVppnne/5
SjUqTG6RllrQU2dKjOqcutONhtPHPuoswuy8xqfMMod5LeNVs/myJft8+ln1ln8Vya+VX0XH4W2F
gip256JY0LINFQzCDPykj9lMVHZ97lGpocvkCvSNYUYY8J2UAYiZYSTj1LqLyVsIAfD8wYiRLjaW
ezT10z6aFvgrG8n95jTf7W3HOHQTgmABpav6iuC2N9l+NIfSjwr6v8gY2AKOcCfF08k6kg5v8vVB
JOU+Ze72PNvwnlbGqHlo0doZc73FEtrqcxUySjceWlMtIm7IO6K8zm7z13JQFE+LsV7dimCFH+03
vEBEUwajfnSjUbJoQ/d7sib3xvwrUmAhe6ZIoA5I59X8Cuc7DqhLPmSvMbsHU401x9rkNrJj7E/y
vDM2fXg52FEdTsVbEm/c1P15XpLratkAA+Wupx+koMqoUt97SXFC10NMzrcDdeR69aHiESsuFxMd
qOIPg3dBFdfo13igCLQDBBf7oBrrC8huiCp83hYHKb4x515S5ZolQoCmwVyK4bG+eruDBc2eDZRH
B4nZ4KBvaTMaV4W1o5L5Tk8ESJGO7BNzsEQd+f96sDP5SNMmbIdHTEvfkah3TUVWPgyGzKvuv0Qw
z2yyJjFVY1e8miA6dUuHzKzCLpBD30Jrgn47l8iXAUosC3Jw4u2WGH1K47S+H6mNAtCKnuoGH/OC
PWcAITugVF7nAP5cxZ0s2ISxZWDmXcGEQdUr0Tlu/iF+RANp9KqTjg2j/TtP7mc6tni4VR7hbCJY
/GCNkGA8WFFGdBL1ZDPndMnSfgYuyn3SsNpy448/u9s3ayWmvDZwzZUJpXEQYrxzeMxN4oyn9B06
YNAWzggNT0/36aI8Hi7x9cp0MVd7GjS6LWFiyFEsvxwKaiuLFSTY49QWCVHvSjb5Xx4TdSdYx4ei
17elHg+/NM9YBa/qK/gWRfgnnP/P3IBR0DgqQBMMM/mNvsU9u0AIdQ7F8hVlLik6vdxYQw8RoNRV
ZpokAIWY5BsadQchBLyEFWdlCy/z2vfnJmyxy2PLiMoqQEHL9NGNYffTli2z3msuwM9IAA4NhGE/
S2Z5a4CWgBOWwZqloirmCHKoyvInV9h25kbqBWjV0aJ9pxb86qDastKaUIQNJapsDK7eBfnQZF0k
cGdsNBIRUICNk1Ozap/QoboRZVVHwJ5Txh4rdtkEalClZpAdO24HlCyKPig3esi5q3Nn8HWxZWnf
bVsM7FNZDNpzer90kfpo1wLiVYSxBQDAqx8g0zveDwopjJ5Lz9UtJ3lyS1IwRoTBsJ9Mhs3QXlQY
FOUqAkdCUS05MjJ32EOLj7K5m2Ht/72hFMSF9f8gWAx+udATVknbQKxfd5QwRB61QMXWFXzWvklT
HI53i7A3UMjOCa8TYhTd7+tiTw8IXiUPfFiqg7oiL3YNQeZUgGW2aGNQAd7IivsawE6heE/GH437
R2n9wky0Y2da0Uxuj29cVH80KvlSj3hZdBxwi3d/mkeU2Tx+IfyJP53ZfNViFlcYbiyN2CxNlTSb
k+2lZQHt42EKRQ+xZtBEA3Hllm0Cu8X3UYjjeulbubZTuXs9zMFnD1NWb5FewYP8q/B3XeUAnZnX
nflwIwrpLlPvUDBeFseloMCknuH8fC6gLEHxBy2mQmpos/83moys2MShYGww1KdBRiSziIhHSbMs
RsfpcqLtLDuhcLVYQde33j0M8FeI9CLQLTcLtkrI+Zh/80cWsS1+HmiObdCKWjSeLKSkt/0ioJCe
bwIRpY+pFD5H/3WyYWRXHUFS7jQc8XqkkY+DZUmjQva66/Z+cEA4U8rkHy1+nQAxbF/rQPtCpb/8
cGTvmvymfRB4pyMxJOolgDmIMGbvS/UMt015CZvHPlPTSC23xOYqM1OkHwd40zayMcTnCr1j6GpH
4VVYNwtA75Q5Ff4pNs3LPnW37HvTqvjOOzGATQN8A38rGtvqRCLVYxD0Yzy2GwJykx8zkep/nlFV
QG0dRx0FLMk1bUefLmRgSY9GDmGC8/cD3zDJSbhPwNaEc6qx8UmckUCiUInJRFBTR/HVBbMQfolT
qhzctpKUmfdnTDSiehdF4KGoXaVFlEpz/yQeOWD/A/pC5e7ydnEvnkxMyEvHTGEPpJbN1jT49jLa
5SyiA3UARqB7tANLqBIQjuCcVA1ZVYJvv3fKVv63G3xsPVrUzKc/J/3fefeBwrHVarYkKFob2lcS
6d4kou0nlHlrorjf/IlbEw2VJQ6R9LzMA4iERj96/Uy/3CufjOdVQBwCsz68V6UzrKlt1a/Wxlm/
U3try6z7HACrk8dPJxcuoaqKyipWxsnObP7re6UCgv8CYm2I7QN5u7vQvbnx+3oJlGkT2cCstUwY
mHMbgPiQ6IJS5ZNO1mVj9YYEdnCuvTzoVgDiOZ5o+DtWHFDnES/XXInF/NntMlB4RoxrK9rTaSrq
WNNIhBK6VPQh2k8H4OdXSdkq23Q4nmQk3TFN+j+CdMrcvLaWQiMySavH/NB5pDvmfJZsEhhrbxCK
0cHt9JjJEthBR0IvpENjPalBa4kpGe/+zuX+8zCnJMAXRARsuk7NMUJDnrBiiFbgOYSD/JfgQXw6
MLJ7iGqKpLlYtO0BMNv0Lxxz+cmwlb1PpTS+h6/S5YEkISGJMYZwZJQT9xHdLeyxXTDrlPvFoQOa
I83YxKXY24KM5haCKiIijykJmQOiacW4o2qcRVEeDVmjaB6eAxszoUApE8KcnY5aVj5+/XuJRXcs
5ckxgkqmioYjG3/9jrTC3dfzFsXknB+he+iNvW8M+QreEzsazZz9R1/8YC01b9dnDc3ZnVN0C7Pe
rYihmKZrkiNSKqk/Etf66sJq+ug6doOzv6vfN0Cv+PhHFzd2VyvApXgZLdYkvgrSF4vxxQFbn0cM
tjG/rS7gC29y6LnpTVGQgFaol+CXgp7SKGv9wxkKtKrYnKb1wyz97xxc1mztc4rcAh+juSLcLtJA
Zz4WDe7NJjKsn4XopdmlXMwCGeNpDOqoL1OYwfgrLNhTAkY1aZ9GZByzOrmsGgA2XJUX30ByXB4F
WPAY6sW4etIQu8tCTHs14v7Ugrh9ZW1opj+u+51+yDvAKSIaQwiG2GOPz35bl+zqIEIBsBIGLDkr
8z7+uz/G0KV0+rANVFa7bQ3dDr4kvPwpUGqAYfWsMcbs7xzYm0c3N+qxpS59GwFryMRa8kZTLi4t
XSl3/QqV0USWg3+jQq4kiUtSF+dPu4OW6yKDSiJhC/EGurJEO2VavhvWylhj6KzNprQRAtn/2UAb
SGU6Kc4ClHxUAMJyuGzApQLmhKjL9Le8dMYf3cCajSHUEIFtxxqigX2OMW8Q/cUSgMi/8FDWcV3o
TsNiPD0nZQ8ihuMSLgGQVdikvwlL6LpC2C+5GsqC3gtH+3Mo0M8dHzE9+4WKTIXJdDJRxSMjTXGi
63YBZnzcQMai4+s+S6m3pER3/Nn78ctKQGPrCuzNCc0Z3hHpJ2krHcyGe/O4XtMjIhSjFfkgjpKi
w/lAY9iEOo+wWU2Jp44oqyf6eUhV/TPjyd0Gn4MKVPrKCJthuqonigfo/dQm4IHJp/snXpw3ITr0
ZFnO/tgbHv0IDDJSu64hCue7YP34GSSObKKnpsevw87auJMcXpHMKV2QEP5dxvw7jrvayBXGR9mS
1LQr9XRNc06FHKgZu1op1wO4poQLXq6GJYNlG4Df5TYQfkvDXeXwbWpTkYcGJqHN+lVI7hdP/vcm
hC3loxgtE9B1M6ZvOiFC3DOpKHOAia/E8iVfWA7unlOmi03xfJiVjmobXGpwI/rgbfr0oGhVdszu
XAZRMb50LRF3bGYfiXQZD7YwcOAmXc8s2A+H6v5gT5I6x0hoW6YvWBwst+CQNK1JD+TfiV9KjTxb
ss+Ez+kaMFSSPSD4jA/XoXdymIaXtPjLTs3bzAPsqyKdlq+idM/TozlGdMgLNIs8m3MfbjRMRi6y
s1e8Dmsp8J/O1hqpg+gHVj73rRbgdkqkM8pwbSZMa5giuNIipCjOYD2s9eg8xw7uRwz2a0hOGipX
O1VY79SvWLiILaK/Pu5Ao4ZQcvDjr1jAKHLp2kfkcISNsyUD7KbHToiQ0dDQ1/ZOhi/T22vSjxoK
c1+PO7950haUGMlV14bLY+cj2SfSZc/J53KZPmpYucMk82tivdqcH9mXgTKvy1ComGyLDZJj53Jx
DtIV3tMRxlSEeeOnr2KvWGS3GEJAALXMyxIDiNjqwr845pzfTGEkolhPbyJKGb1Uld75a60BfduL
VzGsrST/+ghXBHotTYvhATtT11xYUDZb8coyYBOLqf69QTJin1oxqdLN/hsBFQrB69M1ga5jaaRJ
bcldjIM6lQDhz9G9iwASR80GdUweBP0Bz3C8poa4DhAQfeCg72qHi8M4Vy2gLxveLQXU+utN773q
ir+e/mpRaSysifwFOGkl9bg++M5CY8RyNQPs0vEDgWzIuR2MIt3B2thOKO1RI3ziCPescj8pVmM0
1ZWTH7VN3Iz8xanWLuE4MgfS2qjsdVbmWeykFZeRqMOCrWNesLGHFDP2z0tCepLOHPTBHAQS+BY4
onmUF9/2jgKEbUFgeDkoPgQq8oc/ZitrsS8AG9pB9Z9nkKS26Iz4DTkqqBo2gusMFb099S3AyX8q
2A97aSDwdW8eAvxhi7Y/eoX1CUJZiGhEvhzfh3CxjOHAybjXe6sdyDeqaBJGO5BnG5WQqo9GwOP3
YItjCSKA74by7NQyWSqFNAuO/2hm80/BK/7vAHAOYdCm4PAbGGbC86qAfejMPJMTB/dETeY62vTN
QeJpcWb8w3bsk1s1yX3y1m2PYANKK0xUsGIPNDUBWJwTH5DqQ4+bpuxqPzIn13qD0uBwxkTjH5bh
BxspDlzJubXtylb4oMyrdCicumpuePXqfqDoDe2MWU3GUeNObycGColWFWpxWgLJ0lor6iXMajLJ
NPyL4QUT4I/FPQ0E6FZ2wXJHf1rONRKULikPsOvYKeWumOBcqLxLp0GN5PMmxWB6w2ES6lpIzSBW
RT+qBcgjwWwaD0IRk/HAHNa2xGKgd24yHJeWsG/Jd+1GEornzSCgLUOeRnB8VDs119lIamCRUxFK
xQY1+xjTT43UMcEXK2W0rCe76xzKcMtGj/JWXxg1gaqzKL/q45lezfBcL8KPXPInQh3QhRtProp/
L9eeajnjkywJJTa3TTZnUlA02QNfqdZN1c41HgVXnl/YjjbGinLxD9aGzbovMA83zngRJVLSoyQB
BvdyDkb5soO1wtE/dk83Sp6qq2RnlIT5zUzlSILzoJk9k6hrBAzffjhPk05HUsHlN4pnok60gyV4
eDmlvoNU7ABq+JliGzVnUgTEFCOiwfOMtcSITICE1zJjvHA2zD2P7Yw3393rPfAf72c1ojqhIi2X
2IVtFEMc8OLimVzQosPUrEjWYlZVF2N0YXCBtLsnl2ehJLbOxW31cupTdS7+Pl2criGVZThEaADY
BJ9BgyqqFCbTl1b7vc2xncN0vabw4YBuRFhlL8wbKS50abj2XRwR2O+1CWstgUfuEFgEdprzkyxp
n7DoBpOxPhSdrXtdAIUHKsMg3vaYclksYnyqlVidTz6fr9/0E9iY9DdPGLZgnUIaLcXJn4AuaAJk
Pg52bZBVGKT+N/pbXXtnLhevMYyjn3y8/5eXUgD/UeNNyASvyztMb6lJovgWnh4EsJaBiRBLNu6m
YZR/QuYnVxf6RMsdvMT2x/qsTq40gBq2jLoznFiWjglvQldbsw3h9/+ml4WcZrJoKLbDtTN3htYz
NbYfJ8syT1ML+8gHwwDDdZfbgJNZXhWy1lxK3oK4JkmVIzBb9Vtz9yn5bIP7mcMJCxTg1qPCrw94
GBKT3PO3G5CGI6P35Qne6hBSAvbk4aYP+aoZDkFGr9yxvLAZrKiL/CBTWmz0aOr2jBS0njlLGZOj
a2u9LxTU/CrrQX1kAbqLBreP6zUhRljvu40UvvbEt7Am/NmKotmtP8aegIYhIiParVYot0xGQwyz
pjhap+DXfBjjVZs0+EcM3Emb6fAH/RXoMgpmVWpx/Nu6OyXVmA44eJihUJjndkdVCcD9dRdM3khU
ZXFh0sjBghcwnqYAfky1fEu2eKDuaNNMiaseOs+lvD5TCOKg83kVQZ8elfsPvGsrwcJJYTXenzns
BEa6KB5jOM66dfwOTTxuvV7a1HOX9s/t8jDwRc+TShXQHAtXhNZrQcahIyfhRih6gVT7CviviH1G
/yyb7NdXO3JCeQk9l9xQXSwHk/z12ZiHxs7cY2XtjzftFvW137gQHzLIyflG3k0AVl4TM3MYsKa7
v5IoOKaqOoBUFjSMiDUm6tz9k2a0ZbBQSzNZeGjX80g5EOEZfJD5helxykfYXpyT4lQRfGBwP9Zy
Kymcpv2+ApAFwbBkocHhcxm6+NMlbuuv4lGH36QaoSs+1wzUKEQ7tJGiaQFx7icACAIZPtoYKEKT
djUXQzQumXFKrs5nMlmIDYbbv/c6F9NTL/AsQ4aEajYuLd5kLZqA/ToxTJ45sg1XR7WMRC8DYtmF
/G8P/ifeih5+DaAXJHHpUAYlyK7/7KSsga0dCD7xGyxxzgrrds33vh+b/w1CSUTBdBAb+Zv6Bt3Z
f/8fA/Q1Zvm4NMRqU+n2zwO+cf5f3BsimfQFaZVARGNA+nlj8Y4vrFXQqz72CZIYAF8RhDK9NW2C
8o4I5RNuJ0Psg5Iejc4+dqAWMeON+quHV2LlswYqZGze4fRsnxSgZ8bq/dNZ67tSM1SjeF+E49eC
i2eC8QCqEzJS92oC9mUoXFkD2XXkGHRWJ5xwzjGorvUCTI+0ZSED1o06tWITWMBgdxalQUD9ds06
O1niJWwrfFfL+D3OdqXjRlq7dBER2EujxP8/jjx9R++4v1dI7IMG1OkCokxh+biE/Jxi+Yaxo9pr
JlLVzQc3DV/YYfyUlBpS1cXHs+UbkaVJ343gDjGcCwUPwdI5FHv9m1O5ZYHTVpId547y//VzMzlz
giApgykP5D1Z0qzPrq3lT9N9GNMr/4vwN1BsaW3r3KTxGBovJKzSbJFTOPwG7GzQBMztHS8Tvy9h
5/Z9lhbqAGlmnh8xmx9lfQmHlUnaFfWuYZxqNvBU9LuIC4YoiyBS38KKpFoOklH/Eny+Py8b83n2
T3NvX9BxF+DAKntOuPKBKGgnbiOJo97GI2WtrcLxHtdnUieusmsPfo6ZcfT8fUg809BuJ3OeuYF7
dfadfISeCQZ8GYg7b7F4sG9ArQvFUX2zqIggZnk7gFnZbdaP4d5B88eODWjsF8JF/KVElsgOj3MW
oUkrL0Xl9dY7W/PO/cWwhEIKa23SdTX3OEKHr/5TWNC5uToMEbJmjFNWifN2Yl6emQFgGzjHYru1
fhU6estV9h4bwQxImp1KxTdz92rG9LJMh7iOEPmW9fmdmmUQSVNQq2ycV8VovqQpLZjS7yTygLMk
HYKGkPQVoo1JS+vtOVHBmSyJ3XEtyjUQuQP8EE0cRXkOKdmBk6h39+EhS1SuMn8DnoiBA9dOM+DY
jmHjwp6AlpPiKpxpnBDofwRNjD5HWH/JyrcXNQtzfxmslUjtRc9xG4T+YNoWpUrG9Wb2BCtQRGjF
3iiviS4aOOQBq8JE2lKlnJvGFbsi8VzkV5+v084MlA/BkiYVPQh5WhEVgnO4260OojUKtwhfQjcB
gmucWtwVVs5OLOMTvLxOILxkYmKRu9Yk9ha4miVS++nugwMcHT4HNzLvb+XD13sGFT9IbFQm0sat
Zbna0wSOEbmdU3GEZNVuTnwQiiax/2Ue5111A8POzbGFH4ZcImSq+hegcnjwVDt/4KkZw2Y+joLh
Ixwn69lRX9k63TYDZvHZaltiaJntq5Pxf7K4e1fGuwyKegeIFhvUXsSqCBVrIkUkoaSESFeHAgJP
yUUMU1/c57l1sxqLMxj1l7kKGjhJ/oDl0hxVKSu84T8YsOBs9aDjvSB2pjyNa7z+H3KRKez2uZ/f
kz2R6oSB1vK5K+r5Os3tgVuGkCvWmxzkn3CbmBpXQB55qWzE/mGsbrxxhgJsstvLwbcGjwc+nLoL
QCFTIToCrzx7byPBrZKjz9AOm1aghbMXSxDees9TrV//OgThn2CAF5RQlBq7HMoF+GJEnAjNVCo6
HBFZcUTGcfHDp4qU5aX1jr2Mhh77+lzY5XeY1qFEHdw3xdI+w98sOeqjTkC/diTk8qmNoK61giGj
zBf3Kq/z2i+YXCxKxehF/AY58U5nH/gv1mEMBc7a7KARk3NWVD46RIPjNE0pSxR7Uj/1SOGKrdFM
H3awLBfUHll9G0R8KJcl27MYO8scU0voHYyUS+IHwClbbcStpN8az625WHYbJDXPzCNK+cqPzDby
hRFTdL0Jy61xmvYHz85noBJNcS73KSNNH/P4IHzMrKYCzy40xWlp8+bvku/C32LEmoqqnri9DXPb
/y72BB4F2tOf89zj723kVCNKhRU6d1BCPTNrgHgr2wy6qZxsRl7xdy0eEA4hREl/AOLRsBPUZjux
IT3r8ff27sijfdroWS/NheVkS08YG0VBRGZi3+YiJtGcAqApELfFk32LD9OHMKbphP5Q3g16LXFu
Wjbu8OcQmQPtyb8Cjl7BIOgjfTvBmgt/2J+Ox7ZU+jB0rt7hCVn8BxHe8DbgyWCxmvbVMB++vhbL
qPjNVg+3iYa/IEG4e9lmJRrRQEozXz4buWZaCbgUWfWm5reqJJ9TNr+3/rPwziLHiSMqz89B5gKc
fkqcn2IqD1xD1THmVIEG4V/L+Xu+FOUY6ebsoU+0kkPV/iQe/Pe6EAk3RBNiK7GbfK1eEHI/nLRq
lyx7A4WJgpgu7OIN4QQvRb/WNViJytLUaWpNUzL9fAOQaDdzfFtUitG2IkObSpR0V48WyFqILaCc
T0ZuxbCPuEqUmuPWO0b9rWWBWWrHKHQnkHVK3iuLlbFSNFPteBrzgsB5DOGk/hRB7qucxjoPg6O1
LGZhmQU5hSLiMTr4BsqdVA/agbRvBqbRKyEZA+FNlS9nfYC+u0VZfTi5c2HjpzjXiBdWV+qUHaq8
kT/6MCWQ0Fh0ZOoi8hNhOSB7TLsutmPc6I7jX5x6S36GQzV7UJmNrs2tTOQQuQmzUoO+WDED1zDE
zSapogePOlfojy3OpKhNlzjywToSUnybdYlfCcpS1PqfecxP21SCN2TOf8XsowE8Eh/5WIUFsnky
CVHXpagLF1PaauuXH4ZXr4WOJVKtLHWbzNuQi34gB1EG0uODfQApudTsusiNc9wqxkif+B9zMuM9
RPFc9qjUXHa00abS+NapLflRCGxkJFF7wHc8Oa3hJOHF5xXvh3nj/2FyRZt6fny1IZmSwMAMwrKA
6go/6rdBRf+2mYpmCWfBkKgrJ3BcnNT4h4/5KOnMctgynOqiDmkHEJlXXOIF7on+PkRpNQBcfbLB
jKP9gffbcforMCWiITe/LfjnqBqUwyMOMLc7CJv6/PsI+HUT/ewgnaaS6j1Mp3K4pE6tvmr6Nh7T
Vhwn6/mkUOPJzXquv04aOsddKuuY6L4GRh285yTKHUBvBKiCdkF2jDAtW/fqZQE+V5JwwnicGmQy
xY2xfkswp2BOFPXSxp9vB/P1gV0xBQHLH7XpXgff3/zHb0rJ59foM1uRcW+C2b4W4vaXBFV1FypT
GBntQ4xPJBBeyYgg7s7w4ODfaomhqg3SANPgCp19eyEpxGIafsUgjE9Bi3ta3PX72dpDF75V90ki
cXWi74Gkja0IP4b/fCDbMqjaGMZDJZefhcdFpcmaQzZu+w5EBl475aU55DzKwSiXaI70Xrlw228x
RAMR3BkXnEwsxb/uGqRQmwdXj2SJ6ApdPow62N4vtFDMDEOsnnZesC81GwvwJ2NKzp5dEjlIlqVG
VLBpkqAolhKHKg5Wru3af3iqZ8VdhF92GTxnVkKqAmdAa4aAg+ZHtE1U0Acur3AV+4Ou8GxbuwTZ
UciUHeYjbM9oOiDlxPwLfctn3MVsbF5Ca1WD22S6rsmRLgVyrQvD8AHx50PShRpqY1rC4R+dAk4n
v7lLM1RUjROb1LrAoq+VVB7rrpgjLeRjxT9Udhb1S1l+J2jUPkLy26ZTwd80B26vaSREvPLb0kYX
3pNmG5185M4OLHVVz6lDm8wkMslMnCxvp2MkTf4inwH6+2dT8oh0AEe82FyrkENUgWD/Et+1aeRP
62R/ZljdcMS6wkAmp3YxxyTHGsUspUrYoWcLzX8ivZEphx3uDba6UXrikPyAUh+OSZDx9v1bD8D9
eJztiwuc5l601MLy2QMVyBdDo0/qwqLf+vuNuull+Pg7qGLrKlWSJicbJtEWcAhYbqkvThurR9KR
8DzJrxHQ1o5HoHHUCZOR/J3ZyUZQC8RCWWSY7esFxWNrGvq4m4Jv5SHR6FmlE2+c3FVli9ZCdOVm
BDzUvISwIP8rUyoT/2iWQEbgid0x55ksR/FRWmHt25yZ/KAbiv1YNcLcAl6FveSWbnToV3UjV0EA
vASFgHHu+m+av16II+QKk86oZwPzZ0A7d6xyzzIhzNsODEuCCv3WY82SjEL0lD/PGG+s0sQufgJ1
M1BoJUgK/oUJdMlh8k/3r4JqmSCE/2l5xoxWz4uCp7FOTrHIx3111mlzDmMyYM1+bMg/BI76zfy0
agqK1pAbSA1IwCvjzceJnOUZY/fNqqTuwWljNe0taq5TkOkWOd163Y6uhzvduN5w1uc/fSSWBiuS
+cDjsHGd0nrzmKWmigpqnuzELRWEhPLm7VOXArlNgZVoAextnpbQWOG4RJav2rPKcksNDWKJUYz2
JV4ykqfwJf00bwpWxApsQVhmgQsMlWgMaR2JUAPtMFknnef2xpxW1lFHXHv38o2rzuGdPKYpgWmp
+THh/Ixqi46D2FFgXxT+awiJOR2mAcuajtfGb6sq5gAxiO1I5h2BhrSE29hu2ny/myy7Wdg0lqpX
ophbeEulkUi1h1huEjrkCqXlPEYzJxJfz/B7LdSsC7oD9udTd2Pm9M6K1FWg9s/D9mYXwUUjfS78
BbcVS5xyZi12jbsGI1nVhEqPdJlQL94Ja25zjM6j5g6MGhJBOSoNyk+UCa7c80wegcnJ2fwAAphh
xlhGuHQ+OxWRCqGcjob1fogZaX4n6YIkT03i7h0UzFUlVsDgEH46rDYAn98jTbeSEBQyoNrNsnKM
81sZjqLiFvONeJnoLaN43gLkjMVM6x8LDvySXCZIRbR/r1mbMEVcNXv6KWObwToixzrfttHufNAF
nPfA0dvn2spK/Ddw0UGnoGGAWc9bbwDXgOIDxtN6Zp1P1bf3gk+zIXeT75lE/oiRg6z8IS0MYcyF
yaUWvPScCaeJFm7Kd1bRpll78MDzfbJ0sbS8RmIaxrRMhG3pQqVU5gGGGXxGeFFgv7JCoEZWDpdU
UzG2lUFHrefRPfBLphapPYIs3DBp+vBnDiYSizTmOqikUCG+lTJJD8ebG63uibT3ix85pFzog+aQ
SHhqOlQ+mqg4LeAgtt2e+Qyabbh3njQl+YF2BGaVN4m4IWs/sGJgk9rWoZDX2zNXmk8ZqzAGSRw2
l+c+eKaUjSSO2vIo+qpa8xxGAK9EPUONkzrAkDn+ymyb+757PiwetKJ4PJAjIxPc1N7Ee8QwU2sX
Zlo9hhrKEqUHDmAf+5nkkdHUEl2cyX0IQ7T1dd/vpXfNPyLe6DQJ5c1/H/kuz87i4ZH/2vPh4dvK
/yFZNWLkw4fbQXP6u1OGtafL/BGNDmv0XLrDRrsBH7Y9jmPwRaJ0G3MkTvdQJcfTxa4kBFNIK1HI
iPDT7aUmvwapwyEuzlZrTiG/CgtEbTpLYdwBoKQ7RSnOo3rRshEt97qKZ4LtbJlz1N0V5+zgGREY
s8pPZTpRWgac2Fc7+14IwoUvNqZzObzM8va+ny1OEkrnVUVH4nzEaN8M9kr4GsKscstXJWXX9K1h
yNthlSv4Sei+q4TzzMpOfIc7xUOI3jS3XFtVGUlSrnhiNGAsTrVFOc0hXCZ7nhNrqEF+o9dDptsW
CctYi5Vfx2NRJvmS1XHLBSucXyVGNa2q16BNo2OZzq/yRt1Z8E9XIf1BgtnPe34vJHm0ZsrVzh1t
Cqi55ZhatucFJc739mX4iPpjrZ86b61ka9U3Rdw9ymS9CMXaq22Q14KhHfSc4HRPr32LwsPSOWPR
Ob++6yKHKpXACcWSNHWL8d6hCtjVg2JX1bQY2dK1QR8ZlvHZyqAH0ZnISWS6d4qThH/xhVuw1PlZ
QVmaHRDjOH38doloeAL5O1Ds196DbVK2rIdZnvuihG8xJGS9tSCq0ZKCdvU1i3BFwL+n+QAE+1/r
nfBQxoHB4D5sDQ5ORnWk7wV4ybDxPQelgdsW+OFesLUnm75aSGtDhnX6yn/jaOhmBmJ0B1Kww70h
vX6sByzCmlnYp4nXCmZOawuXsTRMppyAAF+k4u023lftQb7wuSlIQzP3ak/LaFxi9Q9mG9mrZ8wi
wq2z5xiBxOK1lKPg79KrdmQjGHXdFDFMiUmoGFt53zq/UbrNAPrmtHA4x09+mqSyFf3toXMVRNin
E4Xwprms7nLi07UMk7NsRlh7G+qoPUWtPicuUkNcyn/MzTAoctNL9pjDEOpsyleSE+UoYvlKi9uE
4lSSjFWhCxSAAXf3rg9oIfIKJzBMrQZ4ILt/bBOKsD5ynHUoxYeIMchEGfYrSHe33mNwhM7BGopp
QQcTsOOZXZLmVbx+z3sMohZhDVdxBXhje0Ad1e8zHbIp732LetTKVdq8fiirwgTM0KpoyUPnhtou
Vl/KoY9+e6lelNLPbPZTDy0jfpI9tnfZAF/LIWTxynqcSVFK/57qYhGt4b4xfKGpMbTHwQ6z1BD+
6gxSYirjZyxQaQFJiUODXXRB0WmHOg+JEmt/eQegQtiaoqYneN/ap3jXfBgf82JqF21r15+G4ihT
/ElXPzt1BlVD9+yKBmbQQLGtglfR0T8rjqTrHGVfQQuq5QvRVaIzhlalM8OEZj7MGKmRkqxveU0W
TXsKvATZMvgiiTkkpTserBsP5IXorTCmKlFJm7f7oOmYdhFtUmXyww+OXBhJVdBAh+oHJSgFt4g3
RhwmpAvMjtTCsmAHt3x/aHs5HDWRiCzfR/L/X1x751CV+TeoQTBGgxww4z+vywVtNgFZF9X8D7eN
x+PbOi+u8F75SjfVaxmFUTcT2YCFkXLqLzx3qa4RXiuiTpMq+rJ6NN9HJhIoVv14Df2cKuhQL//A
b96uybWumFZSj95ijAsVrmrxsocOwYx71aMjIr6EN3krpK38rG1lp3raTd0GrTeaGOV7GgV7h5vZ
YZMUYcDkFYte/ywZd1jthAik5ARBjlozwDp0rdpK8v5hxrzuEZuYi1OtNI+HQuWyjMsQ2bePEVPO
oORf5ZbX0w5Ncn+v0bal1EJ9i4LNUE0PlDrLWRHthJ2iicsL32qeqfCnXVjG+0JCsc+xv6bxegJ1
XoG8JTvwz10vi7EXcWLUIyRIEGb3mxthozedjvZxKYnmwxEaRrrGhL4u3I3+MYwX83I0MA8/uI6U
oPNYwK10B6a0AE3MoTOZAIhLNXan8WA1+SNw6rZ2Mw041PwEIEksq8jT6tQUd75pS+zkP2AlmXDD
ZuJ19L2cwod5r3MgZmMd6yGJDDXPdynzIJeEZEEuhyFQSQTenv8f01DHXcHT+UVfn85ONhbqTzyN
PO1RxkLW0ltcWs1Dc2t5nMYHzpjhdksSJmEjj7yHYFc/his6jHwDdOSs9tKmITMwLD3rf/CL1Wj+
rYBl3iOy98MlF78pysr6F3v4KomNA4fNF6uf1IiACc9jjvlC54tq3W4BbNv2+MGDtwWiXrqc56+A
J03AciNSiaplnYqWw814z5s+wR5p8JbPHm4+JV5N4YMKpd31WJuWBzuEGgNMjFtU1e9fyRseHXXh
p0bYfpWC5JEKvGbjx+mKlA5aJz4duKWL4YqDIsQTN6vBb60PUqKrD9zIihPP55FrEej+eR44Y5aU
w94UwBPVIurWlTEv/Z3Zf8DWpuJhF1B+IjBnRFSoU8ax8Lno264/hJsGmp0IKiO6R2tjGL/UIl3J
zh56vkNeHCmyoFuCH1lswUM+Rs5XAbalgAdfr7Mj6z1J3AcOuTPDcwmIQw0HShnv7mMxS7xtbtm3
l+wfm7u4wmtXAvfbYwQLUwiXTqkkYwQHkYjlJQZy+nIIbB6PSjRPEIKk5WZpVNeE6re+1HohU22r
BFWL9MA96qKB5oT59aALI1mK5IkZaLT9xZR48TlSSFKDn19JbkzcOZiwp7+kjl3z8br8xl2sou8j
j9B2gIHkrctR3uPMLmbS2UP+6+k3vgqZvwwkGTT/ND3CCibGETRxw8Rxl/lGMxN50+kkrpCsJiM+
tFOAP218z5guFEp0fCxEs4dBa0v3RFxUn7bTF7vOrxxllGxo+j/OOKPMWhAMA3onzqfOyBlEH6rR
xLPI1+hOB0FdSDVPth0IpsCML4QKWp4z5GtKi2Bq5FerifPB7rdfp//9EuXkwWmkNq9JvrzTg2H1
afc86PK+mma8MlA2PkzuLhbjNt+5dvB2DUS0WGE+8tHfOOiR0RmMM1lPnFC36vRzl80HJcZK/hXk
CtlfAmed12hwM2o/VJkES/BxV9PGVVrqW1XZiUBLAS8t4+KHHAHAJTnFeHgKv4vGolzRm0t6WFec
x73kbaxac6P7099c63HxGv2B8lMQ+opOtoAYMcesGJ9LRIOcx7QxO7uXYi0W0TEGYufkb/dcRaye
CGo9ZNZYYDaEFJafuN2oQUF6Kj0ZNQDr+iHJXJb0gAPEoK8WMaQqx+E1derlB0FBThmxy1zanCE1
Cs9lShPKQ5D+jwX3kXJIoDHcOqwzsEt1X7+onrcEBkdtw+oSyokfeiKIA0l/p5eX8vXq+Nq3CGCx
WjGb5nYYpUQTSXtkhfIc8+taSkxLDChCoOzZvnIKi7XJpI4q3qSGBvc6Snig+JUyPxxze3YhKeA7
3bWifpoACIr3NHXeA+b4x9SrdlkjOgLZ6w8YSNcjT7B3PeW51PY74Ic7KKF/8DMeBZRN9eTsm0GB
Yw24Qx0IKwqb5I1Gcw74usAxnNPzZTlc/dxRiu5pPSUmBcsKDnkXm8/kPm4DlUmW5/akeKS4fVjH
4j+HEYq6zlHF/9nL6ptGYI+Cr9E795wZ1c0cy8/fzTP/zgiBicwuZBGyUvtrIhvp3n46PNpDJSa3
g3/VpqOGD5+7eOBkEvps2rZrwoPwH889Yb3oCqlbyfwDyXEIQ8f+cnoWK7GQjVfRjhSGep2zI4BF
f0XHcTIhk6kPhEzcEu3eTM1PMIF0uY8BJkVPiRsLDpcEb4prEi9dE2m61HkPebY9JXuE2ZOqhxPZ
HpTCz7Xu80URTYaCXHwqrHAADW4Unbrw6KoN1blKxBLY6CTbPNieLvPRtX7wrTHTkxPNXp05R7nj
nsUhCTLZ34qK2CtyR0O18RIdYYknR3Tzk6FAfH0eNKNggAkiYvqvOj7VkAo1+zo/+mno1ke7fLvQ
+qlZ9FHPMBK7jxD9pcAdk/SbA56kWM5KeEu8du3nFAJn4QPztRttV5L4WvFCjtcyed53VnGwziqh
n8NDabSOwXMS/vlecngAe6OJLIXO1wBbDOvRZGQHUUhtCOjYU5wJ54xJ+kdU2jqbNI7gc7+I2JOY
tekZiQn5DgNb4oDCJaNFUGnxIEWZjpu9WMr4mIQZ0Gs2ncM4S5G4Lb95bKvoA+bafQ84XvU5Dxco
6HX40cM4GufG4DL8bkf7DxoTRuDVVQsKDvXyRxndr7kpY5DSeWigaEIlSW0IMVy5JzlEjswwNRB2
4sVqkAH8kcGtrm8SkhqfV2LZI5zJgKL//TsQmlQcTh8hoe1Pa0xUr1yjPO5vl39NjpwtLrM60mfT
H4FOcOsapTD+TiY25MsBZxP8I7z0YO0Oq/tvDLCaLaRAVHN3UtcnbTQPjwE0CbJMxnYJYZuLCO8X
iNj92EPxDLpQ91cp5HNGdv/TH0SosNlitzAFHXd/ryahQubuqRXy3yI/3NNEenOlsM8kOO/xBBn7
89I5lNDsaLd6C2qe3nX2iBNn/o4HK2ePz1xps/rdoeP7ZEQ2pf4IqpZANf81DFv/UsuWUwbvJnZg
xEPRIT0yZ+AM2/p5bDVL/b8SfjRQMHbNLWQRITcs0HwHxMFvkmdXbQwHdGPi/xg1PJBjlwl1poOJ
vzGPnXPA7O67IRoKjm6X9HZxGvpKCoHWTXnoFgmf/wNYLI28nMH/tsFwjZjmslPqjSPUHyB6NhQv
FgmY2cqxUoJqQVb33oiiv4Yzmb2llRTVllCkpIoJ1fUgPycRSagQVwWFm0S77AzyDywd8Gp5pjkZ
vNO6UxNOYALNCV2Pbn9dSSDtG+dJZRQzUNbIfi9gRhRKkLAQtoMHrNrdnKjNAHE0HRw4oIKIjpjl
rWeok86jkT3AS2jx2Vw8ts6UQhseW16wPnuJMNBLRxHdRg/HooEY6wAWmGO9ZvWoSr3F1XCvdys3
/qENBWvfRX+b3Gm5RGox1SWMMEtFJijePZWp303HbJyd7xNqbtkhBM/2xaxffAKPzAja64iuDs07
8Fl/vZlC1DyzruLzawdJvbbfRsAV1tOLEMPwlZjJxmgL2ibGJlMFrJEnJGgsKDip5Lpn7bhGJCUK
eHtuJcS6dnQkXXDFlsQM5YWkbXTsDhWVj9fL12swsZjksWr60hdltP076v8Y/QxHQK0cVxysxpNr
UM9/VDZtjeX8ilx6DVPGVULZjqgbSebWq1xWEYrAHJ8Wkdn6oXH+TvCwrgsqXlW/2wA2nVChDhJ6
tb2X7woXMcqLb2i9QlYcA3jAsb0HrOxu4EGh93+tepmpG63uebwwMl2d5x22ZAFEpD2fOoQeoLsM
ul5111Uw/SeMQKhNfYorv4F7ofVqVYsp/khgCn+f48hFoJgN8DjRjc7m5Z+aNeodvBhALLECvodO
gAx5ybbSmPJrJoG/bH66vRXVrRz7E9cNw+MTIerRcT7LFjoCsu4elGoPtdmxFQ5KXcsuJAJOW0Uw
VykoXrpGie1+T+DAaor/yfaJa4EPXa1y0NGyp8BdKFdTv9s/qOaC9RDgW9tphDWQlJ7DwQrjZhbh
DpCvy71DAo1ZmZ1DL6mvdFv8RBR20kAQwapbmxDWCkqyFT8S+lOq5ymcacIHnqDdSlb1eJTC6UFO
rpKmXcrna05OtddvUWm3WeUG7dsA3ZukZHfg5jlQxyyHDy8vwfykcexSGcNrEGWQZ8GxHwgdo45v
Fwr8WXBfTs9VSGR/t1ZXOIDjth2+ExLJKEn2hX4eN/7FSmcpwSYx5Yx9qUCXKQDlP7vx6BL14IqX
QBrWWM8hEeX/Or8WBK0FPvLWyR6gC20yCrNJ/x+n9dexoCJo9lQs/zmdQv86m2RB3YQB7UoGIVq+
vfL3XIEEcg/ZChOQMXsxGFXsvDLeDr0sutr1dRvqDlHet/CTE2vOmcHEOW+3Ish05GQwsBNfb8T+
hJtumJcQn3jh5IuQpAgaYXUx7xnjf6dggGDlqlhQUzxqNCP9T4nQtx5P7bBlHzRIQ9JlBIlTKJPY
io99PKfMpy5m2YWjttANjfJFHxwPh3GwIDS9GibhBJyLjQsOOseNuXM8rwhkMJMWdpWgusbhUJKR
0StOrMCN4x50auIPDZKmyA5p3ez2F+kQRUNx44yrHZkbsbXdmtP0dZPZ1RpUTfTUATWG/Ep0ezYb
ik0E98wEP+o1Yd+wb50MvrAoctT7Cq6bYIEU/RYRldZPR3eqyEctSZa10w90B4hHd3rSW8FfsoRd
zNXxAc7kUFowCTTEkXx7nEI4XGclRrWxpQoXhmn1UQtKPwIJUc7/D5pAzL7dPOYoCtWB/CGrI0DF
YoqixhyHukVe6dxUVqB6igUQA2J6kMyESY+X7B8UuIazydJ80u3yVhuAEDT2P1OV1iE3W4BTCzRr
WGvOYRe9Hg52O4E7k0NsuXcTOf52d68H9OlTWgCBHfslJXi77NW2ZyuqEqLdBUIuCQLpP6ttH+eU
3v6jeYV0VZtLBTFA816dpXRBl+8l6wrNwCGAeLR44Co9xY2/CDFvdp8AAu/XR8gssjtsR+1Rimrb
skzV0WBq9kFnQ90/JSZl21UcdtNleOxEnC6bNkunEmWBRdyrjmNzZAVhY7EywqzOp87Qi698P96B
6XBtpbUvq8erWAvEJN0CeLDMOcrK1zNkgbZ3VHwxNOGHhqQkbDK7AnPBbwovtEy5o6rw5m/S0MZN
LPL3nDXsck8cl03f6mdr9QgSluiPkGC7v53lqtzokVWT2jfGxDlhOsB/LW4y6RtagiHF35wt3gBs
vuHf/LXLng5Gu3Eelab+cPqn+EAy6Ve5UoBTymrHdh2s20tSjEF5ti8J1J6AcM/p2hirCa81Xpw5
hFUhrhRMcUhcHD6sp3gsJ7kDN5Br5yJnGUotKxZAcabn5gE6QmkbYmQBveQ+i6livKv4BWMhtbuw
794JPo5muruxMP76owSOir5PqpBNr3PixVfOHS4sL8+ty+0pmNZlBioPtHO0fpuRzanvLsTYnpjF
Y5fiiKzLaHfBwxfAjKvly3eiS5sPWXecEB/OQ8zUn0iLCpbEiI8nFZtZsEI/euE95R6SRmjCHSFw
zs86l5+CwBQSz1LH26rnLDt6GZ68jvnuPo9q82D6C/PDb7j70UCUPRRZxCp7a/NQctHeIlLhpy80
FJjQhJwaB4qxBiRXt8fuHmwZM84XeK+Uw6clgrcg+hQJJUCwLmJSJ12j0fevs/t0cVcGdOh7FHXC
g8bUsdVYQNLvycgPKHlIzCANoBlmLHLqGuZylTWFPmgTUeJwG60yfHlC2THiQLwgetSqNyDzPwJS
e0YwitoJXV+q04LyhsPELMvNYnOyV8jsgB29rXsd4LxziZIjFeLNSa+u+pANzrGgbJeuDjnxVo3Z
+ea7zn+wRONBimtGhuGCpRY49/msPn1yAx04Bj7PBAXlLN8AJavGIiOLbxhAIKGEvBXlSEX36t6C
bBON67SdD+ww0z9f8U9c5Hodb1ej7QVUAtmifivTD7a+gTipGP00bUjSObRWrUCMDhPznJ0unSpL
IorPTAwvJYYeyeE6Fn2QBy7PE2CdIBMe1d0zPUkGP08opeXrXpnHbtjB8c3RCg8fpbR+60Q8D33X
jp5lDttwxkyLzATgPdhThXu6A1vhScMabgccT4HUd4V0VdXVTkVRw7xHk/7ky+QMPP55/Dg9WPRC
APsC6jG79nCGJWKgpBbqEeNwjRPxLW5jEmNH0e5p2Z8uCo4LuH9WuMXF0fYM1YHwkgSIhO2Q4JU/
SgUhKOzS8DfkeAOGptOAfw7oo17CEnP//QAhgUCxpU9HrAFk89bfRS8TyXIr2P+Ep1OUwrmzGaBD
9vAkPr80qa6X4t9gTddc0YYQf/2n144w0rrLgf6d1psSPRBA/6vkDlFeAVmwYtqINZzHsZ8VBioX
qYul2X09+R6B2xljph4FpPfYublqsCwI2Ew3/ww29wOiBI3w7CU0qPLe3VeYh1r54JkGnq5NJ7d6
7rvFZ0kjjeFXvDLGeDuDK0KIvw2bQnsh3KdcEhtNPEjvPm7QhCTA64xwJre5mzv2iV6NYHs0zLSj
ZM5F03V0qiuVDxhRbZUhlAU2wIXahXWtVnAtSKCMxXPX7ugpdUXQ+kClWjb3iQ/P393+OOLzHBXi
sRuk3IM9lCeDr+d7VwH+bKoczw/VgYz/R0Fl56feBDzAX+ca98z80gS1EcswJ1gA0nyDfzgNBdaP
qr5e1f4BTxwZOn5JRkymFdzBumUL4KPFHARVzj6r91AwxCvOxy2NrNYZ5z8V7GfQi7IB3xJvGe2J
9Y1MZ2cWAOa2984Qcx5EwahmhjiYGyr1Y51Kh25K8SAvQadlKCskMgMBtQtqWW4Zy1wVex59JUei
jIHCHeP/DQay1ZluwuYZlLBJVXiNnk5BkCtCxpzynaMTmJUPv+gH/LAKqI4HDKerTbztvlQrzHWL
soDXXvLrRroZJgAmRpvoDNG27OPbWlv1PYaewOdG1kzPrxvsBiDNnbA+WnZB1bAdsjPbsy5lUl1O
hBx6aPMdV5neqpyMteWZm2nBQJCTFKP0U2h/dU5zV3lXxdX2/9K3i7cT67zlIFwVh+n/cowBGfaz
WKhvZEkm8wokZeJyTwYtDGZ4kZL3Nir0gZXy8OwXv2ijJphmtiLmxgnfOJ53GeLNR+bGJ5SXHIhl
2hQHimt4vj1KGDdhHa0Pk8kUFmQVnIVc04EntdHlulMlTINRfv2+PWdowCO1rD2ReWzCHNRqfMlE
SrkdNKaIEnr9M5UlXgztHQcldyoMpGesuYFGFkL3zBP+KK8PriFd80/xu1wVIKJkUta3QaEeusgm
EL8KX+3hQi1NzbpbXxu60dVsNj0313g9rzJtFhP3b7mVH78dqsf6nFAKgJR/NNzC4NrObt6jmSpO
mPZul0eT9RcUY2o42QyV9v1rbrz8l5Xjj+sN2rvkPgFpWY/cqTzoUQYZIwm/e/84WozWllQrVkoR
vTGpJxRjyOferBJc/1XAMuSMjzJascEN6p7lqsErvlgH8o3JyRcBYjrzP8+C5utZ6sOS/1oB1lK6
FVrpsEM9PCWl3I22AATDSqkQ5R39dDzp0IZb1g2NVbtrWAxw8VB2hZDEZGfH5n0RbKe901mBJz14
zGldrZcegi6QMX/4C+eTedWzOBW3cJ8tSjMNsPMfxHKOT+V2B0zbMOiDhdU7yklbd32GXMlGcl2v
bMZy0jD6GVoRv4qunrgBAeRDiOE4XEwjeCbYppZkKf0VpcVaezRC4/Q8rRqyrIZMcpSG7ZNG5dGZ
03b6+clUbJkea6em7Krd5L/2kbU0p9hXmSzQRGeHhzJsb8E1uJjMtC+JHMmRHXpsBXjlNe2ARtpI
SgFkCGnQ+kCSUeL2rTlVZRGm7HxXLKOAKjhItUvbHJoulpt+e8h2QVQJUkWvqrgm1e2Tp/askUPX
Q2a7Ri3w2sdHlnE3YQUtLA3+x40KQosCVM1FdC0t/y3C4X1QhrKzhBQ3kORGTDpNJQVhEEuezA3p
miqqCtlYkF78acCa8nFefTpAReDMELQWuwUQumyhkHHOgKi2L4MuFzBQoh9XCoCvd2Y+fJCXt9JM
NGp7bC0MOhXvLr5RbrZw2V4hTpxczbB70F1LyigZUSYWKO/QendnP3YItUIlafwGKLn3x9Y22ped
uudxM+3ZXh+Hsim2dIRFINuGNbkkhUS4720D6j8cPdvF1iHi3hfG6NPh/KB4myPXZ6+jpB/LKoE2
Bb9R7dnGW7y5/TSoPvrNrjXrnkl0zHxVpeWCxoYkDk9wZs+YCyjZoUbdggvjyOUekI3T66yJZecG
wELiQdjiFD/HPSmnjh2LpZK0+4IMBNPhe8t5oMuO6ZmrwrmHEbJ5k2B6w/cQxwuyAD8qIxBE6Zo1
y/B2/q6nFRReZfXwyX71TrQ3fzkoAcKbDTMKbkBWS1ghQdojXdFreEJYt13x2SL8NdwTtZRmjx+x
3Fdg9TkapEpmmcm9sUHQIEDaoGHcA5Hkb/6vVG8LBxLvZWqgABgH9HVT2fkgVbqzJFEzISRvIx2w
l0RzbFJMnscB9UxxgKQwU7YHeuCVAHwOfHsOoS/uVyH7E7bQ8+D/cP59NtM8KUw3WsLfv6+PQwIh
P2FxgPtnUWpzruG6MOFUpBxUWQeDm4XZ6RvRcE14FkFgSMLMPllEE8ngpQpbd9HjHbSjgwldnY0E
hd6OHnVRRvK5iW7tpuZWe00jglRdQbUm0NwR5ybThwFFyZOApuH9DN0qdVUu9Mminkh+pYs1J1w1
QT2KTtcT+5RaDudP1c6xlPhQ6nwRhtptwPQIcTR8/3UiMJccQ51V2xcbS7SLzCwHQXVUO3qwldMP
y6qBJjhbPdzJQk9Xsp03hIXBEtFVdOlsjGKvED9prQCiVyOzMuI1oxTxxbRQkliAYWq1HzzT26ks
DaydaZQqaPuUAbT5Q7W6QIdP18bfhMOhMr4fFowdMPsZCTCHLJ3SUB2qrW6t4jM9IMJGIRJvTvnX
vYNagpnEnr5VA0qiVD+O05AFEDfKEQ7WsuyMmKzz1heqaZhuthg3UkIxZrFDgIWIhGltAhDiQNnU
u6m4bOAV17coWWYcCP4HnBKhd2bnUQfpo1K4YsPOCOm6rDiIYNCBFa4A/ZRyrMMGRNA3XLKJ6W+2
hf98S26PwhDTkO+BU2eT4NnjVbWFnYuh/0MDK0AUtSCUIOzqwBfte8LdOson0qWAj2tOoOahJK21
4DYif7URy6Dhc1o0oeAjT0xJzn5370iOIQ64r13KdeoD/j949N4y+AXhJaHs4ThLlo3uZF+EWSoU
OGBXFvhKQmOsVM2ZHb4btk7CPN+36xL2pKHXIEKGK4nyrkGx3jnS7Sbs/MilOvHxpSEwKIQoxSsj
zoRW6I2ZRBw8709G6yaSb+Pd081wxEV4gEF8Uux8ChPAhe2uKpFG3x4N+Av4g08IsJzoChJCnOZP
4J63rtGIM6Pgg+5X7uEDgtsPb1M1Yr7w078XJgCEQHus2kRDRyXBATEZKIxIsZQYx2+Ihly964lo
l0miiRfBuY9zwHNw6v9tejdelMjqdWaLtsrF2gz/NJQc3mTIHdn7jFtpKhrfsGNbwoMBY8DmoLO5
Q9/TwaSvpTwyrm9SfMknq/HtnlBGSsNmarjdmD2mnfjnOAZfZYTLJ6ihaA4AeED/HgLZZoKWJbiC
siFW0ycY+0uaknpqNd++4NaZ0hNlFTiP1C+X2RxtixKsgp/GVNbCDq/c9J0HVHdOFwPkKPC0xpW6
SbZqDc1pq/EBZ23WnaOfpfNnXK22L7H3jlKzfpNHupqiZlXvKy8AGCtWU7c8WlYGgtf7njJ+KaT8
hJsz9alBwtm/xW7HBD8g8on3rzrhaWgz3FWjtfW6tfyozQ9zNISDo5gLeoayhBPj1jWusUwPAB2l
n1m10bfi8sWrHgDb9/aRVcyJelSJd+rXP9wQyOSzbnKHbbCEFDGhkIHbGxSWAQXiZgo/GPkoEURL
6X0qcayfMe7WUCb5tz7a4EuZCtz4ZVIDVvABI+JTnK1/7In2JTRgylpowOP+cedqAkShfA+ksnw0
ZVvIhyGVeX3zeLulCAT8q2yG2ivr2XkI3VeVX1+lQdAQKREOe6227jvUVQrFzaAAfkCy/Wg/imTH
V2SCabLUYKgNOSHeFWwTAIgefB5IKHrl4Mu+P4l1LJfctfe41nzQ67eXW6GCUwW+B1xWu6CJQG7Y
qPUCqQt/vBVMzIfd5Maj2Z2Gsg4Pia65Nd6JQT3EwMDnU+10+AxcxSSYLRGL+2ExWJW4e14RLRpD
nki2jguwnUQn9yegPU7+uNy1rNcwVkiPExsP5QiSlLgafPUPyfIAUFwh8uKzMRuC2E94hriIsT5m
83Vhnc8O15FyfGERCMpCAgTAyzdrT2iKlN8z0Hr97Boj2i0/CoCTOAtjmpNZOm6oplCOh9CL2tj8
U340m5dH3tmF54XSHc6L9Oppfm0FTkzUCE8H+dhq+yBOfa8706egaIKgvcuYp5XQ1m3kfFpc1AMS
HdnJoicXPNkh+iU8Gp/mMHDwv60oPh67b0X77Wnpo9w002c6iLsJSt9qUb/oNeuzKWwYgmdAR/Eu
PmnsduP3vqajAnlAzbmRxfQ2bmlCKuTV3RDpPy0Ee8LEPKh/gOypP2u/OqQpkPeJ6XhdrXv2qukv
prkxetIjYYkD801Gv6sd6SlqupWHymJ9rawXaspazUkZrSs4gQmnZ9RujKf5Ov+Kxv3YDv+MXOSJ
b/f/J4+R5aTfu6XQxkMOcY6Q0C72lo6K8RAybI1ol2TGjA/BHFaXDykKnWbHewWXgvuUaB2ZCjcp
5RmYaCwVQOOxXzBVlCix33WGX56xo3+P1G+8wMwEdMWW+4qnwhIzjd42FD2cvOT+pUUL/bBgU04N
6CgQXDFcuB7V83RoqhgwbyGDE0rIy7mUEwbQbu7eo/q70xx1s6oDGU6G5k07quqzxlZcVuXQ4f7Z
e2BrqSqQ50VNnsZ7VBB18KXXgT3GgfPo/1VHdCgWgjom10Ny179+v0fh/VEDoyDW0KOS4HcWHjPm
ozUH22YZBvwrunl5QEYzPGZ4mWLKo7zJIXLxFe+3QBYUnNIw7k90MraVwiLXPotfI6DYDMrrR4zf
niOh+dfaK/2npvALjGt3BUFk004S5YpuZ9yoonMZemuQ0NroacvFONtr6SCUcT4L92eg6XNR2JF6
U07J4xxDNbo2DRds1sqnSF25n8gBPJ5ddu7hy+L4abyXP+wkxPgtn8i3cvbOQ2egEZ3hFN//YFt9
Hr0HsIn9u0LJS8eY4FP95/dJ7JnU+nBdWfK6dqVrnnv+nB2Qpc25UGGpJDWp+yIDLWBj8sOTHfOk
Y2/eTTJa8sWPsfjH4mrGlsbWCA+akSs2tyJVPVmk16SvXA3v+IfpKf561t8Wl3/dIaO5czzJ/k18
8BVuqSRsEPLSK0mi8YSuy7YzD8OZevMP0U+wwGUd02SrXakeUsnRyUumpauRfvmMDmWuWAvX9MnS
8/aRIufmIe9PgCTOmW3mPmQP8DnR0RcBKoJo0yVYUr81mNcYy9OYYSFrVIKkTTc2Epho/WWeFPzf
gE4A6yQGJqkjzC8IrqccoOC7dTX8Hzey6wJ5ICDNAYzaEI8F4WANqJKCnefp7ILpa4Zb4SwVJATb
gn1vtcsi4svdBfp33/AlZHS175zCLZ+6bVQqTCZOLK0TzzBt1Sl505Pmh7R9hNsT//SsOHs+9V1C
6wCu37AFtsk0HXlTmFbzYZo/RDug3+1vC7K+J3n8rMTTuRqIl1Lt0pSAOnBqI+2KB3ZqkrUchP/r
Smv18yl4iO+8JhanwBE2IVi4P5PdaVdYTaio09FUbF4TdHgZiWIKRznSqfoKt2jzHa/zXytetyl4
rlrhnj2yIJxGxrvOLVjNMpoh7pDy4T8kes6kxt8uQGG5tIaffIEKOq6C5/YhP0gFpcQZ4GdvkSnE
b0cfKrmxKGJCUaH7ukUVgMmrOTqRmnFz9oYMAAntpqWiEj84zPZxSawtuWpmG8odUGKA5X1Y6ryB
5eF/XxOCrh2dFQOg3CIyEHZZ6mO7LJ+CzqHnKy6TLiwjwJzuENIMev2psrBvD/PTWuNZ5KdCWPCH
5Zd+jHhftOX12AJ+pQLMFjl/ecUXqElOqCiRAagHqFb6xv5p9j2R8fd0YuyBiIc/JQJa2+CJWY0g
40xUPOaxbTJ4xrq7ijxwLsCjnpTtaxMx5cEWZrxqo7jWIq/LVdkcTX2khNUz8gaJL5gO9GBbKxxs
ao6OINFeSWvBfQ7H9ohOL/H4ha0BG/IYjT3KxkFjxX7s+k7sIBYHMH78Bhcb9O0mTUrWMk6PqgKp
eGX4RyZRaPHiXPwx/1NpD8NF2Yka6y4+rEo7AQWuWs5owveMq3MIEbqF1KUfCwZ3KVf+PCUWzDWQ
LBEhWjJAkIQtxjk6PzULfJNUIsXIRJqmztYsMtfy/Xtbrwx0wx5qauL+txVuOrDsJ/iD1gGwAZYz
OhR+1Muioye5QuIg6qfD2htu7QUliJ8qnl/4G27lQ9Q9N7kKtWqRywxIS9ULLUGCHXaiYcl85O9S
eH17VgwJKU/kyaa+NTR5DDDQkGa2ISRyZcdQw3OsOGjwvWViEbT8+pMwXfC+lVFWyz35BTSIteuA
KVOpl7iGHHhfJC2/zqpTkvEWJUwtw59/JWpWvR/EnXdT9kdIcGx6q1FF6zpG+FzRN+GnF9KPjD6I
T0o5hANtWTe7269YKMdN6hwXmhvLcwmyod9YpZ5AdPhkaZjc9qU8S1G4hIuB0IFIc2n0CAhBE7Z0
kgIaHbwmZMZ7ZN12GP1TIZfcIOwBZnk21KaWB6HNhYRUBbxem6iLmprFy2dchUwEvjNAnlRyKI1k
rNR3fEl0jOMmZVyXRl7z1Xzm7t57+B/qmoDvD8qRukN4czomhze7KBbfsBWX07rdJAZ0XmtWtLxE
aHpobcPfeBHj0YHRvmpYG9uaT16hrSr30uVj+cYin1bYqFu0HKyaeOVp2NwBY4Ue8Gwn2Nc+PxBr
naHlp+65sjwcaNsC73NyxBcistIzJJzaa4n0fzG9qws4LB2wCth2LjXizxOq7KXApK7FaYNpXrN5
7sD9woBrGjNVQcouu+/QelbRZH/05OwRdpbFC0h8ab8G1AIrRXOpCN0Q4PfaGPD/dNdPBlRqYPB+
59zRQKb5MXu3Uv2gh3B1m4vGlaEJhwuICULOo/2Ha71GpwyQSrx+dd/uOh/UFU7ljL8xFTZ6YG+p
w4Hc9lj8srDvS5tuP4b6oAqEwfc2YwjJVDkwu8kEFZSRoJoMb4YdQimN0nknUNJNgCZevYnxC3hO
36IFSEk3FkLxYY7kLV7sBPIDeyXtiA4CO5HQ/tnZ9qh8inXqIN3cBxx5bKWvxliWZ0hYLP0W/18d
XCdy2CcJOZTy80L+rp7rFRU3qVVCyK/zVpXkRm8hvMqMVvjioHZR4hbM9qGWXUeGCmp2LcuT5Fv9
8cngO6Q3E+TlSMdu+71PrgPS5k7GpC4qChHmuxYviapBolhNkA6p7eXiLwX0ry8gCqoRXU5QqsMx
5t5dMvy6FAMxcH9zmVO1JLkgjXjEpdgiv6n3XsLkUoi5+TYNMmt0pqzsnXjF7hp4JfhMnqqAMn19
qmtpb7/ZNZpVn3gB1vkerCV8Sf1cebK3ITVhNDqSuz1QC0mUVCOPC32cpbkWaqgXVVwB9aT23NGj
GkIGRPWPnRDmXufrbBiu8ogf5imhTepq4uvYKGrjeAK1qCbu/bLWH5W0MYjMBLtQtI2ZWnKUTycb
Aoshi219PONChR1fR0byuqTPCYneP7Hd5N4BXDlol53ZrgiW5XgOPFbhvVJrrBIOxDagynBBRFWu
SQzg3MUPTjruzJqXKK01SCCXAsTq1hQ121kDv03tb6zMyAChGrQk7YGmYNghN1+1diUGJkLaui3+
NWsUtKL7Cnldsp2YU+C4L25hC/YUEw7F2/H612enqYNe7+/UFicQCa5X6GryDelQBnNGq8ArYUzT
NLBYRNqmwKuzmvLAnfR5TPYPWlbgdO0tc8fRCeDpLmILRwy4XKkxgvEPn8PG6YAv0zIMPVFMo4Ww
Te8O+D+mHm5Kfed1UDwpSrbWSj0I9IehCHVytpMUFHmFZsjtZz91mu2vLu1hUuDB57wab9JcBSy/
adedbVZzjnIHoTJPLe6kVVDT92KATtgmAZv7hSrpNjE3ftwSXSfNXucYty+Vz6NI6+rvdMsvWXhU
TpsrtfXMZIekK7t2yHx7lOfaAHOfvjpthOwhbF0pO8SnxOdUdBIGCYNHe6ISWatzgA6a8qjsjehs
LuS+nrK7jPn7RTcdRe4qVK2Qojsku+SdAzZMUmW/lNZi2odCuwYVwyGZ/NEfkObG3vU1cv2xivUm
3TVOc9aaYLtukShrBzQcFOrs2lcFKS6imDHfCJ6b5VVRtF5M5kz5RO5zHPO/myIASa4mkDc9pdz0
vBhYqrMAbXq7ZKwrZRkwgWfOuyK1WkS2+RvF0ku2EtZfQb5tyfqgFIcEuGNSQeBPBwJb4kQL6mqi
2+HTklYz6nois2+MxSiXA7fSWX7eaqLNiQj0QNNhfiMw4BNQeZIvPSumPbIdtU80k0CDSgT5Xdvd
PsFI0xr3JYEdQci1pjdaG+Iy9aItosxeL8jgfp9KYMODQ/v7jMb1o/LDFEks2K6wT2MEDxoyPqjV
SVPUbEn8xO3QZzhvHhuXQ1GLqb5vcwpfZ0IW0kRUx+1vIDH7+zLFdWcAIndkyy7luySZdlPk3uRx
Bp+Tiebey9YwRl3j17iWlzEngMPupgFthEq7IhaN0jFUM5ZIKRHxfoB9m0/pnOhKRNCFsMY6//J4
eL7gFd7hEx1X49WgKXP5z4UTZg6NMH4UQrSwPVaGvYyyGwd2We4XUBFnBtI8Xl64cwLsbOjr06vX
3K9iN3RsL5FCDDiCevdiIPDULrwpiIxbdQYgDT4FDsru0hRxUX8Prn0poTSb4PTfqRwT6zuJGZw9
51VKtEmUR/Rx+6t/JOUaLr+HxhSN3WuINI6A9tmCbRIP5F9x/vC6ZU8A5E62257PQgdSbC9Rnk7H
a/E7l0u3P9YzfUbBNWaTbKeHMMVgI+nMzZxB3yOXPRSO24Bo9qkDUZ4iwESAFrkvlG4o5k4AjbjA
9kjolSztMSHi0ZS/ep7TIL2+1UW5oGP4voSPhQpNobir9zP2lZHJDlGn8G8wkAzK9j9ZDbNyxfVg
xT03mPfVAuDtAY7/wI0djOUFnjUyAalJOrOR8hMAOh8W6swN0zbOyearbzZ4raBsTOaurY+BGCjR
iKPUHkJtKk7297UtgVTHYlT/ISfbIXhzHFCtc7SXiNSEX2yGmcdgu4EXb6M4kjj0rsSu8PTegCQh
WGyg4zKB2k0qnhtftKwbQ9tdlQqJ5yNZVXOj7/Kn+o1z9V4+DSRCIt5XG9jS1q293+89TAi3NLtP
IalDWW7k9xfub/pQI9MXexQwwe9lhapGokLWt1PuvNKyqSa8sxIG3y98fKvcVn94NBR1XNEqzKFk
riN92ruc+Y8N5Ia27Ykjky8tkuA9Z30uAIJ+aVfgmNxPrc+FyEN0h9mSKT9mCl3jPHp+MBJVzClt
vwWzbePGtcaWP7mPt0VB5rDURHetDNe+bqIiYVQX14sviCp1Vr0iWE5BFWbt7rnq4nEKpoUhlw1I
8jsvXdG9JvPaOq9hROFnkGiBB5x5QekrqbgOM1WLw+pMTEuiHDbY5kSFCYmRdgVTSycLTxrQHpHz
hqh23sBKqxIQ71yxeEn+flQhcJtLiLATottHzBXOoNvcKPQ4vcxAiBOEZIBXOG0bG9ZZKl3wThTc
ymvLDHiHHbmcoQvNzXkjcGohZnMeUDAzVS2s399z8SRJDXttxmlvpgii8U6pCHVIXRxMPbAgeBUl
TdC+H6zt63srBQakRaWpIYMn2P8j/7AEsxRW93rhf7CwyA6drEdG+MaSw57bgVtztH5WnY+o2ySW
aXD9iKATTHFhJCMWnzpQHDt4ndpKdXKdsdOyaXZmNPYbbVguDdhh/FOy1fiwsJcB5W9PLL2Y2Kec
6ylxe6xD+wn1vxoTXnYIbsNH1ruN8He+y/K+seEnrG4nNynp/UHbO6NrC5VIIZUCT/VgXrkToVPk
Ns5eY2QuoiIAbQtSKHAz5jh+7zqkG9ZQrzgxDuPRtGYNQb4BxvfQhosXkiAgwt7FzQu7pfB40m5N
p7Y1cRGYHPipkAZpDRbAEPg5Yj/eicoZ5ppiPQz0DNx0cfWOx3JF+13XggPzZMm7cXmpTQta/n7Z
fdt9ryhyUlIKdvJ+0np2YpAWc/49CMRSvC5pQlNgFZFPkGdvzyxkSentlnfWsUSu9wKIZW6FptGZ
Wxrb69wbXXS4n1r5paoldpy5E4WqEZSWC7MoDuI1p9VPI7ZcROhHsSECZlFEGUtqcGJRuun1OGZ0
cPFloQ/JB377LC7EypHN8QLBc/rhd1vo9FhTFhlKQKO4jhDRkxc/sNe8BgpLaqGOcE3j6xWJGuY1
qfB+RBk5oIZeGEnf1D3GlKa6Ag2M6K0KVuPOA06d9tK0EfwiSbPT4pMKM0ATY0vtMPQDufotN8Ic
LoUjK4WJEioWtYKkFZEMgiCwLeazeh2GLOtl/WAcSZNRov4G/1ccvcS8CE3/fLqQAIaslN4tN4OZ
1uQQpUMcxt2EL3B8UtsAZ4jGbLBxsSDW76GY1uoQemwqVPsSGqEwAsoYWgjJc4XIf6ovLyOGcoqb
d2Cbf0geRYl0LCjq5rk/6wTLMe/T/Hs9o71Po7+M50VieR3oTn3jMt0FyBoNQ8lh3MUiMDiSRXGA
xA1ZYFauJiaY/RUebro47s6joiOLoJnnJX2w5RI9TKFAtT+mNV7Q466UBB+mXhaB5HaVrgdSF/W5
H8MDyq7AjXykID7q/iasgV0jKXAnzJuTlVZYMnuDPzvyFIUq4zZaHvB/OrsyN7BjMdshlyKixRup
vAzXXq32tmH6vlxLgbGEul3x8GsQpQIrurpm3jFyDvMYcAYielDK6BteKFTw9rdk93D/O6YwyvCZ
JfaTUJAVphdg5NaSXm/MuQeMaF8IawAF4XLjNBpGTv+hZmtUeI0jww6v38yuojn3iK2lH9kJ+2GF
7iaiIXfcyu4oKpaq5xf1709bhHzBe6/52NEV7iqYeRxTlZTdmwQJRNt7gILbvbeaH3jI5r+Pdeea
mdLxKn+Liwz/N/8ehTrxFCUd4L4x1zWkgGZTCtYHLTMOs7DqTXdS8Vty7N9iodkw4BMccDjmS2CW
urQaeuY24xXjh4PMcZtqCy9nalinSfykYj3cnQOEN65X42FSz8sIS4p9guVBjt3VieS00XDqkJNf
M0+gpvP6nH80YRib7V2YCpb2GifCB3ggbuUO2VpVDR976nKIaw9UlnOcd+ZS95U3+IRUFJq4q4xF
ktbsWt4cpYjmfgBrxKkywrIwvOd8K3vlzIl//bi7U9qTqahHzhxstZKWeHYQIcM+ZzlLANZRo8fQ
delxHAqazcLpaamQ9oeHVvd0Gf7FRfEyXRPxTAdU86ZWTu8q1BLqTWjgr9HecjTOwC/dZYoumzFC
VwBtuINX6SaD1TgANv1Txz6Uc46xHPRj2Xw45FUGBBR815qt4ClvdcPxd1r4v9oal3M30kY9KiA5
Sqy83XxmNGQAbEA2JBlEWa9vLyDXh6bCQmD0IEGf+zycoXrbnBTi87wBTqX9viKUkOxJUR4Qim5m
+GkKD4SwpfgiCgdoeNqPqGVd5sTfVBmBjTqaX5kSCxT1qraqv4zEXRjot4b3pZFVQBEp/rHgyPSd
uPpSsZaT+fEUA7FXPpYE1SPcyu3xPk+bGun92PxGmusGk69xD0F8gr3/DrEIsAlEVrg1/PU7Zj4j
c0joA61GIluKZ2wgTwVGIIyZJ+GzKGE/xtoWi8ltnMHehkyyL4sHMww+DzvYhV+QsXXyqRGnE5FO
HdqsyQiZlFWPkM7IOrq+pMmlFmZfZLdW1cePgWJHZRvmQ1BAp1ctRS2/jdgjUflIGk9vBryFlOlY
lKEZW55m1cMN4U5WVhNSWVnIjBYNGFW7QxPaLGzkQUkiDS5OLQSASmNpiLkmY+VDo5TcNt8UfB8o
diJk5imLTy7XawwyCyqNpURMzPILxXbCnj57+4JGjC0Gb/7ReCaaWpHZQBwyP4oWDlppcbmEE5NQ
FMxfduAPsJ2NEpXe5AQ+IF8cmPIxsv7iBmRbS60yXoPW1u3IYiChE41Yf1wMXOM/ZbtA8DOkhNiN
GP3k1ipRvNhkGjmFxJ3KQ70YqzTQTF4hgNdfZCG65XxrB3Jee0CzpsISXUMNE8UF6oHGanGCEom0
23CXtLxJHT4xonp0f7DZlrT2x8hcBdIQvCW9EckZnWTgs0MCSpBg0w5056pQygnHip3BQmZsQ/8E
p0Pd1ve3jj9OCNapeT0zFNn9XRcihPe/5JppWDBR0BDIZ88FfCms7RGbxtfXVDp82JE6jKgdE9rC
efP6rNRV15Fm4cIadnYS9KAYzQfVtKlZjJ3zITJswn9i+hgr/j0Yc/lLJzv6cnN+FPE/WHJobZW8
gHmkK/NNbWdPNOslSolZJ6KrVY3J7vkHeiuGdBjl07MklWscISpntXrHiebz3w19ECv20uEv58y3
A8RC7aAaFtkiq9774dpbRCQ5usKujdONMAYFBenRm7r3Ekf9CesQviMAZdAavChrJtowyGA0UYYe
h486wULhoy/ghKc0tX7K5LsJjnWLwvADv3WCVNJPPWq5dzmtoG/ayN5vP8ihQ0BsaQD4bmRI3CjU
H6cjtBkqjFUsilbobdywsURaGUT8aQJ9o/Sg5Kg6nZZ2mBPN9HXVteRbfjVOiXnE7ywkoHdavXu/
KrrQfvb1XsZ9AOh5hBXGQhf/IRjpqpAds5Q4ZLNpYX2wQoqnjm0Rl+uIti8gbMRHuaNx/szeBQth
zOg0dXP8bkRSVcHsQX+jj7yPqa9zjrr0nSWTu3aCeq26HJ1bhsdYXBpe8kBqW0hewp0J9OXzFIwn
HE92sU76gLU+Q5M3SrfoXzBEUu7F61xOHE8JoloE2gKLpXxcctqRShw1n02q3V+TWebPKX82vTMy
8ltzfzCElvGzzS0AqBUxyKVkWkOC0a5ZUY6EqDJZnxCPvpZ572O3bx5o7+o9EivAA7wDQ8ThYLqY
aKv6Nrp3xps3gf2Rx3c/XPbW627GAejrCq4dytGAZDn9fewogmtvFgxhqV9BG7gfm/kk330PKuxe
jl9m/XiZJC0XTr2G6W4Nc4vC6tza31CPyUs6ZQ1+W/MpA9xSfHtebM7UlPADnlPXWhHGT/cEIpDQ
+I1m5DdKhFbxzPX8VY+N7A6OT+aQgf7p/9vKvVj1LudDzCpygKL9D5Y4D9/Syg/BMYECLWgg6VSE
Wdhbm1ia5EDdFXYbsiYaxwV/xB13WF09F93NOkeE1uuU2rF9OLLtZEC8xv1GP/RWcpoKT0ZGTOlH
l787BwTFXhCWSkEWGiYfHfGBMhBt3d/dVADffqRvkLQSqR82ee/LtCNuzxiLfiG9kJuwyBe0+sMJ
NhpaMwCSaird0SN+3lQJq4Sj86CQ858Hx5QpAMipUBT7UUUp5tg0zy/amnSU6zlnrf09Hhiv0ZsH
m6uqRFmEK3K8T1Bb9feTF+pJ0ePv3Fu2yV5JT4S0aVR48DthsgvgurmrgrfSGztsHUdxkcx/XnKi
DFDLSCewCsnIPSd5ieWzTo4oteBGQQ7KPDYa8wjWf9dixtjD+SA7xge67yUNXBFBm0V4t+Hw1DXg
19v8OSwdEiHFO5k1GYC24owEsj91gZcEyDarNd5fEdAoUMTBACgy6CRUzuQLdsRHD7Z/2SXHENVa
Wq/+PBjBQlDyOEO0zmr9t5vBCVxIFk57VoQ7D8TOnIv3gSP7aAZtzXb3wE+PfVFLIEgbwRUcMA4L
5rE4MgQ/EUpi3HciBkQCxm9Ifw+ZXzmr3home50Jtxm679TPFm+Li0QeWvSMaduEVNTSAqrjiMof
AUphJMBFH1K1wpi5i0vLkqM9V6R1izehKxccrlP7rBhyph6ZYnRC50QibABW5c2t3FceWJ6/5k0r
g6AoJb460f/Ij+YNCW8ssJopQWNr65c6Iesg9y2rzDhYDOq/JSmeHHjBrIiizAGMVNeLj+Uz7FWX
7ld388QdqHSmjA0OiJtw5f/OUnQpB3wgrmaOUSzkTnPjdK0kOMrwMtOM9BVajv8ZplfimlhmuS3D
/h8p7OBASNMQpw/TIRbe01/UTN0RJUnUjSQu/BPqds0HzrM1qlG8S3+XKBkrZ/HYSZxLbwpZgb+/
egrrpXEjUx+xkjorvYgUjj+V+Dv1ln6Pa4qAV5Y75bJ0GF29ABd/spbeyJiN7EXYqJ+Kk4ZYqUya
P3grjidgxkhMANuBVa71wrr2XkRpXlxI694MB8iFhyWo1lzKh3Qa0thNbpETUBCQn85SNrefnL31
R3YY6/X8S1SE0HxfxdMdU3HBjAZhSVFHHsC82DKu3vvN9x3VF0geq0WkM8ZF32ogHdrtO2fKYb3F
EPsiFqXycRoLNxm0CulOxh95AuBQVAvj5av+FmMNZIhgVtOULdMJIPy5DgMldLXWwbl59HtzqZuX
4afOnXyaii0RN126mS1TIXWe1cmuZS28PMVzO6evs0hKdf3gAspLtK+BHiH7YWIqGXd/ES5QZD0d
9N+J0yVyQkf5FM0VIwzO/cneMdfaTluk2EEZ7Gw2TbV3PU35nhHO1EDe2vXRQPBmxFgiSJTTHoht
okL2UYVycq7Q1Jm5ca1deoYpliSJlm6BcpPmtO/fnDwS6eoZeLQCuwDbN97AzGzEeBeeU+NqZFGV
+8pJ7kP6KmEdxJJHNapBz6hztrV+gAZtX67HeC7TDR99+izMVNBxI+6WyL5DQRdNyOYJwy6gcwKB
LwJWLtLI44LJkGVTNn1c4Oi1Oks8fiUzOUYKbkj9OyphNjumfPdgcnt1mAIzwVm7ANlearOt9Ua2
yVXr5tW0eBM9cJHDi7x+zp5Wg7m6w+Sei2jFAQm5CR3O97PKYFPLZjkE7i1lvadyuZXoRZCWDr06
2nwhDACQlBBkCCt11UqtxV8MHsf3x0TaSZOmNzTqmcwqHq1uqJLUveig+psTXyIJeNaj6kV6ExOw
7pCzc/r5V5YnX5wb17tyOtKCKb02gsCIMQxg9tE3Fh5FXZpNBqb6rDCTc87kOdG385Hcayinv6Yf
U2DGrn50YU8cEy11kBezpG4Cl3BL0euF3v/ZypLaHHOl1TCc7ogFu+nIAm4Z+dCWpwhfR1UorN6I
5YEIxzGLELWgbhdm0H4YpPx2EsBUO9EDb4vfvYYnrbLQSGrJkyN85xn/eL4ajF4e5eKl6fb8tEc3
FLv5mZFOQ0X+LQLtr13mU70vWFi8SrXRfTZB2Q3hNVwoVkGgN7tIH4GsfaeNOSfIMu3XUA3hQ8C9
w9ZoVWe+y5eBck8ZSmj7Ejq/28nyrqVtbEAalxvfNq9C/SI1ODPx9iEDi/ZMPu2lPjm502iTmL/5
zP85gn9kWn8355SBtdhPJABVgZe4ebO0C0tl2fQVR9FtqN+2EMQhjcIMv4VlYKDuQWMhuhGgrmru
alF3rcYXy3DAp3/c6FXq5/zBG+0Ad7n/gEO7CU0Q9PE7hXzD94Nro5iR+MxEp7+c1dWOR1pYYHpU
iB2HXpbUwMhKaZTEvhCStmfPf/vxw/lkm5MIhA+GUGhwWh84R+JBM4v7tK2Ej077MYNCTPNuM4nj
T0kibMX3u6sVQjilkaw8fdxNWRExteecEmBNe9/DJvLh8zIzaeYikN/BZFtxnC6YoPTGAclsMAZ1
YovG9Y6PDIwxSLH3cZ2p2JfEgbsWRJq0gJGz+OU195sBY6qA5sI0dFL5SMGRQm2lc9tWvtqhKI0F
eLOll9pfYGrPBD2ABcs11iAuShmIY6yz1mC2RBGRncHbv1h4za/DqkPbnQ/AtxL+6q4laj69S0xF
YPLwlB9ezc8B+959cgpceagW3TNt26dhpuYVr1YAZUFYk0C7O94K7FeRU8PRklNv8DLOzrYHUYfJ
/2oeeQInJICMCK4A+HdCWSIlXg4w0SBNGl7mlgbK7GSH5Z+O3cqMk8wT6/ntswnywg8oB+HP5C77
Gner5Ll76/p11NbDGekBbAjUeWsWMz7uthyhbS1e8PVlrdG8/ZrwkVSixd4ewdQd2UqC1tHwP/Az
Fwmfl4dq40IOD6LUJ1uaUf92eFa5xcFiadO/9UE161vaqffBsbHEMln67F8qct2YB4ePa2g+iCEW
TiJB8wktRERY6h8cZ6KMZhdg0FHZgUskJQQ26a9aoGutKB/eGlpD8MVSPjP4wMziTPNtKGNAa2vo
JjY09qMHfGnYaa0/pf17gRyBNapTBDcJKUjfVafRyk7LrCVRHs10QmESiBFlikV+OnhwqkrGEjNi
VkaBcDvJdxFYhqyDG7E+Yr8NRAxvqAd2/c3kEXHAnQEAjUFeAyjHRNoPaZBVksJqvddeg+L/gqhO
NUMZpjuBS4gavNg0/aDK9YJMPnaERTW0UJcB0006uCp1Rc0ZDHIacCZOT/lb7nBWjhi/Wu1wk4+3
i94pfqT9sAKlk+phEkOLFVpK7OZXLRWzxR6oQNu34z3b9IWTZnjqrWEefDNIchFavPQs/wK8k8ox
0pnkfijP3Uqff+bChzmbzzDjYF6uOqcr8oIU2kttdXuX5jm9jiqdZAk/c+8U2AHwL0s480E9va9Z
DylxEpxa9O+FUSB2JjS4uHoqBgE935cbA21GOcc8vZ85gT5gjpqnu83/AGAJorOUB4OhJe9BOKwB
fulBZY4Lu+9wJV9LshviF3V2oD7O7BjG0B79nqri5h3WZ/075zvLmsuoVMFowP25EccPbNNqAUEr
+IlxhUs2vDEGIRbTJab2SxPZVgtXNJUgEjNzSXMJYyfW8IQ3tmqt3nU4ZImhHtFJnj0C3052HAZG
JRaaBJkxgSMbclt1/ATm/jMnCCWeRculCu5Zt6yRJyjBMUlJMQGE5gFwjNVfLw8aynDYuqPW5kN1
G6EbRWXgqgIK4/0unh/uR0lZI/BKSBUpy/1Wc2zZMla19SNzct25nowZ4SJKd+9nazt4Q/4TrwV3
ECbDyCNprIlF8HMt97Ocrz0+2IPI4ljWfsJRZEbMOEpJ9Vz0ENJaOvyA4Xj/iXWxLmsNMC84w4TX
28VQA67RlgA77a65B9+aCiesYMxX9h5agZBk19ekvKOwkPk8wGZQ2/FBI8/YJyqIcS0BFkUvlKi4
uSBrFnEGBJ7DaCLJYd388d17MYxSg+ZUPrE9DJGrXzYXX+y9EX4zIoOmCP7/huaJ3JqqYzX4TGqs
hSaioTbY50sJaxztLEvoAi1ffgdFyb80MXkEFOx8xgzAx5Pz3OCfdLBYn5xkdaNBA2z52aqsP3F1
I+/cB8tFcgZwVyYc0LFrIMv0xDF9lpx3Lyr+KYYYrj3s379b/Zd1J2bCk83rPQpSBC4tNaEdt8i4
xspbEYgpHeT79NkcP1K4V8gMqlbmoBGiFZamz5EACdaiJicHAtYK9c3CTM1QhgwiHRk/MSXIwlS1
QGhDDaWPpMG2aerEHKtz4vf5/ItYyOtSbESWZb8SRWLXxDXhg0JWmLGOfvRs925x//08TYdV3scP
72rlTQqMpL1p5VcaqqZMFQF6hBrch/N3q6ozcJdTNKfE+3nlFA/EelZmI73TX3UIcd1xNTrxa7Ef
wukPldsTTNBOzL0350X89MsS6jf+cwukAXED1IDj+Io44h1g9Cst3d6kO0RyGgZE+2uiJ44AjBLv
7oWFU31xwVXVdIEBsQHmsKL1sF7sAHV80sLtxDTqS0ZNzMdtY7NXFZRXt/67VrmwOuXRNwva8pGH
SVhfwyHczlzPHoSpOhnHnRc2WPkLAylZTkYf5v5wa2kFC7jGQsaatZuJZU5mlFtp3h0X/0tPoObs
IEXrA/c2zcWeG6VCosQDyNz9yKH8bkVC0vf8qrxJPgaA6b0JFGT9VvAKai0wRNdUeNbTZa8Sn3VO
3gQgpmS6OUWLgQyJs+NejYZDaZVK/50InUJ/yAp1KUlodhQHFrWs+qbHLmMPw4rZcUHyXZVX1NuN
wPUoJzD+cD4IwWvCRw9CNfOwpEoAveQGw/rDvyke6XVF6JxZK/fy4tSvVc2TNPYrNfwrT6XR2z3t
yuKplAx6JV88juYU9PhJbDC6XxxhvLWYhb+hRnyU++1VTBnXqbicDp/7lIeYDiExe9njkYstlbnk
G/yryN1XjRkoULVgyzMTpRPe/vKcsBkXA1UqAr/n9n4/2uo6slZZyeCT8F+zuE64K1MFLe6xotdE
P5apiQ2hHy4D5g9JaMtBF/ujS++N7IqSHgyjc7043x5QcecCUvRB3xssq8WmxS8L4vr1gIGoC5Dz
xuiB7HXgD589CouOGh+AJvjLPWmi5A46a9J0HzkNUMpPgWXWQC/fXE80+2Bs+AZ8lAQl6CHA3D9V
F2hXBK8XgnZvgcfkodKaIU4sOF+ON+fzyY2E9+ZKxv63lcT2tjYT/tfME2Ypu6OjmphEdJ0zQ6PR
BaYzItfSwYaW/HQOc5g1RAccYKyxRYLMjYKcOW4HM6fwbPoDyTz8eHnR9OPuiSIBNtvarNuGy/Zh
m/I8Kq1ICXH9USBKjSiL05eOx6/iGQN0zosb8fTXdLiBJNIToeI9WGazr6UHp3wulb28T2yqxwRi
d99SB17GGSB0NIE1cThyKwNfcAgcdqTcvmIb/T0sFNARS8kH3nW7uilH9hgxmmt+B/3L8SKfRYjZ
2ACNzaD44Ab6dHcit+JN/WKzgTNmeFKje8CXmoccmXWBHlbFtSdX78Epe9TRR/2W/n+nVR8WQTSK
AXOWYK39RCYcrEwkJqbNOPI7CfywS/dxz/9nSSnF9q6DhP0N3qFpxLGhi4rfs7eqimYOJpeNYpt7
EX9R8cU2udzVJrm0czfJfpDbYw485xLQJUHtmdlM8vOdI3auJsBfK2NrrSuEjngaOFPLsZoHmsWQ
8FQTth5M7UCpJQR44L/8VCj0iOvK5q4DgjBBG3nofr4uL+dTdRHLrfWJsPVMmJ2r58XgbCmAYaMi
nG+XulPYqBcGDjVcA1LTlBsC4rHcM8vp7xu9DiGZnMgLUSRdxyxxEikTYk96WV3FXGicDo79v+yx
qLye25OQBCllq0M5rcHcrhgo5qQ+P5xIyCiheRhqyR9CBixHeekVQQtA9qjjYqgOxdgryAuOcHBu
Kp2SOQ/HjpmZGnqJ9i3XHo8b4Qopjf7v1GBLD2eLqBhr1DpcPG1eY4Pa8oaeNpNA8fUy1vyTFB3G
03BwDeU53I0Qnsgy1Ainl51VIVuf1GkJtJxg3XSzSUJKssmt8bV3cj535k2WjnJ34XC7jUxfBYgC
PB/0cVIeplOLS4qMtFZyCNYYxI5+tFxeb6p1y+N0RlU4lqqztoE7IJueGVrIm7WC6aJwrQ2Pp+Z2
uE9HOOxiYrvYdQwbO2wL93iL5ajmIALEfQZhb/aLyrQdQ70g+6UZPURroqaU1yo64kOGc3K3D8/n
bH4+cXkt6NMOnDigxonEt3PDrD+RodSD6CZDxR047Flve/5G4yo7dLhvW6Iw/IdWSvuhVduGgEKT
YUDBsh31YKJ7d/CJQKMyyPVC+t59d7v1f+pOn1xRggsNPAbID/CkcFi7mOO844gJEgLIEFfwrdCB
a+5KNmFfNBxUu7OMknVLg5GHJsNVe/CRfANjcFAu2niBftmPT4V7VnvrQ6H4uVnkDUhA98yBIQVZ
MGc99JE+vEkGZjgmBYl0Ps6wsRMm7AlYD8icmmQF21iprc8ZNCfPwCR0AJD9oJ/LQzLOU1RdtbJg
CfSBwkLbLsh9IP6xIVmYlGZr7tGmzTR6SDj0aW1HhQY+ymNuOFoDKhAIIT1NwqWkkdKn6W2CgPEv
VYT9kljB+m5Q09HIWRY/N5nEAPi+1Z7hLRpFCGf+wGx/ozYW23/Q1jqBQFrCGxTZ05Fv/dfCTNG2
JM/LCaysY30HzIUges7r4tzme+HY8gGpqIZ2E2egj4Y31kup2DBZbZh/u8u39B3xCKsimi2y3asM
Rpg1cvyCO3VsXXnZOIl4Dio1tCGccEjRWFvXIpfLq9OPYSqI4y/qdLCFQwh79aUjaXm1MbwsuFnS
fs/p8RrMKJaGxWhZDr7xWyOuVYGr4r7lt8SGVbfbPlEBSFy8a8TOTmJ9dTqsdHaIt74xAy5qrhxs
cwyaIV46tA0jFfY7rh29EKA6DCemalYgBst6eF3vlOkZtZHWOAqyaX4Hcu1a5gkP7SwplIrT6KQ4
xmxUecC1raVVXe1gsSpKrXUSn96zfZUNnAXsI6KJKgoHHkiZ/F9l7MrlaVnuFR3TkZCK6GqZGS+D
XRiGIbJ8uCrjh89PTCLYWV2dXCXeZA17zSky8S0zO+xaiKQaG2H/Sm2bk8oSXq7H9I/Z7SWsQzLZ
rs9ou4ju3O/y3p4wXNxvG2cYXIKlXDsg5ORiGMqn/ccxxbf4f2r/kr5JCXOYq/0ABg3ejWgajoRd
52732Bi5kw68pM8+ZkJrsEPgiLi9cx2NxpmWDaKBrLcY9wOLYNICTQg6KyjuejRtXB5XNiYhh0gS
l1wNSpAWFGIXuMsp+r4a1XCr0d8jmydBpGmy1nd4MiJSUlRjYM571mXPBFHnkcvgMbTqfOlhHwGl
L/q0JLStF2ctWRJOnSAsF9Z1POmotaszv1/AbZmnbiszMwKKUjIhzswfRaTpuuQy7e6FVyNmULnE
5V0kjiSiGmXTXZLmbbeHXqJT5eDd3XgJPgjQUTJ99pmftNWy7TOT5iGPd+ywmrgAa3g3ob4d9dyw
LYTCgrYHqmPMUrnGCvq2nwy9h0wa7p0NFjcut0AffdKh2YeKIecRixA8v+x4/KEw3FCHS1Gds9m5
/PORn3+FMxN5fBjZInTxVgjo9XMErmz8pkPXJ/7P+crw+JQqOx7A2aAJ+FcbqnbqhacATE/TTudb
rDLHFptt6tZKTTEoDf6zt7Ji7fOecoKqwktJC+oOaWzEI9gJWCP/mS2eQAJQ/gjVD9ItZZNEsnVv
MhDQv6xwIETRPh0RPTABUpG85xF1DF6q9DIHyWJCMfXCRPk6oo9OpFHeY/UA4Q+wrjGKxlhVJH3e
zqCpL4zR6fWwGJiZxMEuUb75rINhARpfqjaCsHZBPwoPVxexTsOsvmq8SL+IMNU+fLBjZz9nTwZG
Ygt8nzWABpoQxIrYDOT5hvC21JmZqBDI0bVpcwhxs/hmA0DsrLP9a2wZiNDqV5a3LFWRm5eRsooq
BmtxCOOM0+EXryPp3S3ZRBsqN+jxHafl98Yi/XAUN4fx3RTTraU/AwHj5QAKSITt76xD3uP5RfD/
zNAapSYH+2ZLStuZd76d6UrjF+k2meZDQPTm/376ubb0BI3FgILC70rFcr6GV+DRYOk6CcnNZUC3
GFsdbaqL4GQIlCyrbxiJ0b+00DQnNCYd2Ei7n/QghGC0SBEeQxdoOpNBGoKuFdcu6wW0s5hZhlJE
aXAOUXuY4NwTvQMBv4BR7JoxzF01V4jWX2XhDHszeHcvaQzGVm/2PWq2v9WoE1il/1mvkRUUmBt2
FiuxlpVKG1a8wBpBwFgLudAATJsFwe7e7mADZ0p+mdvapeuQHsJlwoUqOUSa4QReLLeREvoMm8Pu
TfFmkC401xY008GQTFc8BSu526hlavt6PhS0GEBVnvmry+C/Po/f1zlw8ZVLBeyr6x3F73dL1vLB
/zziexJUI8+WKbLh7LsNK0UFLBU9Dy66CM4WNLyk266711PMejSuMsdJ6vAc4DDFqgS3KIIvCE0w
32c0w86RqSraqCMtH4vE6xGxoC5p2QH4R15JvWLwaDnI58Bp1kqd7xwKFjFyeD6t7UmvnL6lcT2c
UwFSVFjMTez6VsxyXuLWC5o2j9fAJN7BgK05zctCcywsRw6HD2qL4qBlub1oBd2YeDv5LTeX8/L5
LX4aihMaCssinAkAkLXYTIs/OlCI4iqHPhPX44S+l0bDieWDs/POAk0ysa/Prz9owRQK1v0MvrE+
+FE/WA3XK1k1d7NNwl2J1dGR05+qvqbWeHU+RGugqq5mTBt+r8TznrK9VhiVMYgsFeoxUT87xC65
QadFWIY5BRM3bhjrv6kqTHUeI7mUClwPAc/iEqukPZIMQPmSN/MoSBa0NSYjRj2QQ1ZTc/e4KcIg
XScipgNCJAy1R912xtIVIr6yt0pObIRVLrZsC67KS+j9AplPSvYwaMfO6R6U7Vuej7HdbplnvJbh
Jy5HL0WwkH4X3Ig4xj0volgF1kTi7onqzeuRMC/1oAtJJmjj2Uo3c1wuRyE8Va70D75TsQE10zBa
uy08Lc+GSB1FvW8ZyoWveUAp2LQrD2/UZhNUE7LnqOthSS0pRDCLb6AbXQKBzhJSF4mgD6ab00sm
GNTYXrP4kofJk/PJRc3YXtqnu+a/RrRnoDItxiR9kU+0RP4ciJLGbEJFeGR1FtV25/0pCXc65L3l
riQlIcIC3hn8jwkraIW3L4LqT8fXX64ovsVSUpJ3aQ+3CSVJ/y5eV/xPblULZjioYCvxWLqy61GQ
/90fmW17XapJMalHz22RmWaw5vARykssoVts+dosnBzS4Z9kmYS4CXyQwcWzfhtig1kA6JLe/ifr
SPQqUvHGlKUhULLOzx42xSY9+ri/r4NTRtD5m+NcX3i38UAX/3nPID1+3jB34UcVQIZPtKltRN5X
hVACEu6WtpBIMmNkdDci9Su/rNJz9tI4qhbZie9OoE3xlmmti38HJ+lzO1MbYv88vA/AVvlyLCHM
v3vD8irWGDna66rryBvfY1cDLlMS8MQPeA2t+cSBgQcEBSbW97dXPp13d6Ev0SWI5I0DIwvW4dAv
gb97mkQOTzaknn/FWKWDK6OZWXaGc67QR4/+EgxxVJ4e10QRXSpD9RC6IykYOwVJ/kvHfisGxWuK
ohExzV1k/7/uXw2g75/l1SqrgRJ4SIYBy1hx03wBenLWuLmtp4XPI9p7wFouWo3PFHDMeWRNksor
FLChd/WeffDYia4ZqJcEdDMVE915eytkaxg5S3NACBrICAJmrVUQ60tslIG8klVoWdKEOmibX0Do
5RGzQg/F912mfZrGNosGEH7fG6bhch57EUCUTHp8rHJYEJpHlPpLGZ6P77ZqHRfmvvAV0UXBMnV7
WdaofKIAZyuT2Ho1I0sZBqPekyxLRi+qITyQGfXDlXM/0RHtNRFn5OONmcwZjwogsOPWyAwjek3m
CTz2EphvRbH5LFeGCtOpQHIYhFHbS3t16kEZpb3WaHmA1XipB3MDk3XDGUYzjr37AWh9GzGkQ6JX
zZQZv+GUJl3o+rZ/3kYLZgfmIjlAb4AauDQYFkkC/DUniS5p/NQq1lI5GasbYC/hEo2yQ9rJuHfG
4n9ULrrgGBbunnpLML9NC/KKlr4fcpjFcn13u4vlgK+jhNw0w+2D708/aKAHS/bEfF5A1bwQ2/Yo
H0wPl0gMkEZUWaEskWRZ9pOGN4OGwuDqfPGiGzc75aYcIWtcbYoww/zlXJWINX0aeHDIQNXSly/U
UF9Ge7aHoxUKam9lE1uNl+h6Km0nQAsXpgZ9px/mMeAlUwXEANem+qLGuAMTdBVgf9HyO/NI4vBp
1LBqwRssuKIPOhqZ/bl00bVDK/QyL89GE2wxOIpWA0ZxwBhk9VBTAtZapcwi0EaCtb6N02ezbb7r
ZKKaHb3Bhbp85/Kb9pZ1AD2xjtJNdINRuqR4glOuQ4njgqhzuySw6dRZPnuOIqC6uVngBB8UoBdE
XRvs4l3I2A6a+AiAkUNCk8UMnnocfDnz2MOqXN2mlr3A35WA4WVHtF0fvaakNvNC1sPWJI/8z7Mr
87f6d0bSCjvhZOLCjxdoOACBy9MblCEEmC7QIhRCr4ENHN7fWtHfCFmEPvQ9CivGtWU7nWzXAI0p
Kh51wz8gqxkswgVcHOuY68zU9IKEEWQcPIWniWZCvHKbnwES1s5s5Ie8bhkH3avdFQk/xDdzqnNj
rX/Zj1D3nFWyRey7Iczl5sL5VAao6uzFnvIMsc63K/WJjzNqeQpkCrTbzCzIotr1eHyshN+xvq9h
1hheuE6iekTe3ecNXkJryQesISXtvtVpMt4Ria7wpRy6hOtejpmIrjSIpvz0380Xkv6An3muRG12
wosgLvkaTlAb4WVBzX32ykb6+zyZcKuuZCZglBtg/A6lkpFd2WfPafflNitfZtRliwthA99TaLTW
8IjO80q5qg/YK6hGTEPgN9jIgdBTemqyCRbPZp2V5gsJmVVXDKRjfuzitBCv4WwgPrllt6Opooxm
RKBp6L+piafvV9vx1OmS5iT5cGHrrIhf7ufbCgS+5r36s6g6CDNQeB8eUkV9G6e6kd3pFECl7K11
YMs9qPczdFTjfO/jNSLOweMnQuyA/SCwpsXVmxzD8tGojIDxYKaVc9F0ZvDqay7SVEzj1XrlL3zP
5oACPH2OxPYT/+klyKxu6spQEZGchWiUdpA0/Rsdvee7MjGEAfCtMICtL/6E2qcwHEhrfBCUo6sB
5KuAsBh39It4dHHBrem0cJL6McQP8FUJN7tt3pMkoDLylgPlR4ESLmq6rVFuKLTnY6X3I0Wnkgb3
imMAHgJanwfMHPZW+12cX3464+d1iM8Ihq1Y8nylI83r4bbT4jcu87IRJhv0nS3BpqIryHA43EgO
L2ZEDlsiyv3zkMx+9ANNNQfD8ERYySmm0xZc4s9okFN3r3dGgigjjys1Dvsp4r7HzWYmXJOaH0sc
FK/2nLxxB+97GzMndTbWIyXBzPfXgcH/tMc9BwNv7gGbHR0GVdfM2tH6r8H5rOEmJJ0r27ugaKjG
j/JcLq8J3s7DRes+A4ygj1KA3bXTWSdO+142HocUJED+pyz/zJgaPxRSGvW1otpb1XrM6blRzJip
jzsloMsJl0ZNDsZhIpJuJ1Xil7x+0uTz+jqDSKbsAL6CX6L2azd/9OOgBwiHtWneTWse4+8cUQea
Rx7AHkHZtzSVweYKvwFXaxq0DkeEEQNTFfP0ez28HcSIB8tF1n9qHEM/h3+xdXjxBegz4yPOQkpJ
hagGSXp6GwDmkgpFxh9z6ofwxKAfLnqw8HpfoURbRFMKxsC0mOEMsbvXtUYVGhnBz6G2waOgXyag
gO6neAu32S3S1+tnKYbqZeRQPm03+iRA/VhHSJ0jCx8Q0M/w+/OBN3t1q5Uu9hN3mwa5C6qduP3d
sMNIu/jCHSBauR0NlTcHCKqf/YiPcVvWEa2Ck6mqKsgDgG8P65CSy+/d1m7lnWVV/BEkzsnL99Nh
rCHUkmhZs3M3zMZUtzlb+s1CfCYyynIkhy0pswIuU+O9n71ah3hbCAZkunyJAUNY+KxnlXoLLVWD
wUYaGTmlgsIGgaLehaV6gvUUa5BpFb16UH5JK+IxOrbD4jygS/Ibvmv6kDMvK0LQYfTExZW3TY/e
AdbZR7j97KUmlxrooCyglnyOyQWyMZrzu5uIBL2QQVpuBkRcdCvdG6SOkqKspw2NXmKjr1kdxykN
CDI6TScjsbDCRaE/Ppo8teXwEov84M5ReaAQAFoYGQ3XsbaDH5alkAtMi5ESPEaVw8AahSL+2j/C
mvGs9Xxb9hZUbXNC9Ei0P+5rSpjpruzdEyTw6LKRvW4yYGWd4WVIqF1Iwi7FQbv2TOIxylLa6ZF/
Da0metabd166zwbe5oXGFcdRSkvwYWILyQNWj/Wx1r8hkJiQSWmwN2sATb7koF3fH2Z7BQJ9lufi
CZbWYk/R5OaDBcThF+wgTIK72RTivHTeyN7SIcBEKAYoRvYtaA9dlrbiF/w4tYf0nzi9IH6+mPR+
tcQ5w6mEzKP62EZkgInBJ9wFLT3IegxhrwYh0avsQhwYrfxdvn6F9xqtFfLhTqnbZPGKbR822In6
frfldu6O39Z4/Gx1wI11/z6NxrOhqT5Jx/gC0yz6h/9exOWHez60hZdLLFKSCTgrfLIkAcR8JadZ
67SbccEfguZJyG/DHMt8iv3Ngjm8NDlsu7M1sED5cSfal0VZ19iTT4V3HvevbH9FMW+8YgY0n4XH
pWShBjVR65aTLP+pzWoyIG8UQr/n1AaHS8ofcd64FELvnOkNvVmhEaN1uD/jykEGx2JRiOHDD8Ap
rhds3QleydDgOf7Qdn4YByGEp3zIsNnbh8xT+ICwHMVwOC7GmfJpgu83tWFeAhXuH1utkj6dne2B
zkQIpVCOd1cOS6FTc8uUmZciNO87X3Mo+xIzmV2pe+yKTzmRqJHAgBZNxqdY0vpTlZ4MkInSweWV
TPNxsxvVGGRUFa6hjdgmK/BsaF43nXEtbZAS+xOl55aQ121Ok4b1j/FETrrG/UOxVXlRii6AIr6X
+n3l+vwb1ChmjdjHyi3oLGOGGTlMVYZLnPzTGl/ry5Ozi8tS+jdOiLRFWOJ1WjAHHBr8hZEqljwK
dmh3PAdjwEV6Nce55Ap3X4uxsPWDSFe/GUN2dDcnngN1BXO8n8MnakV5tAhVTGYcTxRPAtCF+2RS
kC541Uu4v6kQG9z8KnIb4Fgn0xrtGHPxKbO1UKPk5WcbIqw7qEitmdAc6hye/gvLsGt0U0zvpMM3
VD4K1imulfzE3/ZaficIUc+/6HeeQvRD/sYN07ACbih82h1JOt2Gh+F2KKHXVs42gScp69yNmZCu
sq3OKCGZE7PxBBcXxT676cEyEf1hIErEohN/EVqLDM00ikKNctOGV95K6Sy9ArL7JIuaeqCLIhg/
mxPhJTSIZkUSjnkp/CPQr3xdlDf0F+cPuvz5yC8cr9iU51rxGY6+vk9HIvKlIrrK9tftgXU4dDMe
+ZKCNR6J/dnq96ESaVxsll7Jh5SkJxEjELOmUwn5069dBnt1t+KahvfOZlDRL2MaDcDL+RA6KtJ6
v9/vdI2gb2bhgQ/NdEsMXwXS5u03qh4B0rbgaSy3kT5BNpZzfJtJHUMzfyLqduHvsaBWFEcS0EWk
yfYU9uQA0mRVZUWOPVjnjT9QvtBiB+4jb1790mBlSu6DhZY9PoScc1Pwpeqt8sUBh4cVsykSJc+2
dRmjMP/yckafT/RAXjmQKnRXb20ZXR9HtqSWYeyBnnhefDeYfhLdntN9FNcXn4aD4T89QOiGs276
NKuPPUnQHkmZ538BKCO8kURhGfxERSQv8mEgOObCfDZCC6eak7dZx5Ff+eR7K0EVtP6MEFA3gl5K
IZb0ETETME1R4+PZwbvMcK8IBMnJIs6Az/r/tHFFC/UpBhRcSuiWr9ofjjsCDHYtOCVDWI4aCMLb
FC5ZLoq4bq7fYST/pfd4QiYUZ8hNomE5NtNxChXu8qnBy5McbtNu2egHy24Y4h6xqM/kepmk/i09
gAkPpkjbQOMnNvX1MNNfyGIWm8i5Djyob0JPAp4WTb290+Xe+PqQozyfTdwwUONW6wG2x8bbTGvj
nLO/X+EIuSBnvn7K4asIdtSTiC5gk4Yp+a6w3mPSEntDyWr4M5xbolIwEcLK7iZlTVkYpAqnDD1n
Nww4CCa7v2ZWiTELFqIN3cYIiumQnwsvLjLL1dVRWhQFVuubxTjyhmtrmOSxmlt0c73PNW6bqCjb
UP6zIPPweqytGd44pHHOjVRUCyAGrrRwH3tYIMEshcMt1TtuhybNkjydf9KpOH4f0vHuJz8pctJb
AxWgIPjSqAylKA9Bcts42L7XftZvB3BzX2K726w/uqdlsyfZOdq9PtQMqLejf3FC3WBBHkKnn3KR
JDdC3UAKT7dFGqooAKKhTCEL9JBHNRhSnsBxfeV0XhK3TcWWe9jEnjxnkSF59F5hn4S1QJPAT7sS
hJCVj6Lp5zRyyKKnRrmcf9LM1OJNaVbrwYFnZYaxSK+Ym1h7o26Cmsemg/LfUH3C8IiWxGbwiDmN
XnudiQTWV4DcnKttxzEdIRWlaV8jop8YuR5Be5BUFNKvPptuYukn+kVAtW5sBOMadUp0MLmfLmTp
8rH25vkZkk4at8Pactiv2XtVJhjHoGHulFe8UIL3F55WUgX14UUx2d6KQGQ6LlU3NLiFCbYhZi5h
AQ9fo7P6qEU+ckMlr4NalH2WqTVVZ7D2lDaSoTDC5wAethPUVBGQxVgITOWfWNxNG5YrJXpSJrmI
TZWePkmz5POVQr09wGjlUtCAaGpUfhC3u/zFaakJ82uIxxDOdjpgEA9KgAP03oRmnL7SbRAVX7T2
l8vslAk+PmfzF4xsxMIlOBz1rFap4E735AX+e98QJlMgChbrNlNp4fHhBonQwrC4VAc2g3h62UuZ
bbTT+H6836McJk/s1KScJtR1+4AjzXz4ErP3QkNThmPDUo7YCgl61qkcv2grQZsClr+TNVfn+7xJ
JUw9sanjJnGiUQIiJy/As4Y/30mCTXQrWhjf5MfnSMvpdq/ALLmDnw2GZylPkvaMejk9YHzoKq0p
4kpN0n2vrDofHnOovcfgsQtSyB5fpzu6nqmBjX9JBgYNmbOEs9l1dBovaFH2IYcZRFbIC3PvMlHJ
LvGouhHfFfhQBd3Qbr0Y+lvHXCsgOJE6e0yBiN3mtAWTqyO0wga2XEoWBLLByIQnDLdGI5LqwroQ
VRLLbLZ3hHGKg9XwYcEV8snY93BHIOAXbtsHjmnDWinAXnh97XecSgZcrJmIcAXXng190NSIck3y
K74010hxQA6tsvCH0FmgB+8iuH+No3K8gvt0orSOcsLZZpN0V0Ipuhysm+bZ0OolaR7Cfx5/Silh
v5MCzLFfQX7Rp9x2jP7lSC3dk0bJoMTxCniOjaUOV+8NxeptAQSdxGy2VmDt9+nK7wWvtypevjoM
PNv7X5GUAelDNiF2UYAU5f5q93OSIwtlRGKa0lDZ48tHan1Btr91gq2y2Xzk2JO8mQk/okVn6Bei
v+ISMDK0T+TvkbB0pm6g/gg+IJri8NAo75bwFRQTE0vJ5ChBJQULYITsPfDUDKguo3yUxJbMsog0
tRJSLqxqDNGWKHZjDDMirxVShCfgZGHI+7kiLeWn2eJiu7GfqcU8DuL+NxwjGsvuiqfD6MJxO1WA
1uzKP697QGs/gwhUyIlPKN/xXBp8nf79ypnQN+eSCa0dOsFaWFEjKr7sBkEaytWz9o0kQSkutSoC
JSuLdWgHxcGzoXUhCbndkVLB3T9auKDvEIRpvoI9HX/iHPCGVvLOZ5V7IjK189JxCkkl6Htr55p8
89h0hc/OJfJ92Lcln7YpUA3q/qxPmRSc8Fd7x4H2hh/lz/+sQ8ublMbwlM50QN9+0qc8tQ2DpYI0
e79YcCW0+LJJj4EkPqG4C2ZDrvaMI9qhB1Erdw4NFJiNNu2YjH9hnd4caiVCy7BwE0nhRa2CrfOF
1zkge4cEbgeNO+GTtDMWIfWNiI0W0b/Xgm5/gk8zYIMztWDrl9TAussSUnvcAerMWkUkALXu9SXe
PB28gU84P9px9kAwWcWUEH8FyGZE7Pi+WLWkIHaE1x0qUrvlaQgXgCRdK7X1floflCr5AysRhP1a
2eO/YOvI9ZYfS8JRKe/jZd5BSgYxlyKPNG2dRTW0jxZzzU5jnDtrD2j7dD/7ioQxonf+po38KbvF
7lyPK7EaLUDcuoW1UCh9iTJmAuksD9MlfSb3TwKRiApgDHeQvKVzHLJz6AcFgXUXxISE6e00Gbns
a/y7RGzXstGd8+vitrnGeEmB9SdDv7hCZuP+WQ5Qp8C9vxtCgIPD1f94r9kiGZAEzmWxnytJ00dp
j22t1zngyf1ihv+kYOlmWy/yoJyHwaEMmtyE6mmDMhakpeBSy0YZ7PSzcvlloPOpNGp7ZeEDsQr4
6EzMIeK6TzQLIJ1RK0YGrkiPYUd+Hdt/9kM8s4Wp6yfM0l/fqElrRkcFFvDxJ9mDawMCScZYxPyI
Jy+Qy6Dj8nke+kjL+zvagxRGWHHv+KNW/O6+4ExJaIKSC3c00dqtKncDaaTL5MdTWuMI5H7JQX6w
ZbO7UFNz/Mk4mIlDZDhMC2PNCNOyGWd7mn35eZaNQKc5WgretZNnLMKybSW69s5hGAXXKYMkFe4L
H0sXkHcwdpF8tO73Dod42OG6nFLEhMY1SgnJMnmq4JBaAgbhcLc1icqGAe0YaZOQ1DFPkSgoBW+T
uJSC7ocj2AKCOFnw1NzIm/glBCUC4tfc+eAQGoRTXrzr3YlIWrkJatjLrnemNTnQae/5JYdgzqN6
6wOtw7ic5uQwxBfkDtcSElXT3uU6La+7aAlhXmy1NPwAnonuQqgUSW3AsRRH69wa6krsWni3I8oG
7vUX9Ru6ABIWkpYTGLuC8Fdrk88kQN30CqMZ7cB+q2zkebbEh0fmvXizcFDhb/ppbf/mn7YhtsLs
4DlAZskNuvsjTS1YwN5AFp0l6XGn7lQAMQiGhitsj7+k99rmKkDsZ+XVToPBfjOBbN8WbX10Moj9
xrq6zjlJzBQBukG4rL5ZLuiHto2ZFg4vGEg9ZsqBV8+i4Cqqms3Dz1iCh8RIZ5RwleXdKQemp0+n
MzG1jc61lapA8q/rbZEfBL/s7QKShwZam11PunKFDD6+cR+kSb60c6RlRBS0wDzNNmElborCA3xj
Ucgz/bPnPhDMpPM5PwoSBoD8ZUEWexnQjxXKtVuWHLLu1oXrOjA0gA/v2dZaDthwd2TdgkD1SYnB
aGWXc8pEhFCqMt8CkI+TUuMnqk6jCDWCWuf7+4nUTvNyYgFUobJgjPO6dtepMwfoM/DAcDpUEIpG
bUJsc4mw9baYGqDkH+Cfa5yEDi3R08LdHyTDPaKM+Im/y/hjESVmdbDRoeB3fLb2mctGMXY6XbmB
HIsXrzXJ9oHIh2I37zyCPG/DnFUTuvxzwS8SyUbua9UJGCoYvBFkd0Yq0FOKvwMoPVX60wW6pV57
TYiEFI6J5xSnUzZMk75AhvxTbQYv4ysdmy5SrfJaIEoCI+sp9VziPdOr3/rC2//sNMgDJBbf2kuH
GOzguDmguKJjLUlCW8/NnHzGPZ0COkX1+ijObjhsdLJhrdWzEHm//ELmgufx/poxqY7GN7RcnnED
gWPGe7MFSOA6wjve+uRaernLe2tqyrnfFbcj+285mgj6PCGUe71DoYGIBUmPCNnuWcO9O1RvfVVw
Gkkx+RJ+C9llymGDFEBsUQSs5LikO0mPzHiNMJ/elbWY94zGhso3SRNNMY6MpJaTHLemh1Z4ptoe
RixbkR2jHIkJ6wvjDCLtW4YehpSSD2Bqoebig8K4h26kXFhk6+XTemH0Gd2DAkv6+Wz76xnmL0RH
HNvRh+5RUqESKeaeMvH1McPW29AKP5cYfTIcStBcMzWRCimdDJ+rYT+bU7D7QsYxfSlfHvSUUYyY
IrG5wniLM2Ek7x4yACG01aEQPlAYJYrI/5a3foINNVcIntu0po2k7ZhYxwFKPkxaXipm1ho7ez/N
b0fdHPJIVzFtFb4dEQ/y8ks/emiYU7kypziTGsnMY80UknlfbB5IMWbhvw+4EmLGAAmtqWu5lzkn
g5f30Huf3+GH28//EKkZ3G7jJiPni8DggtN1tgDuAZQA57Wmsl6WPz8UAS+P8LzVBCzVAscQl8F1
2LKbFfr3JkjJrShlra2NQ8MCQKWKgyK9d07/o0kYqb2M+KyNQNsYruEcskfF8uCO/m2lW6rds1WC
NKNxg0VPt30fgtBddjCwC+L3JdQ0nR7G53aqwVnXNj2lgq1xHSuRSX9hyryAWZFeC0Z1kTeMypqF
pXBl4M/8gMAstdsJkO/qU4KmtDuj9YEpx8JjOchA0lC/bhD/v74j2CDoHvUSMbBqZiX/3Fng+hjx
zLS9MFtMDoNn2TZnDNAL1NdTmJNZj0toD8jp6BHvvaTijGNkQ9qC0f6TvjlQtBkc3dSOiBpjggN9
MIDnKZQ3s0savohxqM+icd8/b7MmIhU6inubkOe4f2zlLuXZq7apUYpRQdZ9zyx3YJJ7/9Pka+eu
EDokNB3y5clC29jdEsqNaR8XTulElW/prm6N4o68JFRhJsY54QjFRhupYO461RxCzNX50IT+AHzs
16TbfdNdp0U8yTF38q8+ymEeOwSd3HO5Uyi3i2N9Tdl+NUlN02cW8gPGha4M045M8r3TqclNA+2w
QrkfvXhby6qaM7NU/ekunaDiPp4Q08z2DCzp/vX1NhKP7nMxx3CXPJdtLf9QMXvVBECTPke2Ovbz
DwrteN6k41gle3TgY1A90myF8UeBrwpEJcTubjcCd9jCCPACU/ld4dKR8a6uA1tvBem1Qyg6ED+m
rvj2nwaWXxosWEshT28GFB9GaZFB43ZebdRxuxK8RzGin/q2v/CyXhaCKj00zhVbqi4aeOrxUKi6
M/x91PYaoWBNd9DBaHwvPnv7tusUL7h4xYF+qmBqsW7kfM518Ip9wIOEpqoxpjyQaEk+L4g8Q7YM
3QkBwfofrem70i5CFtdpdIp0nnEQLjKnsRXc4lyr4qWenny7EMdsRvcnTOtjmesYC558zWDPRMke
2RBWapp4OejSP5qNxsMQtH1+fzy2xuhzvyyeXfl0feS6shg4pFoXKGurZysCd7faBTxa1fuoc7ry
3n4kMKXDNSQ33MYHgoTT2FSwGzVEsRxtLb5Dcs8zk33OltsVDBSuwc/m38pjPUl1NEQenVAoNd8v
YKcjFKM1YdyAeUOVwxgCx73IpY7Hp1i2yanFyPU50pIMKTn+M2r8IAT1hf9mbHDDH2MKhoOvT8E3
Ay9AvXX+I7Xfu+WRekCkE2Ukavf4co+FXMo9aWXdNzXZD0lcLappDb5BhEzUxBaR9/qYE/PyM+A6
Jvqv9ozS+B0NYd+8Vem6v2c6y3O/eOFjAUPc1swEbQ774TEENzACYny/zEm0ZcOKQlc6m9JpEhUB
vSO1LRtJqitSnfxlVq1j6ShZdAfOyoK0BNMqH/Lxk161tG4MzNMP+dSjniuwjzRRrzroLjoy7aqQ
4ytMtj51BkH3BpZQZTuwz8XyeYKBK/hdWHi4r/I6eiK8t4LwDBW+F+XwCEC/batfEXnKtV1t+BXG
Wfa7DQr78b130o83TXgxnLfBPAZSASaWTf7/BVLnbZj0ERx+C3F8w+QpS1gKmb5ykK/R4iSWou9B
y0Qjyoc/F6ksFZLmVvlIlcv1UwBIXXbBAEqwb1ES/09g2JhOlymsdHB5OoWuvVw0/pu/1QHcc+QY
VZcmZrMqppR6+a2Lsxf2tcheRSWNHp0HwQTQt/fmLRu+thHgC4iSYWszoJIK0rkyo0W+NKxZVQEa
DCHqeVOi98Jj/4lgsUNebdi+VT2gI3WzEIYlxib1s3RA9HqeWqXeR/7N4PLs0fSXo+GOTB2E7nme
eFmKQNYwSb3x7Dx/6BaHXcCZPymIRZFxZ9Q5IQI1+7ccAsPLw3Z+zu7B427QBlKDGYnVNsHpxqiS
yWAhkFkVFDV9h2DsNrSiiqZeoY7zNHMVlGB/wsjpYo0QvLw7/sR4Yr7Nz45+X1sBZCTDBH4E5WH2
SYiOpbpo4zrLhRstvp0iqxB59qh0YvCvnSdMWrQCf7lIkoqT8bLIoT/uyt9ncUy9JEYURcAa06qF
4PaNY43EssCbNHt68a+9pNUs/isRUKHEKLO8tEQePr3skWBnNDjwdx8XiCKT3tnMTd+c3LD1O9xL
eb4Zj9vwj4jzWQ9xZjhZ01y+DrkbEF89qRqYVFQSb8K4uZ9ngk5IDMb2dtpKOXC+KKcICUQgOM26
0cunPq9jlEl147Bt5+7JrIjUOyPTpPHOY6m4HjVIc6E/nlwOMYDAdO7dHnWkkgtzrW9jxsnwMgNL
iiyKvqQv93ondEuEP9rmyszvZFS81ukRfPCub9BULRX9ceuEogJzo51cC0JpakZN/q7G1IRZIF3b
UBH3jEA4dq8MKYejVp/1w8Ni8FpGvIrI/en41/u6Mtl8prd5YwcY3UlKkoES2eAjWAx3yOGKNboY
YaZ1dAbKrDW3+YA6RlKaVl6+Qzi74BiMQ5Pe1/gyB03gUp1xaEUZcjj0Q94AqysOOSe/vvCtd3ns
Sgogs+U+HvQQ4aNtjYfKwoT6A5dHwh42cff/Vv/KJo+c+HWqrYHYV9niL8ZCXWU8GN0VTdyD/Egt
lnQ9SH7UtrvBarzY0Qje346DUOpwwhefytCRw4thfXNgo5W6IEzUdPwnzSNazhKsagdW8q9FMnA9
2CfnH2cImlTKbC3CIwL0cKbxYo8hvqoRX4boFICQE6o2ids6YV9STvUzbJHyohXA/VBes665HtA3
1zNLZ4GbFGcsrTwJh5h6ILL4+Nq6T3RdTRaypxwxzT7iw/92BE7/V7eL4NKCrdC52xybs2k5LJ3b
FzjQjGmWLMmCPCHuNUTkOnuel792CzMLkVh6fsNaKVKmJxZdQohVmzKLpxXQHF8+n58/THvI8ATk
nZq57i9ZnEWF/eUQTgH4k02c9H5NCJ96jIBUjm0piZ0ZvsqWSia48kaNBqIashl55+01lBhPiBKT
ZU/0jp7Cv1Seca86sxTZUvjutuCjLj0eYUoLGzjtahf2xKIGTcuZvSnFPvT+Y0y39gsl1kvdqAu9
FzMlWpCt8Qg/hcUqtRn2WaIzWjwrXKPdBkt+ncbcH7jFmjN3lRz+XgRn2SuGZ1BNaOS4Wc7fbQts
D3QowgBgCBx81A7otvPqpn7SgknsMUELehKISNqqPWiM9h0vMg9bVPFGUPMVs/OrhwSQuZpJvm8G
byb6RBqUTTpZz8sDBHXWgwYqFgx+auToYI5IdNLvtzEefE+a5B+kipTQyhL7DOuvzXlU6/6MhRKm
PxGjXqtAdXMRWt78yL2/5aPNnLEZYDg/xkV89Ge2WR4bmYoPcVisJkMSoj28nkjnL8LVSMSl16Y9
E0HeFZ7Y41LQD8+dK7gzKV2K8bhp/nX2RkjO9uK1Te3nzJnZ0z7WW1rNEqKUqopnY4Y6VgEQbcvE
0BoUEdcFFdki8rufdgbJ9N/Zh0x2Sa15gUxMW0ilIuTaRy8f4Wuaw3AubfhW0GpSSVHqZTXoha+V
bhRmI1v/L1kRPnEiIVhn0FHxjuJa4Pbc871CEVLKPwumkgHI7V2o6njyYJpiKvBb4KJaEHP7k8wv
7jJEdtwQUbo1gxyEgGk4T0Xc6bvB+iMA3rvSTkmkRu6i30IEAuS7wLff0zM004zHmvh1gkPGs0/5
hB5LVxyOtzLpjVUpAOMj1aCJVf0Nxxcv0kEFr4Jsl01DU9NIpYBHCnBht4LQ4NK+FW6mE5UalVwX
+A6IoaTmMQdYxblkzFJrt7ZarFaansm968Wqg2xKiRjE1dCbncFJ29LzkBvI0vq/vD9dIeQVcLxi
G3pv5vrMIZR4+6Um5lSAePolMCwPqYqdMHlcjqH8xa6CT2Al/0Q9WzFdfkODsZtDIt4k/9rxPJqC
g6iyvUQFaa0lG7T5fEdTgKhDBARmm7az08Pu7dDmpoqnYc2WE6vCHmnoTuaCvVphZQjKnV3amRxR
5wLvMSQnsecDU3uKh+oeg7UZv2ENboyh/mjTuaUF1HiBTb9Qq75EziE+tneKBzo9ju44CJIHCb2E
swa0jA2jtayW0Bf/P8hvj7QUVSo7zkqDkbK4ZItWpuqNBVZvPea1D0OiU0Hf4Wau2Mc21P6jW2ud
UgJ8NqkLXEJDuQPtf1TFymF4tx7CC81Lj2DijYsOnnNJt32UXnkCGy2NYpSSd85U3qjo6A369P7z
9vYZmgBlWCouQTPiZsQqaShd8KVdGhBHblS3Q7IGSM467/a7IRM4kQkR2S4HHHn3ae+eXUMk+sMJ
XYzpSyfWYCQNHVTMzj8hApNVoc6v2RnMFRh1HjrW/lWEVhUyH9KwmRAJGPfWrdlSTzmmro6gKkFh
UGMQWCBxfJmWGTv29fvAOMEFh7o9I1/Xaco1AxwUj7QVHJj/y2yzv07fFsgHlUCw0RWI034EhFqw
MCq+kzephE2YhRFYlXegb9U/4Py7EwEQxL7dIkGIvbCBSrxlUvejtik0tGJg6/vMZgnwPIIty1JH
u3FFkHlPH+mqSsAQe+Xxv15sFOm4BtFNv1H7naWZB7HjPGMuRvWN1Fbm4tHpicR1D3mIQJhOFpFn
QfqEH6wrJEHA5gNTp01b0Z1cNNKW4nmvArOlV9QHdUPxuRh6qHVzXHYT1oVdQWz4qiGlT5U1+cPR
0L7ZMYiXQxzF+Il2O2xhlZTF04gkobT0zq6g89bt2e/7O/LDGNXw90fVPs+ob1HHF18mm/jM1Pt2
lm3yFKVyRpoNf+NJYbwIpnjL/78chxHc1jLWDg0z2Q4+OoGja+pmUfW9A3AWre5cY7w27unL2R52
BLNEMTkh1j7pJ79h1npNhM1qn3a1DGyD3uxnR9P+s//BA0wcH0//hHR5wyh6AEmhRSWPV40Hk4LE
UsNaHLbaKx7NHdD8/RemDjiMFIWebQRvd10aSm7+F93igmgvYYwj26vOsgTubf4BxcXKoTkzAqXM
Ep//3+nbhvH5K928tGueQlAN29ejCBzw28NKVxjquHT/4GLRxOasPDAZ/aR8zO51euvieHECtfEm
DQOQy8f/XA31gtgvYousNrDaaxmx7x17SA93kDv1XVjxsj4xN1wApP/mEZEJ70e5sMNub1UiPgNb
BBWoxDMh6q3oLCEX+CyWkhXK8Jr+YLWGyXNnPugUafCOtvwm7qiPWxbSkO9CwobbVN1MPOGFgaN0
Rk0VZ9JbDObWrMixOrs+z3RVrbp87EOYS8WdJTvRrVkhPPGSdDSbW9Rp4CITeqsyrjS3DKN9f8hw
MapZ/EhUMbuBYQH2MWI+NLQhbh5jbtIozoDLVs5vVS6JdWivY72nZma6dl7EWNs6qG2k4N9ACNvn
CA1C3xo/SNNOu5keNgC1EfMFwyWIlGSzS9A6NcoEECWuunpOxvYJgQwPcfQ0vRXz5nXBwPFEzYHV
ZuGeEcj4NFBkshIc/5y3SMfyWDPmGYe7bV8RPr1xETCKR9n8nrBmTG3d+GUHwW5S7MZ+4STAnTGS
pCMnfxgrXaw/BthRzJnGpMZ24asd5LK8zJM3TNidKQQLPgfcSH4/IGdoLnVse1Kqi243m/fdMSeT
1Wd1amOpj1FJ+WQ9vgPSgOkTjUChHEmxoR3z74BF76ibZgtw+0FspNBF44bxSpnXoggXph/ul74H
rNyyvoXsuaXyPeGEH70vSFgc7Q7gxkm4/kcrVW3blwJ+v5uAdMt8ux3w90vn1fLa0+y6qdd2yegE
pNG1EHuuZrdqJ2fGU4EhUoBWEsRy3jsPHvdakES6IHuHEFIokzOePrQ/vw+NLShHtwKiui+1EddL
XXw1QTCP/g71M6YUWHtcSNnK/sLTkdxkMY3csXvwOt66QCliZtYSl5GyuQAjS8yKUvWAeBwxBhSh
ttPAdAuHjzp+T6Xtsz74BvpgKFgXEQUXVi5/zczMNJXpNSEVIRozlMr+jUGdoh4idYif2KTM4CKm
no4EEZJ+dInj/t7TpEcVBAA/iB3g5ajX4Irvy/PCd0MqotVXLCvUajZtSnVK/vIGPKklVsjz3eJL
B0OLdEUrhkW4JwnoAcMnhaXbcqGJnlICIygGrMmHWo/sMC0bUkptR+/uPWFhvezs2zesVGLHUbyg
Xgy/34a4bNZdC2lTI6YSOL7V10YFshpHh5EkzPFT/DF7uY5pAnhdOaxrcwFYv44AARKA+3O1xdaM
F+AudY3Xp2tbx1Y6jSdzCjxPKfy7BbimKLK0qc3/Sl/0ncoBQnzqamUvzDFmgZgXbQmB/7st6H9P
BSwVry1XQaiGjVvBoNktVJ/hw5SvQ3EkKPZbA1Sy/R5ZdROolW22fNz4TxnoNZ3qTK3aDh3pg8AF
Czqe8+AuRVaoAu25zN0NAfrrGXJJr+57uErCy5jA3CoVO7vfa0JOQJhFD4rY5SKaAL782wl104Hz
pFTEHLEdvHcXQENTA5EUtkW59/B1uCeZG9SNXRzR6u0eHuNdOflq7r7SZJiq094GU7Y1qx1xKLEM
+/t08T/S2UXxTUfOZcQC5PZWi83W/QXFV5DiPjipZzVPkfnUJgLsFP7nO1IH9J8EH1KqZGV8TzjP
LoP+MPGKTnFJYy+z9WFWAeegp0NZFrImnDdHn2XIa875QTOBuiuZ5ezlU+njAIYkPH3xfs6anZc2
6x8QtKK+MhN/ZoNQno8auiPS72r2nT6SGGiD2hMIM+9n7d47IEqVHvWuwZkPyqcZZi8dg+ZReCxa
BIHecv3zLlhsZDHANrseV9caroelxBWQo+kWEy0Rxk/KIFaZl1wXkfPXx/bmwon9Phm8zVYatJwA
V8Y8dUJBX/gXSNTH1mnWD9j/VzWwEYaLp2ZbJnvcb+fWqR2cEq/D8iTn1Nubs1Uhj4oiGb6NW1uz
NLfT1GYpJ5znYQsmZA+npeU5bea/Sh6Zy16XLNL4TRSq4G++gyi7P8r9qLmz/hPq0lvAcxIMlduC
Ed0Uo2gi/57G6VOFD8JQrNudsOu2tWEy3jONb2kAjvxrUKUBOUSBhLaMa9r8O0LgnbSUJN4iUV50
l/urDjlymMqzkkMLiLUn9gCxbD0xDuDGGN07blFDTmyGe0C9NLSBvnQEjEjVenFvmE/xWnOkn7NI
u9ddxt4Pmr0WD65UbTg+N6yKfpJdKHz+WkBEMwfwRpt/E4MVCX4Mg0aEsjIL8XEmcoHsO+7reDQM
NuX0VjCU75jMBGY3MfIsCsb2KiwPIetPfOQ6PiPvPJHy1R0Jl2riybjSuAiLmyU5OMSvFR8JLDTN
LPX6on3Ot8lYkeCq7yDRwkz2gk4jBg7o9NdYOHk4DSh6p9obqnRQBI7LlBbwXNn8kQmK0ksPq9hK
GCuSfiPBacojlTJ6szcxNlDzaWmywm5jbkHZzzehnTFgHuS3ypDEO5YPZaqdntBtpi6vr+W80XT3
vub/fWt17HHspq4QK2CrGNi8goA4FW5zRymq8cvuS1sU6vBqs8iFntjLMaaUPvI+Yt6m4RbX6w1X
2hQB1O96jXosGelzQssCbkp1uKRb3S9uwUSwMACDCOWqSBcbYZhi1fFU+FP0UBRb+VzzKh23qHpl
abR2OqvDzuAK5zaOWM32l7hH218evvPdqcxWh1BtgUoAkiyx5cjT3VPFrE2uudXmh0cixHjpF7EA
dLiS6G8pGxYP5+BIXGPyM3nQPkZkh0jJWFFuDIYc0rT4LU8SgRzUs/cL6gjZFyede4B6YEWiQ4SZ
eVfyjAKDHDhQWTxaWy8cdX3kC8S5TJkFBZzQ/r5bV3Goho6xUYSGMIpWmNI8FpCvy7fr8fNm2dks
TaqIEIxhuoQ9Ezd+bGFb0WhnuWww25BN4j75XgBNon/mMamYoylZEfx6VR+FOj4TyXANiYXm0j6J
/TdXKsONrq8/qkHy+z5g7Y5olT1hX6p+LpxuX38SQOXBQQjZOeHxUU8daBbud3xEYYIkY2hH1Xlg
/vTcPfumHUXgp5O04SNoK0EPhpeVAqNiO0mjI1j73X+N3SNLbhkIqU4/EluNQHl1Kx5xA/l5wdJ7
vVjMCE31PSSoYuNYE2Rzd1fYtvbsqMBeEMjaDsI10V8bMbzqoOAeoqnAWcT4ETCH1dOO36m4U1jn
2cNZZuLcc625Jbr0r5J2nvgHkbLWteeEWW6A/SJsaIx94VY7rJbQqKDja09U3ILYU2ThA1o0yTlZ
PtxiL/lfZ3VVK+TLnmb6fWr0BZQrjYVMaJ4Wj96fItP56B3gLV2NueG7VGWipA68obEK3GuPwgat
7TLta/xBRjakUjXa6IYozO28fJS1aFboj4q2VR/KV333kaZXnjsIcUvBVZtruwUIbFqd29SasDhL
k/o1eH3nV9wcgY+Z4M/MegLCnwk+mlpweh0BSj+rid4UZtt75Bn3x8gSkEkn6KCsrSpJnjHJyTWU
6U/yw3l3X0CUHMbM+qHXJ7GNBg2XIMkfVzfLSbWsK5ENG635N/WoH+IVxLt908vgPlot9stFALsD
u/mAnA6yd6owhn7ZkHx+A7IG3K4rQcciIFdZd9k5UJUwtFaxP2j4gqJioZTwvjFzFXW0Kr83v52/
wvqL6PlC90XWPp4E6bVYg7uo5XF4UNNVAUa2JRzdeVzKtxhZ9YK9pZEJq9kDuBw21aNWuFOwkmO5
GI/g6r1IBzl7AU2sczSbDMpNKuAVSoAp1lWTWn/ZLfUTzS1zxXt7TCL11rrOJeecfQNt4w4zmu6a
YupSHGdAa0lDTg2ZbvOzWScd5E8s92SaBlZyNwF411CvPHAhQvJbhNVULy652Q2B2Mm9AeuOqJL3
cmUQ8aBxSULFTPSZiVrK5yIo8KZGvPYvksqbJrdu5S+ILkfe2I2tmAWj+21N5J9aNATRpy44ozuR
hh8SIUAyoVm9zMUHNsyrJlctV7CoAkLREINWsFjBCuN86soSlmFPNWOmf8kGRbf7InYkZ1hkb5WI
I5tssf1SyqV58x+VteC29y8PAKeHGOyiacTJ4MzldFD/W1NcInSKIx2+k/cYIiaPIYlY9wzGPfXn
MwdYU+A37RhwaPfdSEV8CNwpDDFIOUNnQATxk70o2FSJ46V1n6O3jUaxPNyndoKYYCZfWyy8BhCN
nefiorpbEC9ClyrNw+yDKcHAvG1UQtYt5DAPpHclaMsZ4W+zgHqTiuLr/Ej+Ho5KpOYWw0zqIpc4
6naOtRiy6DqLETaqy1Q9njDY/AWVIzMFdQG1q59vl6pY0Bw8fc13kWCFQzJK7fur6o/NeiuPMVhi
/43pexSZUb6p+Kma3FND3QKEv0y4yCn0Qrjc44XAyvvdDXHieCMd6eegKYOqjFzBu7CGKHzMTjKf
ai7/iJpP9Jbg7ZO6m1pIKBal+EtbtGtVOorwORVjrPX9DWfZ2QF0dw2FVokqt1a+QhxNU1dmfoxK
SgJMWhWj93ra4v2c9RIkmvahg+T5qpJDb1advgW0KpMr2fwdUFwsY9YcRRBtkDF7MXQTRU+KmsI8
1F3F53XKxxILE+BJkxnAjVvcU/xy7d5XEZsSkuGzDgMp+XT23CSwhu1ZU2/vOwNnAVZ7xX7SBi4R
1I1tKcKSowJNS4IzIG6t/Sja40+6YAzPlFJ2jxBHsbX2sJ+yzMmSKWLFG+qz0e8gaKKxEJYML5iw
VudHliAmKFoRNBAfVp661RKkUT52RxINl27z0/DEJlqvmUXh7xxs3FEPt4BClWaRzXpMdZSvByIP
sAuOz+OhWYJbfs+WOg0IjQsG9azRt8S/O/dNe2t2D9VyzWCwOH79xqC1y6HXu5uTtLHQcOgfrolO
BW2HcBlEOabMmYH/4wP/Oeh/cEIa2sxlVBr4lACXEusMh/dTUSQlEbAknuJH5bsCcUuNfmStg8+0
m197YUx4pT66torh8C3BbVNXc3oH4qKBNIYAz5Ga+li0Q8ejeKFQm+jU8hAmfLGsBYdZxwagna3E
uM0ZfWIMr55IlirQeTO9uQOwMt5t5xq8kE4I2wbKzSuthaJGyya2yr1pVhLOSqXNHjRU+56jaTBN
dM8sXr1CliWUw2CIemF0ztOLOj8SUGPV/sbXKtrTv2/oRvz6DlBMbYe3bA251Q00J9oqPdJhqXa/
gkpgyQvSzWFnDU8hUVkG3l/wK7PDTI0uqinDT9tY8T2jZI4pHXsw6od86v4+CV5bCLUewoM+s478
Gz066cU2DXY/2POOzQh9mPi4QvWXOZvZ1hSZ0YeYU8Oany5FezbKvGc5JVeeFVveJlKJrnsRw0vM
oUHfClbClr5mOY/8gWURyWn3ufvNuIunMm4XCO72gPKTYbYE76eIz8Sz9YfL4slz55IikYOpHQBy
+T/4B1wR8SW8j+7AfhF6TyEMm5SkTZqQn16QRdYO50X5xycNt4sK9pBiaBs30ugdSeCn0UdiVqhU
1lSuKxAg1x6GcsAnsWcdXl9JD5A4NEoQBjIzyAQFBougnJkSXPHKP0ozZoBX838rPT/Swg7XRJ7T
IzXlibAfe+2tf/jFTZ+/JwJjqp1KRzXx+xnR10md8QL48XfnVnQ3WnC3MstpSawnJ3R+qZ5tO00x
TNJ3/LWC4Q5umHL7gIOjgna3GRk7GAWaKDGmVN9KaA3talp2LnuLIko3JAtNODdoNTXCdQYqmZ6s
AeXYD61qU6/lfCdGY6BvSt254ERvYyEVU2R6yK5zuQcVcn2VTcG97II9x6+68OwO8jTBPuWRHsH3
IBn9AuhmRcNrSCBI6+1RCKnsg2d0n4vKcXV9nCd+KRw0ytOFnfiP6eQ7bMadVTMdo+frOJUv4kTi
rBrqNPImqiB7KAsHb8qC96aWYW0WPtO0T+tIyYfDr8pGVst+HL4eZBMy9gU+9lw5HAUJa7Ya4zFE
tj1puZDCKqoFtFSgqDNERahAl7vGNOXfNP6ZlY5dnyrHa9RlfAxe44vZTwd9Ta1xiJ5NN8xZ7do1
yZw1JhCyv21++JcJojKaqiNh7bVraVPzh0Tacrb+63yKhKui8uG4/YFy4LGQ772cESFu2Qr5ZSUB
RxftOkLfd3UA5hLleAfocWWjPX52DNf6VsSIOpUg5NPtdry+6ymV/uF5WcP3BsbiICTHRr8Gyngb
RM25GjPY8tTa3kKgLfqkVIvd1dQ3tET/6wjp00TWDJh8VV1RNQC8RI+vr1vRPkidjuDlSsHIdwKn
an4Wh4YFuBymjtoTPZmJ1x7F386wMx7T3gGDjo/7R2lJ01BgRRj9vCY1cc4dJirBQ16us7/qoLqo
SYSoD8PGoX/bL5GbfchQq1Mo0Bkk5+a4ggtsSgtOc9QOPKVN1AEoCL+Ti99MBmRRwhQI7TlyMd0H
PSbULImctf0/hkifjTdZF1an2i/xW8lIkY19J8yQg0xJobarlWWcGnBnU1JWTdykFt7HjP/tbQ3X
s95iDfIo0ged21TL2ZRzKPnZdVj9bGSSiX4tLfQfckbAaG5HfsZf+5sLv1pc/PIcnLjQjrUbhHVQ
Y/rUKD0BMVHL2lQBrVLL94ogk/4bG7XVltX88YMOCB6f8odss6DRPw4BPGGeMiTk4f2ebSDkFdzX
cxzdfGW3hD95hKwmZm8HvSOD2WVPgmuN51N0b76kJSkEEVJK8pDjsZISTc/Ua6dqmSy13cc+s9iZ
MwMtZFaner5eSAYOW4RGEQIKb+Ezlgl/B8IyaaEIhlhQBWb6ze4LuxqklJkH6/MoK8sAmjpcyFUX
gQvgIL4i6qYVeqsZ9G1X3U254ozC7t0Z3TpFtN/pB4e3Hg/QV2fWnabiptBw4RcA+DH9PVpbPFvE
VioMWVtUjo48/n7UvFx7BwrLm6V8UuZgv95xSF8COh5C/rom4vO1shYidNaZcL/peIZmYGnBu5f1
E4Z2/7x0bFA2bj3GEIjrBI344yYPgQiewE2+kznNIvejZhlo8c0+qGRFeXCCcvkoNezuswOkp0Zt
cJaCzkMOdxCkzJGxBNYftj7DGh/DY7saKna0Alxx1XwvuvYUmkOVfzzxyoqBOYBOyT8xcDVL6sCB
rQj04xho4lFgjBlpmUn30lUQwZCvynXggoBxAyI0SZ54c7m9XMfaWIkJ9OjnLXuoGWuZ+E8pWzj/
Ny6Q9Qp/ysZyzUQjv/2s4HJE4DoAqu+ggoVUWcd3I1qOFgSXAs6swxvMbz8uOqU0+Ii/PXxH6xRH
XTHt3cdbWqCKpBIPN/1zqZV55cFyaw00TqdZAVZnpAu0pRsDQc9hSUlwTMGwzmb66nhASqP89rY+
WnKxLGzuhXhEaGk2VRLKyYjIYvv1876GlGFx2ZsjXuSpI62beC6eVksdnZ9Ss97Iq5XTH0HxZIhK
P1KWo9+WENyEg9vF160H63iaaLSYZe5YAe0M7sTfqkJqQVFMANACbtb0S3ee6vXu2+uXGyUQGuYK
IzuH4WvQR1rIdVLU8+09z0koelkxylatLfhCp9ErAfzrry/lpEQUAXEZPzO5aO6YE+BoxUTy4Qie
tNiwjH0gcXJhLWfCz2ulG8YH/nQu4u/Q4wvaiwxg7UpcmK0KYIrco+W2FgXPCUeXdnq+9AD7aDv8
QQjPQi6EEVj1ZITRHcbUXj/9sEcb7Wm+6PymEaM7RCcs+PNS/tUhXOsmYY3giPzxQWq5GMLlDPmQ
gC+s1CF/fR4WT6PPO/ddZSEb42rIxOk14X6uvLcoygU0CQoW8f4M6pZnd7q4qUlOM8D/j8cWJd53
fmnbfdH6o0WAwQ3br38ACXHFhFozcoMZdbf2shD+yFGiHStwF0Jbv/CSqCtqEYVEtFCyo06/mGif
BuBnUbR5vnzvfkRkYk9vv+0P7b1PYob+T1XPNQOSO8mAxeZgPYNfSTRcOH9/V9hrNnYhdFlyJkOs
ZVwFjUToaLzXtdncCJQdLzivxWrBJ/0hJuVJGd2rFHTSRC3FBYuJiNBNeC86TdI++/hsW0bjDrV2
K22cmfxtE5IeBH/vc+OgCIWrJ/POShsU8HaLS5C841t/3NIvb33/RwGCw61V2t5tVQUGg6ygkC14
Ja+CGYERBZ7IN5Gcs0KpZCebSIBcqwefIF2XyrFVxtnd+1WMc731/htkf5kffQ3b/KTPWjzGGVPp
+46IcdWpDPNhJ+sgtDx++UUKwkzIQMTrcTflLfZ2oUL3Lmi7tvVFvZGinYZ9Pzv62CbF/1UVhzy6
6hwKDo55gGIMFCDfhdM5i5K0LgtxQQAeKJJyYjqluXtT+AU4C6kzC+zarQpJNNk9CYS/JKGLYuqx
jSnR8vXgqvZb/4Te8EqMZyDGunbLQzo13+JumLPtZVDPnbmKeTZgiD+ILdiA2Sq9apgfKXLf3FHh
JTHc3kTUrUQ32I6434Viy/gXOEBJHMp0MuZIMtFpLdGmGU2JQ9XyRImuzyZcigVFU+aUb0E4UNyF
afSWzzu48dSwtOB5ul1GNB9+izoE+CC6amGiDvISv/B9/lpAxD/rD0N0mUkj2GLjaxqOa79lb23C
rBuOMG20dcmPAPxuv+pHROLiH/9jCi5HKpx6O9N4z2vjf4dnAiTlbXyLAlUfXFXaRXhqgh0sVnIL
z/hjZcRtTGmkfjVYDXkuR9BchDw1/m9bonoFMsp5cj1ZAQqnyBZik10f7EbSmVBphXiTkfFE+FvG
oq9hv9Z+J5VJy1VXZJIBc0deoLm7fOQLT9DSEGkw+Gar8VGNYKsIOaXnyu1ZNBAGY1ZVxjpQvTgz
w81lpOqtYyPUtuALYrJxmVW+gF5caXCr0kvbOsooB7ilXLtoR4xOYZLSi1TichpK5MGbrsR0zRdU
uxuH9ENde/e7csaZ+gqAO06B4xFERIS11KBcCva2Zbgs/4mXuLH/gN6NGFbikbG8+Eg6cvN56eum
jxP5jvlfYXe3BcUIf+6b1rH9I2FWTepz7WGPPBNVZK/EXflNg+96Gya0MMBkryFNbbaMMXJ0kcci
MSgo6snFysT6Dnzf8tSuwh9usDH7e0TsyavlD48G69xl/IVoD0oN+3r2rvw/Rd5RGHZCU/3ZLNZ2
7p8yVO4n34GUWcdKtPMSnhlI8+yWO08B+lxzBtHG8E6akl0xN/ydlN4KlpEJPJVcyoC4pW/AkPVX
3dqD1trrI5CJJAi2iRXzkelglOsOc0RRnQAHRglpCm3kKAYo2uW5DVSo1DKAnPEBeHjH2Is3xZze
kXKP1x80H4bCHRhKFKl1DCkJb8bQQB/XVkBO16xIVR8kOQtdV/KinAVcJ/l9BTcyaKPxLo9mXhZW
ZVoIV4DCAOvkY7XOnTk+JPrOKSsJlYyy01AToUn0PI+o3bSgJbx4cSBBi9hswyujPsv2Nc4Fpvy0
5k1PPAwcXW4Z9Lm4ozgvfLVVSTXQ0cU9bdH0ce7bbI3mLKp3Ium3CSsupLHDE6yD54vrT6Bu8SMj
vjrZQZrdgRLA6NMaCc0M3DLcwwYscboOW/QK6I4riqJ+OG5lcTIr8SUUKZyQG5Dc4JZusBPQhYQC
vGKo5zTqbczXe7ToDwT7Q16cf/B4vGrNi7WdOMqmKaGdcjXaHPtlLV/rsVqJxweq8sW9tn1KR0dS
jOj/yupNXF94yBI3cBwyZRKZFWxayw29DSAhtM2h8bfLVTxnnMZZlTAdLXGLrEAoVl4EGRS4SrXw
na4hmGfr/0et0uImKcpf7c7/DOPPJo2ZJ7patP1O3miH49JQN6r5UKyE6zHJRho8JHDKUescWNv7
Mu9tUrdZf37dDgoxglKAw4yO5+lPaF1wEu2YmAr3078wBES7S6cT5QUA+qQpI7wYu0WhAjaXvrmw
HIRAZs97SbB/zmtHzlwBW4C5JjEjOAYzhm08fkvo9+OHwQcKyEHUSgMwRUQkyWv2iI7xS6HzGYWu
iIY5OZYplt3kvrch9t7+n2GMyl2Y1HKL893IayzfOFRHM+QqAKIFr8TlZCSAx9XwWet6XtpecT6+
vmqqPuAu/ub/Yw1scxt1jQmLGcniNQWwhhSS1BaYHfEp6jkMUJ1ObnUkvEziZEn4SdnpKGAwPGMK
1dtNJyfEVngsQochQf35ttiKkJp/JOszmKdnDbnn+sanhXdFn+AXU2CejZNhVsIjQewEI+ETHAr+
W7zOlEO/4zVKNKqLey2fAc3Ip0fR3tzfgPSxjTi7r10lZi7ghIyJ9ja9DU6n46gwRwie9q4gXhMA
XDhJDYkiBVqT5eZHAg5sRndO9xezqVXz23FhGyTyKWOIMUINwxVjsfi6ld0JBJEStt091HXZC9cy
wRVW8rXJ7qRryDFZBCHfDXbQSSm/8z5IXsmbr7LReWHltZjvBNXRN6KFs1+2bbIaEOJPPZh/LUtE
8XycWDzkktFSSDHDZXa6VSMlVAphcXb35+j6RVukNjnZGHTq0lOBEbp6Y7pEEBvomYR/6XvcfCC8
vruh5ZZvW/kIQfE5elzUQKEQmnxmMfGh3Z0GGmDzSZqBcepRrbxmTWkDjfz4nvosTHPTzfqehR+p
I1ANNMQz07gYEjZd2NVu5IRo5faeMN5MGNEY+lbCgsBo51DclsEyH8S/IvBTFVDMbg3niOjuFaUZ
tivATmhBccsmF8GdB/EyWNMtJ8jlQx2Y7i6fu+YgyNXVpNxVHdsVqbD0XOcFZUPhv+wDPRac819t
swrOZylneX8EvVa3LhluQnSpPIr6hCcny4cmnOxBjGGTbRE3N6KblffmreVKdVfxn0xbKa8hSXOB
hVp61TPOa5J53fn2+iwAbwnSaa7H05tX9kK6oggKZMm7x+H9ffD4TrWZPls8HuaXYEVrZu8ThFi0
7rcZuDeBdrjENlbcOfMPsNyKF5hRsXamh+EOH2TOA0bOeF3f7X+tZXrwmnyGVTDat6i3ePPyfB7Z
vtMFtRyFFUO/IxVFgfD4SyWWlUT2vr1jlstoreyWxC7eVS9MyrRprlWYE9472S0/g1+RZEznKjba
nutff9cV+OhAmXfgmaYznq3+RA2Fs9+Eg7n2BCmMgaManZtXUt5et/CSgc6V5I4uBd5VlEXi0/I9
J4r3l2tbgGOiGh+YwGFVMqviaOFQSqv8EcC0HyIXC4BH9XuGdCh/twZUP7QWC7zLSoQetcq8TFXk
gfHUUX/pqU/2zqGRX4MniZsPtksDkszyz7hjTY6f6TxwRwAkG/qc33c8oJqpozXQ/wy6W3FmtGTS
EYc9uBBj/Ins7TiOjm84KnFO8D384F0HUKR8AWEq0R1SrJdkBfc5ih/Jbr4FPcZAiQPXFYvxUuFt
tf1z5UrA6GUxUIUQIzCJiz6ZPQHUZmIMf0buHvNxxegn8A1iBP/IVZTNkN7gswP5x83EMSimcOTC
SjHNgL81i+mJicHBe9RHTRhC7tHRaCuiIWuvAvNaLsRqYa9dL7VrkZA1Q4+3rzFTc3O8dSXZ2Xvo
Uptlv1YoX3BmrV7jqFfBGrmKw00stbHbktiVuUpAyk+q+aZI8mk15BBbQYZtyS9/06A9vOYsHkeg
W2rWEsAvTFp15Zgg3JyUe82VUHeXH6FulcopiJ+F25+5ieTICx/6/7DrMMWNuPoO+4+P0zPFOTjo
uJ69BmO9WH51C0tX4GBPg0w/CHV6GRxy/E01g3JgrVzmPI6fwG2XYxMfUBQAkaTjVoJ+d796sYT4
7epdBhdeJpm83q9jN5s4+9VkxNjjexJcz58Jwgelb+ji47nQEqeNqjkScXW0VOLjFQtsSLkn9+eT
qZ6QZIP4uvgZAnwdw2Doya6XK+Nz2RYUe2FNTpQexC/KWNd3Umr2IkGjJOXN85O4mT/raSE9x7r+
VfNo3gmjLmFSozeskoAtUEbpzd64PTi34b1FcCthzsC4vNfw2yPArBbi12HLVkm+r/SSVbGx1+47
y+HBcu9MI4vFuXMhTnaLQW5Tz5KCP4B1v/vTpqrshYG9TODICq0qfWs/gyoYo0LCTzJTvcLRFmy5
1cqR59pOzn4Dp73HTu49HwYuAvyx3hyIs+l5+WknhPG6Ygik/XZ/rOuQl3zhdCb0swvBNhu2peHW
XuTUWcJws9k0LBw9dzfchwzbcEqsOrPdNKr07O3fJ5bSsnWKWF/VoskAB/lBDFpM4uiGJ+MgXdnq
P+Oj6eZRAzmCcmeX2d1oGstjwzSnqv1Fzod1S0wqTA9XGoF5ng8vp5w56RZYX1bYtrNoR3ctqx/2
bwUrd410Eks8Fs1LIH5a+QQ3SoM7B4h7MqhXzdamflePG0K6f8+ZDvrhl2C7Cby+kPlpXCr1QDbZ
3oF5cKFV5OlIGaYFb4Of1kkP9UxVUB2XoDojT1u+07A4/DRKTBbkIk2FNtWMNWYI8ujS/QJi+64p
AzVQR2F/N3tI8APErenG0Z48coIRWxgPil0tO+JCqi89GywBPjR5Bm73cz9sZHuicGaIMi83QL/r
dqKncn/VHXbfPweNZJ+cWt7/+6yAZQ5cnVP80shujV0h/OczA49IhPWvZ8Dh2iWiU0H1Dsc/EIoV
eq2VjoT88rW6CccHfsWpYYc4efxY3T1PfTVJ6Czkul2Qushso7HNZnWtRFWuwukuoc372POpQgf2
QPyo0BLGOuTQ9cbTZQ+kEsBsg65gE1A3MFEmm2hDd5rFLZ3v/oMPGy2b6eXP//sy1jeevtZ95sCy
92pxPxRnPZrH9gzZNWu+O4lW7LD6eYes7G+1n1PUoWqp8YkuehZqsJLspKK9h526YSGnnj0kMpzV
C5/vDAyDaBGrpMZ4laGeAu1+X4ZXHZxPaSKKjuU8fB7gGJIb6ppN1/ke+JM8z4McvQUHfqECfWhj
e897vMQ7LDxPvlHQYFkcNTIKTHOrutKGxR0y9CdPeGNXVCNVXhg2XtmXTYOJU9Zx2fg8QIqb/Kte
NyAWDcShZnf6ID3tAOFb7rbVBcrAbc5KBVcdZ2Be2rOS/OZJyR5yDSX92lwSK4Nt4YIjEQ0wALjL
pVlf4mWyEG7NoLJ/b5NHdSNEqcCcgxpg0hs8PvZ+J9Oik722ApsAYGnAyHRM3lSRDIK53pIz7cMH
jcpsP/FYy0qSXYWevEuSBMxACK8OOgpQtL/4tQeAPSm9QWp3eWbQ2OCaT/NKn9c7K/WdlJ3P3XoX
XHTZXwhRzdNUVsjNU7FK6Ve6qhps8k2wUhG3pz2y+xJVNJswzwryXt6F5yc+4LeCSgeVwgiTrA7a
gx2IWXbCkdsJnLW7ZuBLjSFtQNQQVCQzsiAe+s3q2hmCmXXqHxJXfq4TF1mmRY2IfFpFjep8oRRL
26xaCuOvcbJjcZj9PwPDKH+zYq0/CCKZJK4//tLKH3F3X25pIsjXNDOgbSS0JB7zMPMCwgkxVmA/
8IsDd5LLKvd9tCpPaTtMdBTzP/32uXnYTl/12WIVfQzlrlaUuBHiAtut80p/Lg58BI+KUeEcuONn
E7NRTtvdPT13+UHuGIOByuqDGMWCF2gCnpZT2IvtJnXbRmslXET6T3Cb760s6b7fiJNo5drI5NF1
Rnuo8uR8xYmL5mv/TeJI+fjncrdpcXyG7Kfb5nHSDUZJEslM76wx3ih3F5sZ0iVqM5w1ibqACgbA
QhL2b0cO3NG8zAn2hLIUq8yaWkEror0ALg/eMCHIicj3zhqpDUluxfz/ICzFmmDAgrl/1Hn//UQ2
M3xiGRvZQACB1sTxlSK9yktDwH9U7mlHWXbAzMc6RzPuKZvq79vLDCdyznArN30aL+9S+srNt3o1
jWYE6qHIgNLfzK01v/MUhVGvSnSz45UDW55R8NPbJXXa+YBxuofQCe/FWiln696HJOcaDnsInsyG
41JeNux7mFDR7CJQYYN80kw9GlTeuFQ88uaWqjTZ+KPUbpdIZre7aIAS+mdg2mZVthpKhHMaHaGw
CyWW2vtpjSULh+UQVa+wmR08VzVNw/HLs9u2q9jT7R6cUTxaLFVMaVCqnyoIsHAURc6R6yV733gY
ti1/9A22mX9NNm5fzKlEDEjtjJBuleYRPki9Frc8ZFRfKrJm/Zn/oGnXSszyDqF6dDyDvBSt3/SW
XyNv3cXENjKt8muCgbn9UibK0b5JJi3HHe+i76yQOe7pfTu2HWxIXvcKIpzB10/XLtFsv1O6RydL
kG1/VNiYnVPrZL3gPs4yl0qB6UBw0cJI5+hUrIO7ymjHGuy4I/ArOi3uYKWdiyfDa0GGgYxRW5l6
N1HmYtMxr4TC4dDokclDFcp9nPqcSBLswJzATEfhKlOCWy33MMBnIjV/2gnCm57fCHKmP6AAhi3u
bfQBfaZu62YbdqCdBl0+Q4+9huNMwb63AlFZwG2AK2fNjPGd68nTNpcOHb+t5VP5HIgPy89l/v24
cIggTu8vC0dUhHZDR7K049ImGunVYYm+RsLB1IOSaRTv9cW5jfBonjiqL5nZrNI2rbTRKQ8WO90I
CFXR7WaufZkPWxi+dkeRGcRhEQJ0lVaBPIPqVPCOvFIWV5u2Wz0Jz2yE8UCW9iOls6ROjt/8n1/5
pYOFGam0h53P2wdyvQRzvxN2ElO35r4ouL4fBAWsEDN+lzI2dJN9AgmhcmFWJDdTRM0YSpMh3/7c
xgt9Is909swP0Up8YRZ29lgNlnqtnfrJAw090nXwDTax6wgTqWRwkhmPtE0VAxOPxoCeRpIR95NP
GkU/4TYIMhJMGof7MkvrAxPjG2vIWW+CZkLhKqTzSNiznVUBuRCgIAYn22zqvzYs1i+RqTn5Up3e
6vsrU9p4VjxBjlXlads5/aQ//lWUB45bGwL5emaPW4xy1Vb+DPglehrq2dws7q6khIEV21A1LvkT
jlMqr4xb01/pnYSgEwUI4GNrt3vPhRNkMyLB5KHtvxahvls+zoK1fJ0iwFX7u5mmtipSXjY+AJUX
So9iWlX+FFu+2a5zE/OAGy6o0STfwqBA1tlx8kqcHm+scYaW5CaO59em8AnkoLftC6CibKkV/qSs
j32Nat0DjpVdkHHrpd3QU4EZWORW+CdDSjxYyNCDWtJxQpZo6UhvGOawHff5f+ckctnBc/EqHjm4
WIylWaVML1Iz/49pk3t14yoT8giZH4T0sjG2XdIfQhG6VfP5sZfDfr8W7TauJ8e+xKsF2BtlrMPa
7rz1AHeFN5CTd8fNsIwSzvdYlBZmcvDGojdmrfbVxhHWFgqdPDlEVTkN8IIRZcRlyyi7uvkqcwrh
Ouq4kOxGshik/n2V/BmAfX72Y9duv6EcVjp5lD8EMpQSan8p7DJ7RkpXE5ea2f8LZHuoEpKkAAyK
OxNCx5z4D+l8iaPbp7wgSObOzUuQkQrvJpKa8Q7DZoCevLGlREGQhlVsgQHxkuwlehu4ji8Detze
MGfIodChLN/riD+7/RhaG0uDtbOsYJZJxhW1A6Zj4b/lYivGW0hLuCcu1/CtIQmFH1h13JzVQNP7
BNeyBK/jA456G9tymYx46ST2uz9/m4N9VQJmZxOzD4EUr+Bw0LmEWn4WR/wL8hoYU38oLmUYbE0q
1QGUFWIAmhjWNdnJlkB5VceRE8zliFuQGOJB9CDVto/iaTfAW9VGatlq/BuVS1lHUsWPFh1Rk23Y
a9mylEZG+ONiXZROoAbBK1cT7NhCJAK76FXjR8e/u95XNkDTWCyuqzKbHqS4ZjC1rJEfW1v05d8L
L8MrJhqNzs6l9uVTzhNIru/ii7ar2TH0rT131ScCPYweCu9+g7eq/EHKYMK8Es+s6Dptob3Aw6Wf
dcetRQvMdc+5BSrjYn3DbHs14ba0R3zkTHqm63MGDg1Mxd0tt66bseH48FeheRQa97a6bqeUjhrf
OVAGZqPx8a6gYnNu2201mwXjXPmjQEAlSd733OqfB8Mv6OEaRlnbXLIqXZiEXGZCXtuXT5x7wGyy
6U223t/lVo1VLeA68ZQB5QY6aczzGkCoxvcjBq65loiB06doBlNZkZpvGXp5hp8TJfSSAQdA3FaC
qMTqbe7J7PilddRFRR7fW+JQOWb43pZ8LUl1QgoECFl9uBgyYnGp05MxDzVfrthfzuX3KEex/VKb
J9zK1LJl2ofJxWcB37UEP6IGtC4DgnBwspP6bgwTiX+D+0laKv2w7tqk/C/JV2Zdu4BxYZ3BJLgy
ttK+cKMG90zAmMtSzXBX+9RAwRemu2sMCMFdPiOWuvkA6/awdZWC3bStEi0aGg6+pfim/7Je+Y9s
VeXbBnuw8NowW0yhn9EVnAVJZ76Isci2V+BBY/I4KvJSOGWNfRRnKYA8lhy2qQmALloe5/IFR859
bx5kVtbN0d1n12tBodDsR5PRyvi2Qy3PEDPsJ9XEaW/8HQoGlC2acjzfGmI6e3J0SDSE6xbapdYc
s355drGkUyh7L7xa1GhtZGX41+XiLAkoCbPypXfth4jkzCxmYi6hb4LYjatKagLlQgmKaDIvItxz
3dnHV9d5aJClO8LoERDdAl6ZCo45f7QPfSz0j1c0rQF3Flwtt0LElz93Af3umR4w1SmRq/8lTMTk
hhNSP11FI8+wS4wUIE1+4n4z4DoFq3GXxBH+RdvV3tCLEZ5xdBi/4s7zK8/bOgs2gtQRyZ6yZFpn
epg2b82CXpbD5NX6ELLyr9y2PHOlkgfp2fPri06lAiDxyY9CY6P+oyQ/MQp5bmnFXN2tCvTHaJFp
KJYL3CBVIqATpB0PpNJwkwt47xJ6nuEIs0H5TevuSwixkFJMGJQMzAOlCtdDiwn5HHhJFzAol7OU
KPt81VGsgAL66vbEDobXAwDZN33LdaWOfdmoTlh0rL0juk8czg/904CF2ZSvesIujimtNC0IkPvy
KohRmmFp0EydysRW2adhwgA2AZBZ+GeXElGOL3ZgkFB1xs735HpIzj85Vs5xybMtK/wL6oxf1752
WmDjcIZjzDjgyKP/basN2mV0lyGRxNswVWdEMXxwP1rHAXeSJlkD4Rv6wPRd+NQ2OCLdJcAgwyTy
NSxkOL/tFecJr7WG4/a6PxYBfaVe5nXbFX906RrvBzD15H7jC94S9+fs/GGU3CG3w+4r4Eah+6Yb
OrG9xno1vJL81sNkF6MpxPEwgO8HQfHmZD/XId1BHOYbsr4SozcJZaM5RJntnL3JHyleceULmxZ4
Zt08iDPBBEvb6GYfXwLV1Mh9FxawYr1abYWVAe5U157jFPhJSdn2miEEkaNjDz51FsUwVgVHMM8B
me+2E0z2NgLEMwfseY+vcn7AAJThSqWmlrinAglHvlv9tA4PD54UjKXnvF2p5bXhK2ggTGf13mx2
+r24V1Qo3Jy9hX1wOU4WILcfA7PQaRiBHF8RjwUAiO861XbtCpKX9Je75uwUCtkGbdKWSS472byn
E9yPDw7aFQ7BdYlKE1lfiYL8sa8rtOeIxD656uebJyQYsEnVa8WOBFEyYTjznqpf9RTjeBKMGfBJ
YcDyGEw2Su31z0JFWVZZvr7sv3R0qhhBBXSdCJg8R6Tti+AaPAZZqKEcyXZYOZ6atOEJGqxPSYp0
+7EF+1hi9cyBOzKTY/cGjFDh9mLRjVba9MiYP4GEeE0V15VLDNCDWJhAwryE2rO1j1cNVhk0IX+f
eKUl2YW7PB4/0+5MKSdugHzQ75Vc/WcnLgf7bvpOGMxrqjGUDp+oTmKGIlK4T4pgK5Km8+a2Oh2y
EjN/XRgenZSP5lmRSjkTOoSX2mVEIR2WGYegRU//m3RcChZExNxSs9ZZ4y21p9JmuHBWYIK1iif1
VRB0f6hi4DBNAk+G1IgAxE7BPJv3gskVSPcktB4QxmqT9bSGtcAEPD3TjG6C0YrE72EqbbGIvuTu
r1PsaahJpLnW2b2NDB1jvD2su+eiDqZhwjSeHqnarJD04mJPIwFnDZQYF1UQPY4xHFmYQtc4Ugso
x3MEb6EgwrCvEBjifCCeHkcEKcHDC97VoHMrVHlIQgFO1XjKBGB+zFa50kHx8scK15VvXca00B8j
Prme3OrX7VDLRxd8sza4cKQJOyDmnSb5qfUxX1zBZsdGv6tope/L8KC6X2uygtKktJDxUk4xotzG
YRREvDU92hK7N3WuwPZmdt9Y79Op7Zsk+455IpfSM0U0veNROgD7kfQGympfbNYJJg0pbAr306pE
Gxq9uH2dFZD7UdSn/K41YhHyuZotj82SNgsd2YViv7d/bgjpOipfaXAiQiXSKf4d2fdHpWhvAW+J
JmrJM5R7uDlYfUFiCP3EegdmhizuqBqaFzw+OdZ4zVYIkoZcHbLi4zd8xyK5s8bIZvwy8uJFH1jf
hIxCk++IKMSxAD4AbOqIp/Z5/h5ZDYZs6g9+++11uJeDyx6JuWU6YzivRNJ+n271AEueQjzGpVz0
hgUgBrFiLeetYzP5KK9pbfH691k/ppQnNjt7/mxj5UfUvuToTMJ3HkXbEB/3cvvhPfuC8ReDNt4d
4jd4suNwwp2zUpxwQ8+KzK9uBseyCyiqJwt0pOK4/3xuOE0Wl3H7zn/EHanrQ3uKdzHv0DODXz/L
KuimSzUFd+OeLbIHsV+Xp9kdN8+/Oeorecx7ROdieIhynkf+tcjtObQwczW3WN1zBPIjc7T98wLL
Xz+3dgF7+zQQeT1AKk3EypnJdV0/F2nrYdJvPExhUnAmIkVyQ8pLji4tdwAnW599H3Z24xzIBLth
X/rl39aK8c4fxJMHwEsQLURsCmiaoUSF9LOzACFH1oyT6vFxRv72URlNbRTajODEYv/2+1P90F5G
LHS4NKVJC8BVjy23EN+7Lxyt4m8y47fIeeG/K1TXGTN49qlf5tCY+yuC4Op2loIlVrJOMDO68bb1
aqDNDvv7vFEqj4f/Q/us7Q1GJLlFfA2piSZ6odDq6a6lNynlY1o9QtRn7vgKx5Oc/ZjroxUdW4Cn
4M/owN9KKPZqBtavVYjD9LTfUKU5AVBW4AaQb6FizK+yltrIm1vxLDLFAjDyiEQcxWxsvVTlsn0R
uwPlq3c1ghI4+V2EF/PrgxD0BR0mqiqy5Y8J1+kgaiawuCStVNDFUTPf7KNz9dXd0jCdNKKebiRW
5NpORmW7B6J7qqnr6F1qKyFq/L9e4eTEykJu0fkGD6rKzWAf/kZoRuAaGpZhkENuoz5Yke3mix7P
3NlTWz6miAbJuUiceshc8WX5Jc1HmdPc40SfV6EAnXwjB/Jo2gGaS8JPetkjcbyiJnXMeRGcreQ5
Z0pAgmQCR+xS95O6nBvOZ3ol52ClB6NDCn4pXGNSpfY20K/qH0JI+ZEDY3P6BX8ENMOudPP4703i
Z93Sbu+rCJGyJVCexcEEbqz4ElKDVEXtFNIlVwlMJmAGbQw3s43kI1UdwmrPePnx9LDzUrDeh4Zg
5e5pPt8pw+zYaFvZrXx/baaHJ/IQQq0s/H0vfdtzI3SAFPxf7xu7g2OucAM9Ufendt2kC1iwLchp
eSPngSU+wLIHVzmUSFlxxiUZTZeGBnrBqor1+crZnejUgYnoy8rsYPWOCSGcOwMSg8i8EzuBTDYo
lrQx1CAHtC7MdxJmuelAcNtDrpWqiozO6p3tJJScIGKQQM25G+jLv2/ep5mWs7N8Bca8tjjavOpq
3jSHWKfYNSbgz3OVqGufYJXXp1jWCv1l3nbSA32URftIEwqERlL3CoIg88TTg77Ow+1yejmyWp+t
szDRYs9Nq6Y8/ax7WxO1VK1B7ohjRAnaeVa5AgEEBS9Dp/xDvTSUH78Nk/XCpoTqvKrnjFa2/4Zn
bPAUryStnEUh3KJQrOr3Nhrm9dY8VZHIsNRrAXkdvdKUocPmO90zPQdOZVwmEmwhc3GqRSpV5h7h
oDKTWaiLH810fxWUHpjk0kC/JVIY02POYurHav2o1q+9VPHz88fUCgegw0lFQugjGmNEzD3KPD8G
KcqYy3PVmQYnNY+3RForYN9Eb9CU2mK5OS+y0qOtgu009OpQen3Yl7M9v7AZ8rPNYemTCjjbRwn6
vrH/wcGJjcLJIhzhXbauTbI18H3GupXc1BeV0+mOPfp38PUbYsaeIBRQ/GuLT7/pY953LZQGWjeS
9aMgWbvUBsEY1Y52VY6DTF0roV5jWMMJTPgVZVXpRZuuCEPjuCjbYvAyEdMQBaXzih5LDAniWiN6
/uNElNsYUpG7y5ZeEnUOXx89Y6cAfUCHgeL0KA9xD+mrPgW5cOpc2Nnx8VSjRH5utWAg5DJen5dC
+ZsdpGpvmTACAIAeXxPG/LUKhpMYkWUYchwhWC8KOdz364IWjmUQ52xb4ibLIDcE/PLU3EGcexE5
JvbvoMVOYts927Bc0g8+dPf065yQnoLkbf8+aHGPHNRa3WI75dxGQzC9y/6O4PD3Sc/gfpNjzE52
xDBOGns9tN5buJjqGMILawU5epvT9t7/gOAbTvdinX4OP72llkThZCDuAi2zsWpb5Xy00Wuht/0W
XoGMs87CTZFv9gT/Ays56rnamxseMJnhzCXtbtj0FGHrfL2kVn28r5U5xFfEn/f+bb2r/BdyE371
1MpVeA01eWwSbyVKKruZKeznao9zVBca1xy0LMHH6m0+VFHNG8eKTTsnP2bYClbYcfEiYW6rFmzr
kddsq3JJQjgP+NaWjlXRG4szAjdAzuKV9noCYuLZ4dLieVe/pXQmK1DiUF7y48FctnNWsmXh6yN5
LI3/FBY04fiTJHv/3EDB7lAsaq5+kCSWxt9ATY0LbUr1+45qz6p0DuYBVjB+P0M/uDP4pajeLtpy
6w7Di08fz1NT/vUQ+3HXg0V8vj7YHW19iZuNDVk/WKRXDMP3r7NYUPpb9nCCtchEMJlvJ+66RbSo
n+9cMTxsY1ZCNZQ4Vg1p6W9zxX1S2fGS6iq3Nm+QQcKn+Lcsr38qMyRAPFTHA4cyaxSdMkzl6cz3
CKPt/Zn3MlZCo7dGw6rih4t4sulDtUjdDBrnOupnXnOx8M9hQtCnfspNj+ihlA9OUjz1aVS8nYuL
s3+fsEH3qg4+eMrHKA0LuFYI0FfHJdfffkWbXsqKEFbCbKieMmYhFYXfhUetZf11NztY4r1JNqve
Ltu9zxfAvzN7KPOTnEhdgMkPSqGHSfD1CRa3H8zl/scN8c1hoqgxlbaL2r5NGTn03CegohPEhM31
F7kXAzvP8vkhoJLmXkJnJB0x1HiWfEvpz7IptTQzbUkt6s35vFcy16TePouVJbNhHxPz3OkD1Nuv
Fpfgz4c2tZbmj1qHgDki70EmkpgG18I6cPfY9Ufn6ekgtufEKC3S0N7Q01eOTnmtTJ1pwfWDi1JO
9Wf1UvFZecSFDQ5q5CN9EGKHYhxOVtVzkHdktBv7EkwcouU1shr9esz3vLNAZnMmahPDwxZH16eY
UI1ga/OtxfjWiOJmpVSuIERt1tjK+Cs+gqIo4Kqb87aBX5IE3koBrSYa8RRVlmUCU+gGkyQOX52G
j0q+G4XP5uAk4Nj4JKWHLd12UlDoVl9vaEAXX810XyYWRERlqcx3YN2ybOkMqyicNu5bdKzcBerG
5G8vCG6B0Dovif9ewzCR16Cj+ZILmJSmXP+ma/DxJgzS3Oj1tpoy4quJTAnarWizlMDyxa/FmcqA
9LKSbG7EsQ7dg/jVdEGwqrbZjG2ozFVBKcZMIpNOZBtgc0luFdwekv18glvBrbIeqLhq0c+92cu7
1kUlvkadhxTpNFBmbH6l8GMvCVBBhDzAqEZ9ukfL5GPJ9UZiqgFf5xIRBR9tIWUYxfOqKj41Nuoc
OZnZ/UQAcOzfKDBok5qMm17/ZysaQIvO44pylnXs6rFjprgpqHaSqnBdKpDXHYCNbsiEPL9hweu4
5GOHkeb0fSYcu8BmX1Jn2dPpr2BR8UDBlrmDmVTS53ZApXaGDlloSdETkE4YlVpz8b7UdzqSErUN
YrFIEGhEHLRVbSDb7F8T60RDkXd7LUBEB8PAnL8dhkcKCE+UPobBZz1VIaur7lLFop91Ear/knVx
yQhZNLrGm8nrKugv5CIuDvLsvpG/Y7IliolSbOeo7au+9FI1+xcWBA1SKCsckLEDxtlBgaA1O0NB
nZNgat1+ffruNaceSLaLcs0Ir447o0tWo6O7265KpDAYSlA4ZY9TkfcQ/Swf92HcthiyP8znRj1+
cSwu1GJXKIdZOZX/IMXOXAKnXd8qBKH51hkVj+3C2z+m8j690Viym4IemqKtp+LIKk/QWPSb0wPt
oIhMX9ET6spANr5QSl0z78JubpNdTA1DlsC3otcZQUVyBCk/aKZIhqj2rD4qJq1hTWG2N2cTU6Lo
BYuqUwqgZRtXC0ZjZYUt8PkFNrzaU4Q46NJEmz3Ro90x2cJ5ZvuE0ZqoM4CIoVpwMRoD83G8QjSg
LWB6F5QHlxx5F2nWUOAYPmv6l28bjDHHG5BWvvPN6aXuyick6FU0f1al/XHqys6hdYbgctofBrdt
FM1o/oBkj40FKQMUI/hafmUTJhTAlobEthHO9ns2k8oePdIuPpyFOVMhbOrcI6vBS5ak5i/vGAc2
QgIRwC1W0egEeetPR3qr8WMr3JflbH7Nfto18EdgyWo9Prl++sW6LgBUE6cbkb12lmQZnUOMQ9Bw
QQDVNsUe8n7b7PLBfgaCEF74d5QurfWA3fedRHdEg8f/ATohzrpruRM9VDLKcQqSInAKi20G67Yp
surnDibxstUFRw0ivSo42USrDzj3FtcoxI1rjqIrtfvSOsecKmI1Z3ykyIGw+kJSJtBlcLUSSq4N
+C+8WIiakgwld9sIBGzrRq3wViRTtx540kwVX4HZhVxwTsuhaJTgrl1uBED26564FJNJMf68+APm
6CABq5CGXCHiPN2IV5fkbzWv6bsTXxjkl0iaX6mkKobHQIZ5rfGcnIqfv1uHi/fFLvYbeOCtL4+4
5UU8WABiW+tUmZrJfQcUOQIYB3g+pt7AIUTOYxqvQmE9FDvHgWGr5A74VgVmqSOEdVKoNoYenxRh
t3D9Po4QB4yJdv31dZj43Iamrv7WjKGCW6+ey/gv7lUWKAMhGOY2dzbwPgzWxB3wlvJsATRQfQFM
qkYXO2jayUnart74yq4You+4+sLYt0DJeVzvDpKrjLMWwATRE5cxnStCIvh9l8pDvsAATcNypLIr
KuCcckyGHz1UIkD1tfnk0nUaqvcFPs0Gy2u3tSbXmfFrXr61ydLr5c8gESYukt4lVedrQaV7Baiy
y6xz6nLQ4RJc1YwGmaAuYyoSOFCT6MqaIaiL4EyGy1jSwnNyq+44zKE8GQ6uq873yzB7yo7t3ULb
74ajcGwdkpDTVV1YWrYC2i6GmsO9Vs+Bx92bXzCMtxgEICboswHXDYHAM+n8ywfigs8Uk1ffDmsc
X/eyhW85Y95/BvT39Hj11Plz+UZOF32UGor6qftT3xJVuXK8KYxQRu1+cHBIqI2Dwy8vS3gBTSC4
tEh7HFeXUwE4eI4fcmA//GcOe+U4VLdotexkwfjr7eQouvBSbH+1UMVlhws10SPP7yzT3mU9aqkm
8VBhNNlu1al155mwfI/uuCbumBLBsrIHe0EfM/cJZou40Cf6YfZmHq5afqGb1fxOCxm8cHlTbIlE
hG/CeXKLRPSvGvySVjG4S0gNJPiSCgeV2DV8RrUT759DklPvvGtVsreROqp80tgxSlKoVaOaujSj
3b7pU7lIjVOGdC0T4I37bLdqMx6oFAofeOITTxG2HwaMSEYr9VYCqMTvTokOZwp0UQjwIe2MqcMW
liIKFf5ibLIensy4x4uqgKqa60FzAro75wJUKAd88ApRi3/Y8cOvLAk+ctfsL2y+Dq/lQRjoAUI1
uxdOTIAjG7sdFkD/TRMdeYbH9nTLYxW2HcTvNE390dA8gg+JwYvqpcmRs4OxIl84r2uWzMYDHkvC
sWU8+7uscgmK8VholviNi8JWLXzp/KGFnGbnDD8CeaA9ETbELNXIeHHjUTEgcL3hNuwpkGPbDJBQ
lc0NYYKt2Om7XhhbvLEQw+7skww9KjEzrTnu5YtaP/SP3gxkvkcbawpo4Wqc2J+JdzUmfMvYu4Ad
qHw6xT3tih/+4fHBkUkll269GAl6nF4FXzfh152ZZxxNLosATlV1he0LS9mvM5/I8iPYjXrRxfyt
B098Ryctp6lbQMekGCBbWXkr4iisJLWaQio/Hn1HILRL2Q4WLLcWfjEratIR/Hf3lRFmWr0riAuB
7nf8hP/yew5ZdNB/CXzaJzoBW6iRb6YkLIbeDh7ENbJIMRHNqXwfRnU+bV0wWZSCFfRAoiqT2YYj
Qlgg93jlF+P0DDUGnX4O29syz8LXwqBeSNx5d9CidBoNnmYLdSQU/M9FyORmAuDwwFiCpwds4lor
3vnMsGshOzWD4lHbBO7HzU+bqmGTMNhdhN0kBJ84YWtC6d2uIc1HHqbBM9iwf6KMFz3vdXf15qSo
mGtFP9bXxQ/JewF9ZnyAu9CMwgfSC9ixCIMg5PnHrlBRGHVcI8F/dje2xYq51lpABvSfC0TkHv1c
bduW689HrWrX9n/3JekTvrcQEmqFAQ0KuK0IzIFdecUhYX+eeWmTxa8MdQg3za928kS7prIE5u3Q
Qdv1JTm7qk5iamkcFSYTgM3lUHCThSURR5v9oq0hJNHB/q0Ej1Axhq2vCNYJdzR+xzNGBk7wMLx3
QcZ4dBaXG97XKsy68DlWsufQjf2Wp9FBo6C9AMG8sNppxFfTm6TEIN5P8yr2iQ/G1aEmyGE5SWW0
u/duXcDPoOmAbOGPnTEKD6l0v0hUCFJzfs+gJDHwJ//00NovvcCZ7lGjwn1wUa/L9uwtEgLLG0d1
HJ7cxtqQi40Qic1YTJKaRSeOh9uMLaS7GwjU+aFL8mhNGX0QgayndG9dkbdiFeJ3aEc8evHCT7NX
BIG5gcCG766pqNHlWorZ1BB4z6WN01hrL5brPDHZIKcvE2U4BSuwdq5M59q9eylbzNILp80uqMFl
rBUpj+nE2NeIGB8eWBgkFF4TaMm+c3JE33E69C5tSVgrzzniUC2NufuKO7e+hfh1VWbuMb8v8n4m
M5vrEoYl6tFXgFqmnGE6LUTmRQ20N5+ByXjXAw76f6CrDjbLliF2Lvn8s6A1U6ilB3V09ab94j10
LF52Jgs8/hNFt0OoTHW4VK6FTqSICIHGo3Qp316civu+SbQ0MPB16oNVjS6pUhgmiUg/bv13EW4P
bzlK94TUKzB3cw56LII/Vx8rbk7aysUPPHqo8e1e7I6liDffYdi6h6ogn7w4/dIWWHTmq4m8v+py
BN3a1nVy5ClFS6BFLUU8RxNOTbA8YGYRgfZExLaedAVZLiYtTv0Mg2K+72TmBAkeiDbmkL2yktRf
OfryP6SXIQycr3KALV3KT9HB1v2U1y+wnu/QMl8ThRVlYIQ8cAKLWsSwnDA0BQd3bdvKeqEVdXDU
f2VFw7ybhIZZepRf5uBbjfJGW9cMNRRxkmtFKj5pD2d5xBDuD+jAODD2eDw0fP8sOHzqIccypMCW
dhfakfMBPnHQdxtZ9AtD7u6cJPPWePXf15fCuHrODWtIXjmhOYbNJpQWEPyQtc0m15GYoWMtaVRT
3+RQp2p+Y1n8kGc9zftJoYv9kCTvi4+ABTdCojPWzALJbAS1guc1WSPNS3HUy1Ifxu8lwqzhDV/F
JCLK65QuSTrcpGI/kReER7Cb6rwaURpeUDl3iGLqfz+MAMRvkRFMCau/Y//cmu050JiBlzyHmQfA
Gzp2mz/LN7LiS7g8V9m83yVLTg8Bp1EJkIkCHdYZNtFXp7Vv3EHpD/OlfW7gPeyi4y6DWKwaZv/q
UyJt+cpuIk9Rn6cBLulbmZvsxWfzMJ07fg1gcygYsXIjCG8N3S6e/JfJuRYdnsHh9XQgpwxILIrV
rC3yVzQzD4yc9hOq1618zUQqpDr0LnDCMgqOKglJfepCLdhDtPUCq7VEZ6U2XIQUZQlw2fk1pxZ0
hG2G/Qwn87VuCaKnaYSvxP8aLL3EnN7lKJiSistY08ZzIKtlHaO5ly9lZmp1tOfOumVTl6HM7yTt
A1Upsdox2QkT4d4tfVbr0+cs15+BH9XS7APDyW92sXjUCq8EJx7PIn48nQWa4KZ/kGE8K4A4DXVX
oXH0n6bWA1tUt071oyrzc/SQd22vkvncgCyB/F3QUP+id0wIr6LHfPa6nUxQkVb4I/TkVUkr9tsG
D3qmxEeKocbPmxvKX4XplAPhgkFs3CTvXHNgnK97ba+n+0cGNmHkNuXM9lKVqrB780ozmuhXUEMt
kAaTAUvg0tUd9vBwuCcC9tmcTJnNxeNuSNfFO+cZsZjzN3MV+AYwk4PCZHOCZ/0y6O7z2gmSMTQc
S3nkSW1IfGLLm3y7GiP7yoyPw5g2AKyOefF9UZ0aKkd1Yn7bJ04g0r1CR0bQc7ITdXsxEDyAbQdi
6OxGaJmvDB0KcJZ6VOd98GFHZW3qenqjV/uB284Wzlo0s70vbkF1P+fNJWtpfSjVpLHaeb+zv5cz
YIpFW5k1NXq2WvV+v2Jb2tvQSrptO7GV/GzfP1Xr3nfesPIdIImTldiCR3F3EpwattOUlqvr5MUN
lQ0YU7j2bD6VMYzrFpGp/LL3JZJzWxjx7w/UUItEE2uqnLTOMxrByOehDRzKQ4TMhWjPudgUB6bJ
6N/vfbquXUOsQ1vZ0W6iC2jWxjA1WHBZbnXRSMpH83Sm2QEC/rNbfLwlSLdQq6qxugJYwAcE5DFm
cnWsSEuMehxiDgrltnmkzD0Me1TSMz2clYuV0lp2sS9D9kdFZIlEQMKtoDiRpkJYH7TGsPteK9gk
/7TouKtnAO+Akg+8rfl7vpi0Rf/U4qvMxZTQlqq5kDGIajUS9APvke/cTNcKzKwKnb8KXvhaZ9sE
qmWFdepkH6JbHbbo1ON/O7gBEqt88O1RhwAA0uu6RMR9/TUqoNKmgWY9G4ZQ1QvxweH1USfb+TY2
zLQPTPT2FBnMD5GpuQw6PgwsPq/ZenQ0lCh7IhJnZSbGDcfTfS/GtiEfMzvq5Sim+M5hrWaFgce4
5QsjZ/ILBwJGCBdYdZxu4B28gJhKW6oQYBmHWbBdfCh4YtM8jay+W3jnLr3orwycgb8+zGN9fylc
Y4zOoI4XpsiyogDh2onr6FhSpg1omruhN1I0jmQVx0W79RxS3NjnmjnTdPQ7ShU12puVb69g1eCs
rorAVIs4Po2ELA3Fx1P/M1af0oiVRk/cE2ep0iWQRHCRa4FK2U8tXB8PGnIZCxqS+LrPsVcWcloe
Uguw5K4YyqKeWDt0DwhtrEPEyz86tayMna57kr46ctuiz4gMfAu+z2nnI1F4RZvoM0fL4RQ3z9/M
/HvFjctuH++N8Run1Xm5aWu1zs3M3xuu3zO1p4oDZ5usomxSaVwcH70YOEU0DI/hHU8FT2LF8Py0
Q6cJJDv9ZRK07H53v75551OSsUp9zxlohnHxIjuRIbrSe/bast9+67MvhxU3SmAIEs2AD9vhukLp
4elwBD9Lo7sbZbNLOUXuMXx9TE0a2tgQU7QVSW9iuYEZg1jXhImspaeXPLxDqvMA7/7sodazPXTq
oiqz5IOBgRziKEUi3Tow+Gs4iFYEHG2FhxnIaDaLRbJoNcV1FyiGSiKRE7mC0Oyr+6fHh53WbCV0
j3DlfwnwuExxDB/2fawFTYkZGevsWestVi7vBa+Mtuipev5JfEvnyQVhBn5e8fmOajVCHN6vdJK3
YOt7jTy6niAkPGHq/rcEPZfSQTN9vNSEFEH+xHKpe6hkKOb3UNS9AZst7j879rY1Cs69HcX/Sohd
Nj87zexWSsEPuE3+54sIcZWQZZqcLk45uUuQWjkL48D9llNz9R9y0U6IKrkHUu89foYOEUaWjuE4
p46LqGSlGI4G3qx2dmBojelsFVkaZh2CQGvDRRKUPJsYY7rXPkqBTvWjhdf/aTfnHBW3ubS79HUA
0Pkv2ZfYucQ74DKxcOJW5Z1vuzGeyPreazaPWLBr+b/ywiJi2uGg2UtQ0upZv1OuLIWbi13d+Qt4
Nj9NJJws/45jADu7xI7ouJTcI2ZJxQCw8z5aFpxuKzzdpXPIb3JbuGbau2qewXEscLdt4Ba95T+Q
Zuix0747GVvld8CHaciYOJqwS1iwZCuVqq7Llfp2yl8CEIkYAQm5I02CAvk4zUNCZciXfKaAVkFf
9+QAFB+WpBGsdYeA2EgQpS0GG1NPlOrSbD4Z9LUWj55tNh4C3e8Tck1Er38Qr9VpiOHnumBCPuH4
Bt/KGKKli3qj/I7shYhMFWhsC72d1E8lzhJlM24Rr71Y6cHdC0c+7j1kzD9UKGfAoojRb3UNcnFk
czcPUdjUuWP8IQKZEWAq6uKQS21fdwQSFnJ8ICIIDfa7yESWn1NfgKP2SMAIoRjzyGbKp6rLRUHU
tSXvGTP2rNb9UlKO3UPyVz8rMXHXjEQXsk87+DvzX68QQ74fShnrRBAdfhLIkdHj3/pn90bO7NSF
EjX205FigvhXPPPIEdw3uv1VOgTMg3TtHRk6J01y5Ic4/lik5KiB+UMKJSeg0X5j6D3zIgRKmBSH
u62ZS8xqf82m3LRaSDnsBkDjB0K2vdvypgFIPVRRlEM5owFHpmIs/ytzt2BHjbcY/RSQ8VBtKUMX
/E6V3WRBqbqIcyKp31Qlnza0D6rKLNXaTyHh2eoQQYEdwVozYbZeyWn1AbSJvSWWv08RBZGIsgBC
ZR8XqfqB9R8ZVhd9UxAhToK8zHYWLO2iU8g5/NYHjYRb5p7h/zoiupftc8VKg5NzRrP5ASCvAYTw
roETVXo1ccYm6D1b/BI3R1aTConpR1p53fpA1FHDufiyitZYwFe4MtBezTxObSKKirxF4zyX5j0f
ENcVtFSCn5ogy3RRuccROokx7YK/1bvd7jvTavPTyT416LJfUW35TsVu7grmJoBGipdVX4ObRjvy
405b1/gqZtoMvX67oFYMcgAqANpXU0I0z2/p0sW5GGN3guwt2oewByaSDhdRF1Q0P0ap/cEYqKiG
+QrPam0Be+HICvBmYl0yAwRcm+ggYvXBzzydLTSInsGFnxtOM2MsOkhvaElPSFhWE9xCYRKMoUYU
GJYkNp2l2fjFz89+zFu2SrXh7XFj1GM71UfAYmtMJz3jyTd8YljnKNB3fYBtG8ThbMJ2U+RrexuN
Qjl74azPhD6gZ6m7cFGlkIQg4y4B4zxlFl1G2+RjXiQRMjB08yL4XMbEzyk7GS5mqSZkuwnpVzz0
iF8pKFIs83Gx6ky2/HmtLtoJ0kDckep9dl0Zxc4gbfGDHyPXX+/tRhS+qwBTNxPuukig1WJcFvEa
YlI8WmX6oCb3XwWlgqK/PveYiZJ5xvhX8ebQXswcecMZDLqLWc1zWpdukgK1JlkKSsQ4Ohdwdh9N
z9qJf9ZJzYYt+VyXjPodCKESdlh1lu8LRyKGCoE5DwOjq0iRA+BBFZ/cLbY8OuBMpwVXyQPVKkT2
AJcZy9IUfx6vr+ttxYG7vH2albM9E5XCK0TpfSYvaqmXzyeDYHL28E5kaSgtp2WMo296epppCfcY
UWb5WoLQCc29KsUhwZNfa5BilWuYZpULwxiqZhBfKwLZp7NUjbtK0fr3ai7ofkeWPkvC1ZeV7+It
oO/7oo4g5c5r/i7KeIgiaqOuPcVpMvko02JhhF54Q7+dbUybPQTKqrBuoT6ifppRY24OTg0tBD/Q
Jinl0043nc3YWLb0T4TdYayssuzzAKRvFKge+3vuWwoZJnw1PLIfmZVaEZvdy9u129hVhr+o1EHv
y+WV91jZdaeJsPphyzTY6F1z6hxWFGTbTvWwY7cqlCn2AsTR8lXassD9ZWg8E2rPxZ64CHEbAqw8
UZjHTBqfoDDfbSXQeauvR3MSGWgk+vaIp8W/y8hFbqdJzdVsabQX5bSN1Fo1JOL3YPjnALz9Ak6q
v8CNdozot8cxtbmQmmVndu0t5YnnJvux8xNZxwF/e02hXlokmohaddsimVE+W1IztGasw6eC2W+5
gbqmQUw/ptI/Mz9/Efr1iO9StKNLajH4C4C8SSqPE2D/itlxWb1QCsnKyOVaI2ZKcfZR+l1Gz5EW
f3b1g6L4ETY0MLiusNAQa1Iit+MNsoaoTonSYt3L9e3OSmt0YLrp96HYYxJWusjeZn81aUZGjWDz
AIjdeJ97Mt4vEmP7/K1Yo18CaiJvq2Fe9/5M4BIkcYkoyN5/ZnzzzC+8TgYtv4Oh2LBADSMQBnJ7
Xn1Nm/uJ+2M0CCKTQCtgOuc5ZH0i3DERmHKyMbxl9ARAEYcJMW3XZAz2Ij6ww1t6B+aSzujurCm8
KBZ1P7YtA/mQZnXy2f8wev+WQFdaDsz+K12Iid2MKJSpgUfp6ysWVNXrVO0stOrUcUPins6+ii/V
6JDAo4/grlbZ9gKzJCQNO6pn5gN6j4QU+NIFS03hFB7dtqMe+8re5WL2XUwgRckQmQLEodt4ehHF
J3jzeS01ZsP2/GmTE0M3rW1/rPy0eOG0uDR+3NwaTQSOYtP7nnPKJZzXJJ/4rLlD+PPtfb/ynmej
ZmiSagIayAhcy/c7Wb7wiFOCL1iZEV4w7f75qa+HEFZBW7KgHMrJBiqLnMMlhqzmMVWGgzALpooB
uhq74DksSH7E2rD0X8gSghL40HiIWYCbIXD2PsueQiRqDln36b1HCc20A/vneNFh/fS5RwE/Zp3n
d2Fl5tPE+8Otvf29e5spj303aJ/CwAWDzJIIrNfZ7o+WlT9iEeWWomiFKAIhNUCQp3dgY+C8ufTy
InhvktQVX7DQvNXS6gAxGKlaIi06YfRyArOlVjjgXZ+waVU5KHC57pYpkuumTtgw/7li3DouhZUY
UPWM+tpUzbiPC5UyHni0msBqAASNBbh+ScfNqs5VKQWfYdW6/PcuryDbALxUR+QGZfCo42fz0bDv
Pb3QJIJxVRYnVOOEYFJXLnNHgMG0f6n3bHzSuECv3UPCKZHF4wzJ+ByNLahIMJmRGlsU3kB19hv4
798MdNQm/jQbLfbqGVqkSIQTveRBS2ZJQZdSMCxXWYi1G4AOH9MSdxRlwMdpU0nP6URMnoDGZiKi
zx2BUZWtGxOgVJTK8qhlHJhUX4gBDRNgCiM/KcGIVXY9Jv9Q2RZsg5k6lK66BoELgImvzZzSOzT9
ZAf6oJu1YfNVOSGv2OVQcUDosz05jH1yp+Vai5Z0YXexdwqXjDKle53hyYGz2WnZlB/Sj1BB1ABe
k/EPFv2WPL7hzUCEZpgbiHV48/hqq+m1B6iQU02mqP4765e0m7NdXOi0cLO3/3vTcoN3iUi5dPkj
9BEwdMEosoYfTT277lEGKSZcu59QBp/jfYN0AGXZEGnpg2x3JneeGDVdtW9Ra8NPlK06v0XbFNeq
rzveSVCBdFhZeGaeTc+NbuesefWnPxbh9p01UoNfwJggzGotbdiBYRbfslZGVuXfAzAQmmEGDDfT
abA3UOIGgG5HHCEsnjkYWFv5yhvXd8kYTsCKtBM2qQu1+6WLj+HI/9gtSFWwSXwqp/ySnizxBB7N
LTNXY+ND2BlIc7E57exSS30sdghcJ3vRz1ubzy56RdGheMO0gRwWV508zBJkSQLnCqNrJnLzSsa4
3qHYHB4/oDK+N7KsYe5e7JRio8AyD5scdX6NMG+jCx0FfYL6OMKJl4RoH+JHsI+G4h4ZKoXe5d5z
cxQxK+99D2zeRjLknsl87JPrgLCJW/x562vHDZsP9enGVq1qKVo6rsUzLrUCes9JRFHCg0L+ETzx
d2Q9ecgHzpKnoIWX7iMsRyOk9aV3D4yXmNW5uMNT8OESQLyX7QUNFLWfy2djMP1pdJCBXGqYMLFL
nQvgfR4MKxgM7SatEjiZLY4nX3NMPD1jMk5t/LJfa7NK0c1m5LBmIFm5jpVftnKTiv8IuClkHj48
lytEpWHfulkdCsNHncVWn6p5OtXweqhTUQ6CWYT8F4X18nfDJuSXZn5THOuiXWSb8hKKi1mUenUy
cRm72OWWWMlBJi4ZtD+WlOOTC7TtyEKeXGvZvidZqCCHOAvGmSOdUDI0qohgWm89yLhWApx8nv3a
e++8paaiGeXr08nRBxd6kPTtvZOc6F7tJvfRoFvRh1kzcb+teMuWPZDZXbOn1Tuz2opPwKdnP4Ez
GttFMJPr3whoMQT606/oQOiZjUjT4AvixFFxW4h3gSzDCMg6PWl3YCZExE8TS9Qu2kRPhkl6PXB6
4Vpq8VxvDX5lc5zHU854S9r1TWSXNMAbtMkF8cUFqhr01fDsBodh858R9+LNuP7rWXQH4C9yOxkN
cHGpk0i+k1ImMHvcQKzwXWWjbKjGGbgMJHW8dpFx94PqCbC8KV/KL9LLxGOd7ihKxT5gaQ1TAZsv
jB+Ju98qew7v+0J5HEE9Y173t2+KD8xZ3up/xj1ExsNa81gfnQfVLBGFeCY+VXTIOpXoAdHNnZCu
bSSXKNqIBeE3nMjmVxgPUqSAs7SnMWtlnnU7ifz5kN/l4a/7rXy2APLy5a+rt+tbWXbsYdt8KXvi
46p5/0GCnSl7b7qGE8o4IVxwUTwO7k5XWlGh3Mri6nLi3yMd0HeYnq643ObYnKnqh5sW5AAQe/2E
SMzHR7LfRMZgOZese2kQ2Sf1Xuf2bpSNVTZbIu92hPRif/0YHV1etQVCZva1QRSBSSYO8S66Mw0+
aXzp4ELUtMkKB1eEiNBid/J2bwm+OA+ZS4jZROMWScmlYrJyr9URapSm7+1Rr41spo9xOG6GcymS
RZRNvJvIGVrsPLllxPItTkn0AKPA8CBVOoNQM/R6ktRk4Xe3eal41rAkYnljLxMOCSlsmPRwzFgF
W2Vc1SpZHaHXUpmrmoZkM6x+AKwYasXnE/ibXQOiGykXAYec8MnuVGCVuhuZQWMvbaM19Q4vJqLN
qXjC+PmcSktPL9iLz4D5GDqsQXTPOuOpu4+eMsxfooRISRXvPviEzuxXHOA2Ejr/oJC3zoA5k+IU
Dkh/z4rCcvmxQr7GFPHDW+kSI9bhADnVjYRJWbrWgwMOvPqGklrq0+6cpARvW6S6mWnhStr3OFia
EfsdjnvXIMzvEAn1+TBMMJ4ihGMs86bgYFheKVwvUj+vvK2ZLOj6C1vPNH8EwCfUFLT2+7CRl8bi
0Q+OBYNn0s0i579zE9E8pQsUovv+0ByQd2zuwzDzfpd5BgEDWlcK36joroI9aXNyXaJe2z3sFt22
i2yI7J5ui/PZOIDSoW1UPOymtjYj77Qngalt1+QzosehcqnttcKz0EQ4H2AJDdusHYzeBqHIlvl3
Tx6y6sF911j6HVdZ6z5avy9cgJ2+Lih4hC+WoAmHAUq58oI9L9l2yLHHzf6tur9jIQbUZB5UDiWK
CO0cA1CIUlOrEJePpUkl0odDzZeWI1/XbC5SDONBc/IiuxaU/XtebSOS8d6P6tpLfVg4yb4GE68D
lj8qDpxBC0oMlbNTT3QUBFQHqPtE2iqPW9ELjm+DZflbOelvUSZFhzKFDAsYpoDp89FFIoySEhvy
XATYMHKgeGCTJAz5N1B/j8VFFyBdcid7xXDp8MQaZd9dIpTgEkjHcUU2X9HvwybF5iu/isqLEjON
W8R7YPM9rCl9SvQSDLk9kuW1XiaSMlSwqEu+Qy9/4tPqYdrHXAq3/ZxPB7+lM3N8OQydVEbcNapn
veAfFvOlB643quDgF2liujaSpJgKVDbHD0ref5EKsAwE8/kHl4QXI/Frlkgp091nk9FI0yyeGg2u
H0xd9SEW8WBZUfecFfdYeaVu9gPsCpZwvMeY66faJuQo862EVgZ4psa5vrY44f2AHPd1i5YBJHK7
qaOvSmJ19jZlnMvKXFStsUlPNxFTfEHJ0n2QGFlp4s9mQpjw65MBFcIM1xLZL2VfuZTyrWmhk4O8
xJ32Cw3oU91s77l+B+GIjLTqmZpozx4i10P5OpMB9kXKmYiMIxNdv/c55WUOG6ol/f9to0hpBjI5
KuS/5sGVHZtfDVQbqjP/xK0nKP4+UoaRXt5zdN30LY2nK7U4YZlLsTwQPLVcr/ZuIaGaJxmAVuyl
2mvpCiUzFAS4z1WqK8AvrTcUNLOA0Q2sDRQ1/47SXBgG2EMAu5MjjQI6DcD/K+B9W2F33lx6LffS
Tk9SpFISNUDcCsk2WLK1XaqbO4JWXVB6CIiE8BtZYGTVf/ZeQvtpQGzBCYZSZ5LLCH9bZop9WUE6
LwbBTqkZMoU3oSUBe6osh5t0lkPGajQjNv97x/qQsgo/+c4oS+0nPgnCJz12rxmFuIURkAQNazvL
BZKnF4LKh/UKxMTAbSy6T+Houm7pcVIrBV76fCe/9p8aBRZd1s725bOicTxPG7vZxtG8bTXldqAP
j/Qg+8W6Zqgyygiif2KzovQFsieMS0LbohpqXTGn9hVXR4mHEOSrAtszKRIMEzjxA3Ne44QwWxgS
oidw6ki9G9B3qqM2y5Fj5YPCQZhxmYeUXNjeP5chv90uAu2bcxq9D9ol+pPZDqEFuALAykdXEt8U
iPpNkeLc9RFLnedhKZX8BOcqInKEQ7RJC8RM/ztSryDkvNMPAfxi2RtR0h7xuCIyMjQG2i6e9GLp
6AH6FvmVLOhpkiwqxGX1NqZ/pAQmiEY8WjfjHj8O9IFTtv6+3DTaabEKwJpQEEPMds1oVmRMtMRO
/54YUaxssp4Et6iogk4ymq84/0cH0brNbz5gKaLNH/JJjEQVFNzBgYyZ9Wdf+6DQtrCRgDd3jb1/
nvCkpstNANi8KoXL4iA+MiL8c1gO8pknOGQVA/LF23CMt9jWpX4PNFh4auyXfbvoPh38575Y/E4p
1JNSkjmvNF42tYuPvNGH2iEemNhIXScNQ3B1ecHVmDf3bt/gOh3Uim5lAYUn+XTT37w2btG/ero5
oyTTLRuWpnUGeTaaNNmP9dSXhY1elFVbrqVvMhxq/2gC8MFy6V0RRQUlZyTjc9PWea3/79sgDRpi
X0zRD/4FUR3AumK/Ccn0OQ2xdE6jEVWUqNY6qtYeknDNCT0PCoTztzmjoRqTmaLQfr7ocEzUhFDv
o72QXEZ5VcpPnTi5uGJxhjfOzRvW+W2xvj7ItlZyVMXKmfIFBZe62NJBKUTd0TTRS0+Gz9NqpeSh
SJpOE2uM9ErXulnBHQVlMAbgYPKtp8cLlFt0tcSNqE2AnryI8s2MFch3OIMPlWa49M2AjkeRmUHH
i95toMkapFF7LuzYkPJZmkWqi7AoM80//LX5qNZPfJpG+m9hpLPkycTbbzjGuDj9szBZhrre2ziN
nG/QL2a7FDLANoHbynKe4T/Z/Xk3imfgiT6tU13ofhw5WWvXl6c4z1aaT751NiGngqS1WYGEjFcQ
J8f34g9DzumHyfPRcB673E/q+ZniFqZQLd6Nb48PX1t9p1xjQbmwk5Czo6GgXfAWQ6wzHW5AXI02
gPRyasB7gRV/cxBHUQBpJQqyT34Qd2Vr76ZpXjDdolkNS9F1th0nQg4/S5mZ85ExPiYEeMzdMa34
onzVtyVpLGq1f+9w4pWXybaWN0aZFOklXo968zJ/5kwm4PL8CvSjah3A0OtcgHNU1S5h6SepbYf/
DumBRavUpLDWmuYkuWJgZp+vn1zgTXrrTMmWbTo90FzpEkMJzE6MBdeN9i64awWfp3npOtJx88aO
lWkpX7pFyV/uMaRS+A/D9BSl51UedesK3BD9uykPH8MbXu2+UJckcTsTzYafej0Vlo+NzTNWOApI
Yxp+Bdu6h79Izgvqdn5lbp5HQ09G2Gm8M2lP5rbFdqtg9jwlPJ+FTvO3ZxHeLKfF7tlsB/Gmyb88
PCjsx9kq8Z0dCZi8h19/BnqQOLtfY3ivsXfA+fcplmtPQoRpkVY13L9I1Qr/nwXkfi0/Ye8i1DxB
BRcWkOKcFgwhV3ANt5k6Nwsclzw2k1HLcmY4MmEdjeX0YlfCTXTQMAy9K9kskWnR+Q/t8IDc9Zpm
3uDB7jB8dv1XfwQuZQAn7/qFPbTWvpE1NA57Zg3sboCPIHjR6dnl1oDUDOpvUnaMeMTov2H+LoGw
WdDM5okW7k8LTKOQPQ9FFDTpLf1o3cvV9aLDPfOU0dAzEu7G+mblfF+lLhKXg1+Yb6VmGRdWDv/u
IckfuT6ul3EGoGHBuA51eUlpeGf+qTn3DPJuiqUwZFlvH3KhM2+hP2bxxA9dJA3An5SVUnWwaN3Y
G0AbfRoIo71DoAqhUH9JVb9k9EgG2smEYu2g+j8J1B/T0TOvtOmpGdvieW9PegBFuRdAmi+QS38/
fc5sRoEGI+QFuLCSp3qDQgOIUy8ephA0v6H/JCUP26a2cOT/0TBe4MIwmgrYZUO0tiRRta5FXqpK
zIxcWO2NWswLml7mJBKvD8Zk6jWfMfmhdUivmfpT+dS+jvHAy7oRgQ4SACrCJbzXGpVXRGZnpZW8
WfDdKgdY4YyQXO47h9fF9dkN8R4WiWZZusDoYVFnjkve1QF265vKsGSEyAGuzdIuc78HsX04dazN
UKG0Sk7n/5r3tf6v/FGPgFLg3vou5aijutkx5gpFHVNhNgMhlz8jKfmsOIk55VYRwoz16/P6W8zZ
YX9ot1cmiHIXqVlmHMmdkNdcXsGNKZyPbi6B17v8rJZBb+T7/QkBQqHJT2PSXxgVU+Eiu3cj83sx
VTVWOCbgiQ5lIJMqfhszn70diBs1VNQL07s7TOrgxfvfSNkuVWkaU+PyJmGtaHD/NeC66p46YGV2
/rVIJb4741s2Y8jGZTNj4IN+m6SpfpqbkzlTx1MrXEVht3HDe1h34IkIt83paucJUSxPzJ/ZYeLs
tL0n2X3asiZ98FuYvvF7Xlq9l3erL7QS59f7mim3Rf3F4WaiOozxPaHveN6e4Nsj0nfHvh0pT4gb
dW4/150tLEhniOf+ghqNvcKu1u1zCUSfwm/RwkAyudaRl8HRyVq9J5GtMmfbHVFfNJZ+KYmFomI7
BtnJFuWE1vsbE/+LY3SBXTznd+QTQPHS19GQc87pXay7up1c08g2szoGikzh7yqaOo7BcSGrN0rG
VWcn5+WwRAVYoMDRdwpAP5PdkP+D8bsZglr1wZBgxR51CUbU1I4l3miRsRg8ZvIBUTnz+b6WJ26N
PnS3D8rBmIWbqp6DKsyqmy7Grj+oK/jVIDhI7yBjE9dE6vNCPC0aIU1O10O8yXQnmxVvrTWUqHOi
YxKlEIg/Z7WleiAhU4Eq2jIV2h7uWsBUOZQ+vytGXCfY2jVqRx3XmX5HO5wVqU4T15lG3nI+tl3n
3a3tLscPT1CZMy+Ms9l6Czsjj7McHOj93TNxr5BF0W66aBx8cezR2uQXyuVlcQ0AqMmOtY36WevQ
L8u9zl0cSCmPEi1uzv9WVbg47aqA+TVcQN40/iRHQHjziaTTRyJxpAdJ8cEe9hlETORBceWdSZOP
ZK7Z5DJke3Ysh4Wf1ybOiFLToD88WxEk/gpmwXkn5fGGpQKoLkojXjATesstzDX4+TyHXug8/dXm
z+v5tpuBoeDv4TH7J8tFsrzsNHMn4lZYQuVyOzgKduonkUfoIghXQgkMPetPZmpoz7SzJCLhBXlj
6gB5q393cjFH/hw2Ct1UYOOr69ioOzSVFSgVYbJZ7Wa0mtHdpKJTt1x2INGQnPJYj4bvGuKEXSin
NJzgLBg/rqVmfYJ4mS9tBst7+3pYNhiK4N1qaPEK0FsTeyaTNLdeaxVxTSmOuHG7rICof+3c4la3
+Fkakh2+3EKNHTsDz1A3x3N2lEr66SKmF67QueDnE62PJEQKI7WSbMdaDYm2LN8K1ZnFJnk9iVEn
W0piXMFGB+6DRCzOWCKHFrH1d89qxihKYhMsHhBYnobUVyb5V27JGja1gypw7ntUEXK6DWC+Ps57
VyDBBdDIdIuo2d3mILiiSS+Xt3NX9oDCp68qOlqY3f1TcpIfe+w5JjplbjhV2VxyBWgjqNgrCwvr
xSqkf5HsD1dP+TQOBsEJ2zSYdGx33wtZQJ/KOP4+sXfTxTggGACOByAHdFgbg9jjJVfEV2F21OGO
MiYVeklIS+6cQ8RtW3yUHBsSyzthbU/QnIKky3LWfrqlvjHGpBwKyvfsBPCWukWxZxLx+2JoO+bd
fdDxbA9rXml7IDU9bpMnsSrAzrGWifmAhpprSFxRCJq60HxG9Sa7FU99z0DwApcmB3h8HlcuCtiO
sRM4v2dfTWSD6HuL1aKdIy7LwLwDgDfebxrVmzQh/Ym3/E4yP+kdNbeNfwbr3so8JQ5sY2vnJxMM
HksFBfdTaROg/pJ7O8tI6xmC8MNvn7D8geQYeu+6rFT+8JtysxPsvzP16/3ym/9XMVSCvIckheXR
Py1fIC07Riah4Zl3DFLJATf5R61C5FAihXuxOi1cRTomy/U67yM3lcRwb/gVAnT9D0l39wMMX9p6
rIFBFJM1jyry3tDLfNEEEPKdv9C3xI4SA+uwodmR6IXAih0vWriiG9VQE6XZslOCtlBxGJ3kZI/2
PQwh5om8/Hy7FFkDdX9asE5u58PypWLrnpB+DmoCeIljzfFIxu3x7/AHj/j2aM/5HaZgIMc4HDMM
xTl4yzH64xnQ1PpfROaqXl4PEoToV9QMwANJWMSA+Hrakeoi+Mrhoqi7KZ8JPDkedgEuL/dlZ5lZ
UQT5yz8N+9NmDF4MUuVfs3QMfT4/w+40UnSVRJSF7F1+/2+ngTIl4ojYyqzZVyScrpa+xW/C7KQj
TDguDLfkb5FyKp28W4gzXRG02hLdyhnYoVdMSgCaELM+7TMTGzXTQXO0+xCjtIx5gSM5UjFjOGEz
Fx9hwtODgAhQ9pRlHzhbebsNN6PiuBnhXF8D/2CY09/R27YuoO2LdiwbhIr7MpEFW9dbs7cty3Rd
lfwhzpgPABkkBBP+p7P6dKoZVpskIMdtUxnyMOwShC+bixO3854gP7hOj3m8vcdSqFtPOfAdBF5O
hBLE/Rg+ut8zOV7ImxMSXlPA5LWlQ8VVFQh/YX8mr7YnLC0tG0ysx9+QShdigePISkFkgCs5pA2h
LWZDLGDxu49JuoICDZzBj1nxyc9oLq45Ijp6z8IK/hMLR1+RGDSaDX1RQ04Nw8pfwm3nPpyOdMpa
5GbwG8/Cy2+eVVMs/PDPL4PdI62uVV1yDV/7kNGTnvfElv0T4PbJEIYqnxB0j3Ik9ljxwy+jAm0a
JwmhTrDaoceA4DKb9Vui0lAkvsCPcoPcETXxC03besgYxYotnmga2eaOWNPEF0HHeH6S8exx//td
qWbdjrSBVoo1d4iH5pKrKEqb9vd6T4FsANNEvPBfqAA87MUgtyAn9z25/sgdLP0fsSscDBwYCI3a
0PQacqOsOwHhlMoyIbWsqEmS5U1LccZTJ7FYI8nEn2Gox4kKjiyRZMgj5IopPHmKSWRdH7qdYprc
9hVeUhqYTm80zUM0L2PuSLNx2Blt5rHtYiCYCQQQexG44BlI2VoerjKhD+PZEr7ax2WAP81PbBA3
N+N4gmuHhMiH/cvZ7iAoCyXcDW5UsPcoS/uGhFPeMX2uio5luNiECITwUzoc5kV4qrTdgBBJ1+Sl
AQu2C/xjNl8UHBFkmxUNpgLa8vcvbvR0v7A7huFns51lgwsaG2EcfLCfNi2oFb0r+8hchp+r2hcm
vbp7n/J6FQdWvR56Tn9CP1/lPkG6OaFchoMlq24ug6grTfH1HxvY6ZRrC1ZIL3/0OHw2XhIYPmWL
Txdro3eeTNEs5fyYLQIsysHKXbs+SBmRKggbWJGmS31sXjYl8q1Ckr4h+0kgAORWChJooHCEoOk9
/Wf0uksZNmsOunj9/o9CXVq/ISqmHtQ3q6O68700nBjAvJnk9lUdRdR8R6iL3r5DoAgXKMH/SMfB
CHVcPNcXOqe8I8cEhwLX/0Gsv5UVjwDpGEOtJWxoM8DkENjAe6QoYo8jaBuE14Ba3oadKmT9cIzO
gp6nF2cTcTJ1HCTgcZhNGeYHzGBxkwPU3xqc+o+6DMnTiQIE9fgoXWRnvMsN2M7G/jLkrwJ0aHbw
LyCo90RZTlAk1uehckoDwO/2Ou/8sCYkRYelL6w8LKI+S3Pgfa5w21n3CqaQUVjsea4nc1QF93Xj
LFZnKfVUBLn7yrichuWRSoIjTywBNvBxB3yBmT7Fo1OKhgYW3E2Cp5WqNDWHbjtVdc0Atu+l30mg
6opcye0k8grhQXGxyTG3OubF4jmBGTVdSxQb0HxGM7kRliLf3MycpUaJyVPqOa2ImVzLXlWYOOmH
ju6bE5lJjc62O0DYZLoaLlBfSwWOPGM2KMYX+pkBY+NHwvhKZg+/qT2kWY8IJDtWe56XSx3Qs2hL
UjpIvvvJBK1Ad2hINyvQY8jZTCC60NMg3aQ8PkwdwA3fewCNm8NNnFGgOPsix9ntH6Rlt3IqJ8Tl
GnZEU6P4AmWQxYektWoUsXr/yV7Uod/LW/BuqTiHd1fEx+QsZd3jdgTeaq5Wer/wNJoycTNRUBhb
pAq2aP1j4bWXtUhhaTxi2fDNqUh05LhrAWmTF6KdNtC6w2Fw4a4+ZGHU0WAM1Sj1T7F+4Rpu9F8E
YFUnk9cJKLANY+5dSW667A8BnMZDP6zFvi7tCBLxTMq3HNOR5dEWtAZxKJzr8XlWDMTWh3KH1qAO
5zwFJSKPSOkLVg0iKcW3leF2b+ABDBjNqh21LgV4bsSJ2+zOfkIbZkXKsc3MjB6icfB6hTbn5otp
smasoNojwOj7+z1i44Ll0BPafUNUUHcrJ3MK4FV1aSJOd9CmNqKjbV11zNGbMTeTWzqxtO/4E2f7
8UatOJK5fqN/UXq3v4plhbJlMWQyzV066oheMQ015Zry4Js9qwmmsAoTKoLQfrSIIIvBsHLfLoE8
M8tYVzxjzuGrrufVFgQ4+/kWoHpYoMctq8z2Oj0+BoKXLzX4dXaF2Myj9L24klOIlRGC3tHOV8hm
CnjTlkNNpprOrWoR7zK84hwk+0IRaXWQqlY0UFcKtBYd/jsb6nKehLvoVey7Jx7GxW7ehM5Bverw
RERKI7EuFdcAWPYcrJ+k2Q3t73mrpDpnygx0VzyXdcTuryMnnj7aYOYwjV+27FiWnEPoklRuyKvT
ze/On6H+DTqNd6OuyApemh1VeXYmpMYxbLFPOchSDKm8NkhDnwwu4+rPgK5C8KL3Gd+O25Kl44ku
LQe01izKe860OnD1WZM3tau9on9IGX0emEE4VlqlOWTyXMfMYYeeOGMx0UQbupfrrcXlRUIhYqvw
EiDMr5ncsBX+o1A/ebraLV14akxMiD5Vq6LKdqBsAhyY4fZpxomYNTj/I9zjFBaZYje16Brf/32r
vGRNbSlre8Z/mx3AovaNr1IksDPeNVDNeFzo9QGtnoJsmBL3IAZ1bWlmBv4S1lYu7i+XQyrlRauV
tjLOoSJBz8plwvjQpPOp2dXQOqbLMdpyKFBI4+W7g52D4jYaeM7LC4xPBJtaFo5uH6pLguSp96lS
+qlfG0kLuYEF+vgpiPnyxr+x1x9d7cuiOW/KbWgQyvsKB7rWYsVrPybM4ICV8GV//L1vZsRdQzoZ
7qWKC12eZAIrDEsbqrF4ZVdsMGpkaIa8qKgCaGwswJdOwWhTWacyF9Eg5BBagf0hAnN22Ilz9Z8O
eWDiLBaB2W712aXtM1DMi/mKqh31buR05gxMaUxj2jsqxJVIwlvevfZAk49RDhI3L2AEMRWX2jlL
OB2MPAR2PUV+OrU/X30JhbrUF/cmV5mWZe2rmcpJLkq5BE61/8RLCnGPGLfLNyk7VnF3S6Xx2Xbv
VUidmFjCiotFk230V0wDGxrmwVWgqUKJI/SQ5IMBhF7LzlYkw8ZKuRvShgGJQOytV8jg4na1h+W4
BlvSdRqR6by0YMMOF2LolnxhjZU7O3a0Tn9AuEIFZiF/22WTE1SNUrlxnbBL03CctPWq+tBht5ao
/abEc66i0SdGKt28MeZ/DuJSV/pvyor9zODeFuSWkY8+cpBaK7NsLyrjCTpWvVWhZPLMx6P9O2Ze
h1HX+YcRzc0T8nulYUg72wgcQ/+hZkPL4U12taHduwo50TeqqPLTVsNDd9G6AcUViqCqqB0bWLcJ
BwyWO97lF4pfFpHVF/HN2I0c9eEXwo8evEOqnzGljPb5VyG54xG2AvGc0Shpo0zbySWtrGqJ6mmw
bQvcag2lFi5+Sv6mmX0FYkjkPM3nbjB4RVJO+2qFozGhyEXkZ6BkbdOCEw+LWjcybmoa9TR67dir
8n3uBt6dNdU2Zzi4S85WAzkOf08yS8BGMz3YwiknnNdVslZfqp1JO6vOJJCg7FjJ34VnrfHBo31X
zR3ZCoPjU0Lk5sUlpgph9VVEAuVu4OM0xrBN0NPuHLklG8KfI8XcArX2WToWaGZCIup2mSGstLh0
YAzxs4hCKBMMMs9ltAjDrL5QMGUgICH1m6oBCqTBepUv++nr+p0gtrEg0Fg39eldqTlPoQFlgf4e
UIQxEj9yIqhuVt+Ic4OegHV0bKBzmyD9kziQ1iZRn6gLQyZkVrW65q8LVltoAX9ZuDShSnXCP2xA
j9ItC+jomeCwibC3f31dck8i32WnhIeowBFoXseyTWutbbmmiBmuTJVYmGrhnHwH+eC+5VO3G+Jq
9FTmc00wViWt7NxEccqdpgeM28YyacwwVzkgFr/5P9LppCMTTBQzc6FsyQEZatnk2S+6Hslx0mu5
vhrR5QbCQwhsrHHxGKFFauC/s/EjhFSP/znj8iGmGCQSZsSW6OmQsSyHWv97EYrQjxEU7eZSZ/hH
heAf8T9Lg1fo4eHlJDyFkYTzq6KLgHXc6tHBcDx8Y8Crsv8NEzKeZCYqHQXaPCKU4/T7bk8nssZ+
DdKQmgKh/KDb1iBmvpAY4mduCR6BEYXBmJlR6UHP/Xrl3f80BlZegEbtwfYWNYtkwz+XW4p61pDT
CKEtWZLbSRm4Dy35jGFGPcb7mJtB/WzDVTWeFsIZfzUWlfeyYTe0J7/GJkvzzhKDC3z9EdNR97ct
3CL74NUkrZbDmQN8pKgkynevoYY2f6+oyFNqJmI3KuqnvHLfr9Gi40Mr+Ehzd4uRMc2MFcnfkxU5
59mmuTXiUVuz36GA7rmoMqNIxQxN/jhwLOIs0/1upzmUF2AOCM+Gs8TfgJbePoR8ZHQ505/mxRnK
Eqdz/6HqXHc2N7N9Vn4ojYjLDZZ8CGIzcZ/7nywQrsACrYwCUNLjqoQi1KWD5MApU7n1xUhSM/ib
CkyMkOejR48u/Nulyzpj7Rjqt3iNZn2ci2hwsEXwdMJ6rD0l1KyvGzZl4ClGdCkkEWAO2lB21t3i
UvRl06QtzJnBjrpS7+AUIgfPIrMuPt2DVsFEqvF7pNf+0KXbpKrqQTf4yRzC3JjP3QVsc8VrjcX1
KHR4rfOhlzOax/jLeLHxvfvY4ABk6DDy86JFjudnM7SP9hFaxpQ3dTvAAaX5T3FaTXBYWs5F4YuC
scBGg9NUeP+XNgJkz6xurG7F8mnEsif27MbMxMPlzRd4sTCGWmWtgp7gOC40bP6qVRgvuuthqod1
EN/XiIQItlJpDur2wghWkxSLXeGAajjWG0L3j/ZAeNBwHBaSM11uLccDDDmD74+9evpTnDl0HHgT
EhuJJ05/yR3JIHc+vXFOvsJJueoPUn/H4KpSxFRhrrS8RnZeQhgzQBZMIukoMUqwsQ3qJe3zEyLx
YbJKsuQwBKbj9hL3LaSV9KFyJ1TAfYfuAIQAQoSXd9BF/ni2nRmrxAC2EZrg7woZGhMo1ptbRGu6
y30CrhxGSe7eHRC1FmwEyXE+zUDXLZ3pysUL5i85CmXRmwF4Y3bGCbjRq0+PsApyUOAlyU2JfngI
Hp+QpXaTVNTGIPYklzX1HIcqgT6J+XbZyNYNVsYZeCxqX9R/E9aAsPEUN4/2OXP1AUoaVB7yM2Xl
Wd08zbmKgtPUdkqYUlfDCZ77fXH6J97HUQLGj1D03bvxk50TwyASOszG7XvgwCAPDz5qSLL2yM9/
rW9HRgr/gy951t4yIZvG5Yw04wYIPAcmsFcUiumW6A5FgL4DUWn/McH+CH4l39Rd1YtHJYN9SdnJ
OacouciEx14zPxRIDDJN/1CD4X7qxIoqR6ZSYng/aLknp4RXqpoKW6dM4dLbiGpwT66whcks7qVP
CvQ4XyQ8J+d0CCA6+kDuVgZ94nw+Bg9WbZUUz/0gFDT7/ZCpnLP2ZkbW0C66fGpnlZ9NJtg0UyMe
TEEyHptuLLauR7e0/1hgr8wtDkjbLD5TTXy0WzTfvMjJiba2hvNIVRMuReFrJtZ+6ktjx185wdFc
MWFMAx1G6Wm3FPv2g4/UNvQrZ0vMTDYwExPbtrvAdKvemMX4O7ec7NOl1GQZLcsgPr8xMunofNL1
nkz7prKqxpdLereKC+XPtShVC1sjjlvfc7rw2OMvrF4X6JZM4m5OqEk7evNmtR9RYGjfzHqf1a7v
mc0NfcshpdK/ft3F1np1BIKrC69lM1OJiW1Q38V9C4BjPTNyWLctbqg8DTFZ644yeJhUxermkic0
l4ZtWm5l+HOJHwpXfZs7KXzk2L66uXocNHIF0sgYxyb2bF6B5G8nZ14qW/c4m06IH7CjuX+5rG2e
nYud7QC9vY4DdtFwfRHY1aal+36qkVvDdIFFMCVJD13lBf+vuX5ahrRxV1tAbMa7tTNCtXzgZQTs
P/+PbArihklDTsP9w5Nt/MEkx5YE7F0P41sPzHL3Allul0s3tf5awyVPkL6eTw9xa+vwdMYCsnKI
rKiJQ5trD3T3ZBIhErc462jnxKHZXEOe+cPz4VGrWYgP5nRNBEm7yoqMW1IWNpw3Vqdq590S25qG
Zk4Q2Gikb/+KLMgba1iqied1qPe7DkMLl/FWA4Tf+70CyB0vZ7Y2sgwN59Nao0MWdqL2gtUkMEQ1
pAqIM22XhDlNBsjN/NtCx/B/hHkq45fEGdl14vqZv+gqcH0M7ndYz4CC2m+jJNBkNJTbyC5Zfayv
NAeGDaoVZf23EUWLVjGbZboNZQBCTHe3fhu4ZvkYW3OXO7tMj1nI+J6A5ZpQkYPZmpJQpWJpSyPM
OfPrihDBtuTwM5+KUZop+q84LmbJnx/lzyKnzJqjHJJyLUK0S3t1y7fXOusl2sOaVGRFbZ8hHRb5
KgPzPZ+o3mRig9R8o80THXe5nkzLWOW46A2hQsZPXtETZWhhSwva8/MVBYnewdu2Q+sqhYa9di9t
yVzQft/sturG4aIvbGTwxabNlfYT5YWQMuDYM9KLba9OJ2eyBM8eCvdaI4XoYwSoTknniwzOY+wC
t+ls62FnIWiEK0ChsHeU7rKsDJdOLaMzmlQwju5VjnS/Ktsjd6cm36/GDJKV06MrNfcLW70fZrU7
3ZzXynEwSk813tlyj1oTxUfBFQR8kCW/+HlIuPOXl5XFvUN/3oz/CNboNK57v6Qj3SXyMxUgAZhU
zUi5iY2jfrRRl9Wlx2UyYY+ZsdGmcwOK47kRmhZfXfIQ2PIa6+P4CNxt8ejyWYvMwzd/pvtI1wjD
7puW/Nq7avK/mXeDrKJjN0XapD9qwqJFE74sGZkeuWkm2DBDyfZphH9VZlRlDX4j3xGsASLcZrqh
x0+8q9R2RPn2laSmPdTyJH/0or5iEdPO8M2vT9tM3Ruquw96GL1E0U3ZeMnwSBSSyyHVU0AuSW3H
XJyZwSU1EmvuzezknRGU9DjHd4e2NRWQKr0aG/tiZULTzzqgdBQ2rjITOkQyzPaNTya9wno6U/gH
E4QNnugvKJ4f0CtKDvea/nS8NQZQRKER2s9Ql5kjX93/UkPH0C8Cs9B1kP9ZpGLIfe/7xDCNxn0v
Kq+N1mzIs+KQ2g0WIa31Ac1bzHopFk0XANi4poedzgAcyOox1j/MuzRDMhATSXbOnP3cABu2f3Xj
zMHZbFQgHKtXqALsqktXI+HdLv+Rz8y74BA+leHnxFlSXHdemjQJlIZJMDQjGZ4mpLk7vh/Jt9fA
f15cjKgSZCzryqJQNtesDZtNeJedcOdMVLzV6cFHC2oKBmF27/ey235OBYbhbxxNY19PrOcXT2kg
iih/uas3xW0c5Y5rjmJ4gxl6uvdHByaj8qAOd0YwYx/CPMfv1ihaK2SgCTAXjAqekE109RHDNXPi
ZZ15cIqtgjxR5Vl01KWU3Q40oq9XjRX5YRaL4cct8M2K67tGfcDk2pTTYa68mZIor8fWA+Rn+aNN
ebxKWTEIgS9c5SpMoSfdaDPUHetmGN/59VA6k4zAR+qYma7teSNwx8xrPsGfn1aTGb02c6FLa87u
6WjSno62+AKOul/jenfjg+C9KOHWNmmc/TOQNNfwj+GUypEs8+yeH7UcaGpiwqVHWKsCutS5qMWm
LxiNMBVduvvXlC7zM3Y4Bcp7RD23PiseivuYIJvO5pDCuNM4pmS2ezvJNxSZwEjeSGNDvWE2o1Mg
M275oL9PBTiF8YtXdtRgonnstzn9s3SKw1sp83Ssi9JqZhdfD40mEtgHTWPlRea1FWQHuY5bKjIA
yIYIBBBblkN7IaDP+hN5Dm60Tz+IFE12EiUCzXEcNhIAqNTCcwaCefZTYsAnhjp3jzf/olq0QPBx
8Lrc5vNxlPu0/Xt2y8SPJSX8QpfgulVQ4TVCs2W4yUlkd0JS7FcVLfV1ftMxtkb0WADdDXRFJhS1
YCiDEbdYJ17vVqpL+pq6hWsBAPXH+mGy/0Ssgdjlcu+teEn7y1R2I3CLJjDqaRMg8jj/5O6upoI/
LMBtxRlcSfvqmbRi1LIVe4FWd4gA8H7hyro3NLrHYh0KpMCb8XI3jqPriJNl/JmSAJ8eTZLJc3m5
zI6a+Qb+pmVhEH5TlNdWZULY4hT0/2hT1cmuHncG1c9lHeGCkir+k/kDAcYIVIBwwobaBuWqTnYq
bRMNo2fWMlnS1UFWmAgLwOUTBZVPml+g6dfESUK4jIJkJNWrVaILJk3ZMywx5k3FTxteNa7ZdKcT
f0b5bDPfm1LsAFPvjJzyP8DZ8J6DdKz5iAPYUIbMhn+A9GzPcONmC2D7aQJeBBWoyAEwTCA4uLJC
bcFJESujaXA5MezYQyPzmbDVaXMPKfIxt4q+1BnkIVYnh2hB5Jpcxkl03YIrAQRzIMnn6xX3XgnM
jichixdVN+8/G4dnrx72k5FDePpu2vS6mYAMQWn/YTBXQbeWUE/ur93GwDClOgFZuf2s94cD0gsp
heseHH/iEIN+80R4I5EgflxtDGJvInNbs/SonpFYI7hDqFfXn2LvfvTsygaDOt/4IM72Ss9brcSG
iGEUWEGSS5IKPeiEh/IxtXLJuyJe/t+e+E+JcbV7BvHZIcQZADs6NCd507zXmqPaDxkT3cvZWvke
hR4oS9GP2c7rOjtFpfs4S0ekL0UXq4ODGZFtJ1KUKv5xBXYn/OyrCibuUwRuWnMuru/HoUYeZuYf
6rPxKNmQ0/7FmHAiUT/aHT41h3ICikMzyE3tF0ZCVFeKu1Ul8ywcb02lczTQH7O6wwxj9QDm8J9f
0POO+CGwSqKPgllQ8hjJgTlhDPxcqbCB5HQ/nuQD16XGD1gJo+xkPsEM+mkU5+ImQYLwkk5yQSip
tBG1SXHtrksVVxjOq8szh6BdDz0pV6hwBOH5eaa+LWPz9plsgGNQxYfFzo1CMF7TXcoH3C1AxcrE
pcf3CjC5TbDass6kU9tN/i614+FCZ5iB3TU1QWK3AyyV98jAHiUSX9huDPKw5BUf9LYtRgGCY6m9
jShFZ2HJ4JTmZP6eLEKe+1ynWDqHgbj8Oa7Pe8USTfqi/ai9MMWYcnGtOqjIgmR1Yeo8PXd7Khcf
v4vTNr2InXT+YVEPcvqXytBMv7TNeJbGHRrJNKcDfInwQ/LBW28KlCO5/2bCeV+9XYWO+47NQGb7
4vd8xqBefIAR0zwt3TULmwKNZ0ugl2QVSdOo6gxOS8cPC78cIdlM/XWh7z8pXmheXcu33e1thtr/
KoRT6nhvIwCUkMMbjyqCyc+m0DEzfZJxTWB4jLz/u/G3W2O9pCrzslB7sAYsbd8iLQE2X7pTmfSD
mvjPoHzxEtx8Zxfrl4NT7cwFPTuxpC9n3jCCxMe7+JBtGJhtSDSFb7H3IczUuvPhAjjQBptZwuCf
qdsObfspY396dBNoRiWYFM3Rs5Doy3+ug2U+Ci+J5pFEU7Zr0ClOFdROwgSOq8sJGkL3ilgZhypB
i3W2nKxeJ1H6jOomCsKP0+t5StRJvJx7+tK+2FK0KVkRGVQl+scetpxVPxQStuJyd4AmvsSsk6EM
tkSr6tz5a5eGtuWt6wvUa/Pct1OhaQUD4kf8lBitXiuBDC62Exm3p8s9j9d8tPbLiONtj8PEU5+y
E41S0YzEYrehMli7oZxekfJrVL1qgYdmAH2jx/8r+WJnO5SVJ+wLirPriYSRGqVAvdxmIjYYnX3Q
dt17/uN/ETLCiN47bguEBV6zcNRl3vB1NnWUhuyhO+/+2aIdlPHYwr0cTlAwHsKEKxZmOW2I1CAX
LohDyG84cE74BTLALJRNAz0U7DuOISIr5Qm5JJKC1kIGDmQdaQBx2wceYVwe+B4man7N2ZLaiDkb
QaqUq0ZgduVYE5yYySv0pIGUdLu8d/4MC2qYk0zwwFt1JySZMc9VotJngWYVWYc+U9sXnyVsk09t
La6r0VISy5fn/0+Zl84QqzVo233HtACFpevOYne1AoVAO1zLnfT8Vo8SFgZPyjZa4GKkUr55EMq0
IEFiWO00kjI6p5U+eztopXfjL0PWSBW8zCsiGhntcIycFzm0Sjaz8hnnA3v1ZNsv/C93LNxzoEAm
MDd8lCCHuC5Q/Gjfs5NrJz3+/0v8Mi4V797s65b4gtILPVUByvuMrlXl2XfyVoXPH0aw/eewT+Kd
c01GcLJ4Grbic3Em/Q6wX0gfNf6exYKVd068RWV2qmEq3XMQNYmmLAM7dA6Hd461HWgePwsU6YJ+
HkeNzcQodZXk2tIjq6Zazh+/f0eM4wt331ZeAbs1eHZ16aPr+7Ta+sfN8hb1P3aDDpkQnPZsGa4H
nEoEg/u9f1v2Bsjc4scEprJBKIhX2mQ7O/bNc9rMl6+WdhutfvFS8pyHm6oOCenlRMyhhPcEfG+W
rRZ8I5dbDkdgLHdeO3YJmwbKMZsW/ZA9iVlJRTOjSma4BPKe58YYng0lsoY7qVF0ivtb/xZY+o31
6yDDkS2+9IO3Lrt7T4zMwai0RSZvrBrJaZMychF3VO8GV4BNlWHv5Zybky7uKslOv5RGNtNyOLYI
8NksM8Mb7wOUAd2u3HuboTxI8dGCRaw0tKCReqdUGonwhztGqkB6FURPSvumYgl8kqyoE0ckwkSS
dPnZkUQJJ/bO0IvYu1y4UdFfrhHw6CR95V5ACWPX+8E3/yeY13xirqLfBgGnJtw6ALBkjgJz+6ju
UMh9IeGA8snBPVMdffw+WG+Wc3NiO/H09wj2buMA2KplQtjnqsdfxSHv4vPDvrb/5MEO2iLmza2M
a16aAX/2CoGK8B5WE2Tw2emESLlzfC4xj08GC7/lzE6LvVe78XeSF60CxCj06TCdtgeaxh0RUKpu
//C6dGdmVGvTSh7hEMF4U0ea7R8LIrEoevSQYOnIpYLaDKEJPl7cxNPqLq3RLj3YTTwSSzS82S8H
w568nolRyWAPrHpBCETLbhVqaNmSrceRvJDc2n6KaQnibBrYiK1mfb9sL4QfPqfnwuomZC974/aH
ZEWwxwfYmQtl89pxTERAioLGMgb2SdKXkopidNXW0qEOpJ/rXobfrU45G/JF8FRDy5GY8Ok3Gd97
oEZjOt06rXvqT/0xQ+vbFpPQ9VLW5Luh3XSA+kqKtb0tZVrHpkZ9fNKMgsNU8CQtTTYCSJEQ6bSS
ea4HuX+kWqTWYO5WNFaoxilFk9YpvyyoxIeBUk3jhKxN7b0b3Lr1jGA6vs8geGxdpCRyimg8GgBC
JBxNuuJC/sWfkx8TjqpUnPcbLMmW+3o8QN3NZ3iPOTLJ2PenZSLjEgXfwjJlf5jGK438FXxaITFu
yEITKZajMyzuJob9N/5cec3xwQYVsYV6e3qzy0e6sruzq0a2P7Wt/zxKzTKFbMpYi/I+E/MzOiwR
QfZWTBwmqFjI731uPgloMtxVuQn98bJils4wel0V2CQXnMSxVVsTEDMakcL5gwf2/J6kz8ta+12/
1ufUZk408tkzyKLbaInX3o5te0PI8YnNgFIwHCKVOfe5r/StSH5VngBxKvYQxPgn/2E9xn1miNIz
Te8F90ooy4s16I8f/E3ira+dQ8HCqpGJeKbxtndHpjvVGL2krFP/NaNsESBO8lkXxMXzb/D/O1Pj
BZ2kvxgR3ixmRwWIDWQt5XNQ3NEAln54nvrcvHabHqdXrcB1HdeKtGaOV1mkpEup8PsolRrOspMl
np7+6twBdDew5NZuifuemDMT9oxi+Qoi7TFrcwS8FBlVIFfQiRUmuUVp6P5fN1hEoH1hbdI77gjo
+sBf2J86J584+q8You8/v+Zao/UNYXzN/JsRPwnrrjhsCB5Ns6YLm9J/n17GA+QGywWP0eFKpsC7
IpuLUNfZOIvCGI7BOpXIlR97f0rv4GgpuJqPyZFwNxL3FEGPDLpPtPx5DiQalBploDqGkTvP10Zq
YC8obH2VSRLkv3Uv2qjuqGSGMRMnxhe1W95WCeFY/6Q4aELKXoX0yKr1hgDwFeRQoaDn2H1f4Xdc
UokuyokmTLcEKa/RrK38l8c4fxS0rr87u4tFMtTlNING4Ua1uk/lxl5jqewvUmaDsYErpuCSubC0
sjyIEpun4wD3b3TuFO+gM8+m3HZLmmlDJzyzw4NrKnp+DANx06l3FP0Zk5DQc1XpBn/8GvknGTxZ
qkL79+zXporXm6u+5+AGWMIEoKURy9ohD6y98/ROgoRurM5ikZlQGxm99bGa3kKAHbsNvHPKbm8A
+yCtKJsnvi99Ir9yWqy0LBqn9qOm0tJCMEggcxZG1rwOA7otKX0x3Fx4xDVcuXAS8+hQp5uSZ47a
cfGhGlgquiCqbJlbsq1osSqZQvWuyf8R9z1sB3IDMLISDEI2oGOEk8jW3su9dR/rEuXmW/lY5QF0
J2QHMWHTn1+HOn2kTdmnYM725WPU3H4YafTsn1QEE/P/hR0BsbHQQldZgJQnmDgNZLZjW+uWAFtk
NsC9fldGb9e0Y1A8a12NlXfBGmf+qHljQ5JrOBzdmtP2B6qeCAn4gUIN/oAraz1wY0BKQyiGT0LU
atM36ViRjcdrZKs4Mdi70LYq1NM+QA4uB1/8BswJIkTN1DbjlawgoXS6hcTE0DjQ4mlk6WfokcXo
av2zli/dg8FmRIGA2Z1+DruKUhyMI6roUNcHYVhLmpd2OEV6yR8KydJeWh06iLAaEY4x780FWNwD
40PprgjhTrP1DPGT0Ya138ywEIUaczdn2mE4MftaaBZwVbxiZA6WdvrWJvsWuoaTRbrKosGY5nEX
hknVVuuFMX86JGE9rotRoQOwlnrAnYRxfCsb8+ZCBsWbDEv7sBeW+SbojvTU3NUZzR+5S2tXFBIm
INswLPui6wmzjq9QF6jLvzCWnUo6jFmfZL4lAHivEFtn30FcE8j9kXsg8KEhOcCu6qDOtZP+iPxI
MDaqIEfxSUJY+9MJWU2I3/bO57on/Dva9MR13ShaGjX40NLgm5JunFH6TB6Vo5FTuIpoMjicFMn6
aDS+aMjZIgQbkuayqCR6HjeWRAN9iR91daKM2+rkzC6XnuAFVkF1CXWxteu9ELKa+esVPAqlPwaH
G/wv1PpKpWJS4N2JCC6ZxVWmiiwuJb+y1EX4dXZnUoJoQ6Ma/BxqsCBIPRMc0y4aJpxX29uetGVJ
l/Ocu1C8ozL9BVj1qYp+PWpCiZpcs9byDqz+aLUJUSCv0vxyBZGAamuIsFIUzTtq92oFTRecHe03
Lu5PNQIEBgwY2RCK8G9FtyZVCWvjY+dDewJbcqzKK1LKh32qwOn5ACe/wIpRJXYD+YFWbB2Wmcgs
XVhyqzGD1uksIBE0FgeGQAwgLrEkZgZsWkOqjb4PG5ECfOJjlfBv3LxEKhymLGr3XH1k0CWs9VpR
rcWv6bd59e8JzamtaZa79n+JAuWxs+bSV7lLxxZW6LBA046tGhMhtYSY/AoDPvqwVs+D7uHDSFuj
ypiEkTcdvEM9NUy6o/dFBIPXGtqcYuZuazV15canRRqv0XTeALM97YvnKMSAtvaHvysGrTDE/hy0
1V9c/vKY+f51Tk37kWtdmrQhZV8KyPQ39F0hT6FSe6YrhL7WWlBehPMHOZvwToNpWYY6Dja8d3Yy
uw9PAGCOxK7z8EB9/ZNI0FdUeAG1rqCXcqADAh/MV7L1xmAU/b+YGwbRIgGol9qE4NhSYZe65Kxo
QWqvx0B5vKE5DOUco+TesY1r1M3rjYIv/spp9q29O1SaAVCoKYvhRlU9wr0Wt+Khxwx5dQ3QYigU
S6Vy8yb53yXbYvvKCYw0/94341prStELQB9z+PoOGMjAeALRklYgv+9Kinl6jcBmFxlGFCBhYJge
NdD8gGevdaczyuTryVzOVFcyAd9Frkp+Rk5kYT9EvGo0p5nxf+gWSCZy6EpQOt38kGQwalmg7uOO
pZrExHCSmMDdOV1PbDDMVuInwncjNhZ1n0sNmZO/irMdajP0ZchNSKq39H3dUhsMYbVnWvoMSHUw
PybHz1ONanMEMAlbisdQDzvnuyPFlxQ4fh6SK/Rnzoc7YgNsIyq+oRBYVLZB0wzl1lL3cI/Hbyjc
80KZFd4zyDD3xdK48NNSZhHr9/Hr60h8NvEg55xlldMHuo3ZHngalRyVFI9wwUx8biaoBSowSr0+
jVtmi0ZX735yQ4p5/62OX1XR+vxAN/Aa7VbqrYJdlOeIpJt6lT/zqGsq5QBPjGEtqxRtQUQBRatq
HIybjdgFtYgxkebTti2J+0b1uPm/hKI3+6fUsNeCOtyBfnx0nKMvBKhRq+OF+uiRsP0UUa/5pw2j
19RRj/bS1Ugpq0VRPhChL/uIDQRvW7T/4UNVALcVKbcU/z6IZ+eap4oMVQC47TYlpDVTeuF5zA4X
v/T2lpFkmBlvgvpAR3+lpjp/kxsdAe7isQ156q/YPvY/BemqHmSCntuiHUrJC8P/Ojvq0UC8J5DA
cX7LYY6hXEUtWPjxFkbkCFCzLT0srvGoiovplXyWIQI8AmpGT+1P4wGx1GqBtZmibLxUZ6svlOs0
l4rp+htIO2if8faRSRZLPd8JRvdhOp3FGSWRVx74CiHEX3S8kTcOQkuIiJXoL2bxfvts1y57pR/m
JNoA8GSSKDK90NSb2lqGORCndtUKRK7YddqI3F0COMEImsUDn+QJvJ/ey88t527imzBqUHy6E1Tr
BP4thlICUi0Zb4xHFgc5d3abjNTt+e/N8OhAz38KlarPOsmzdAlnQ6EEAH3DQkX0ey/XbKVXeh2/
u07yLo0UedChBroZEtFBGfBQpVzxfFji+0wgwtLG1BcvsTd1J01BEFcUHxNhS9cc9xW6cAGdo3gz
YohUpQLlsDRy7rKkO8bUfoSR5JXE7ecvbg3UUufTpIjZDQ4AdffqTwNak2dWG0HnbFZaQ9tCOiHW
rGagho/JhKqnjqwUihv/wTaERI9Cs+bTNlipfeZ854XQ7V/GlLwFBL62obm4uQt+ud7CB9yuxOed
iVlvYDnn+YOFvJOQ+iHoyycxDW84GxEZ4zJ2DQ1AzDu/aEmQjOd8yvi+Uog+5auOgXXQmPoFnVOY
cg2kKx73A8xZd5yheWzYqImCxQPdEB2FNYNFXV4M9UOBc7XkTONdw02HGu5pIEjO/Qo3Bp3n2gGh
AETXzcj4PUhspNISrqINIHzMyiRyPOlvBVJzi3bS9/RflACKUbhfRq7Uj0AbHqPW7vQkNVfnOvPR
YLtPushU0B7z6vHmrYp87e9PSqHKmdHJMoyrzqiolDUmu6Y4pPdHHZo40w1WMYrJvXheq+SiAfUk
WeOzSHlucA+IRB9JLcv1PU8FWDEQL8Oqgh9QMWZa8M/j0F05dOMeN1XtEjoQK/h01Wb21Wv4H5wq
11RtIuLb6vkbWhpO2MG5kC+2v0Fiiyn34Ek9oUrO2uN2AybGMBCAmpPVXKDWYD4xpqu4D67lZEB9
HRjZ336iDEoufcYEeFkuArPHcdocKMvlvCEaX6ApqkJLApdv0VB1XFd3w36bShj1plV0g+R77pM/
K2cMH9mWnraq0zoQaanggNsRmJEAwpfJx/4tjjrMv3grHaeOS5pDDeJdOmLnzAzMik6AoEjNDQ9s
aXXVWkSGsqdDRiz6VLjym6RlsxMC+JKptMNBJayzcM1jt3RzA8YIqicuFESx5S9ipcMelGl/4oT1
wego8xxbnF5uW+4ckwWOEWzVmdbIPiFvtNPpBh9b5g6SNTMmb3FaRZ70T3FW5x+bB2G0l2KHSTyP
ILddrvSeF2JRVfLOOw6wCDPeS+COf4EN6Vu5/0jYJHu8G5h/55orjeiveqceDYn2NxH8L8uj0ahh
R0o1wH40ff5Wx+k4NHA7QZ6k+bCW1+wCzh7RHYjBcCq4qryiyM0NXL+KQh2ybDXELDF3iTriVKJR
bcp96jZTyl7OLFy/qV66NkORJ6XNTSUUove8NA9R9Y5y60VRhm3tNwllMc+MiLQKtIWWicjGD+H8
z3HbW/NtBBy0cyB10DCdKTmu5DVxa+c/RmU82kEX/6vOMt1pVDeq1NY4OeSgJosp9cXhaeW3GL1c
Fsbf0MSGpRSFRycWRAPuMEYkB80LAWFwc16ZOQZB2HHEaZkp6TqJjTIdOQSV2KiC6H8jkCP2a7PZ
LvtMovupifP36V/ecUGdjlkbIZ9SO+VKfIEsWKCD4/ESnoVauPzaFj6fLSp/WOtGKSd5PksPB2Fp
IFqUd8mxH+VOTaBBJF2mAuJhe/PQCQEs70aSOYfil8ziKsnMls4OLpMk1+Gg7rgR/2KHRV2kMi63
86tIxKEy74Ki0lzdC4iIp1entFU3IvwJPbwauI8IVIrlLyX9GnCKvgvvyfSqlevkF1CPoTkZkQd2
Dslg+COQ8SxIFPAE8EGgAx6K6t3Hvq6FIGp9pZXiP3j5RwD+dzRLWDhSU/o6eAGc5tn2R0yZCj8w
h0NcGY+Zs34FW9FgPThij28x3E3VAu+XWNY7UU0tG+Xd3hFYBnLf1s0sCRPEhP0vOauwoQHQiPuT
eYiUB30/tdhdOCnmpRJCjWeAvXbUV7atRzCvhN4G+ExnlpOWtBHnEJ475fQLX9mS7g8+HFyDOskC
hXSt6ZxWdB7WVdhFz4asTmJw9FkP49Qq70eqVkLWmGT5QoeKkgj49oX4KFj/16eA6HpBpS66z15g
IPGeEMwxyxL3GZLfpnKfzI2cotU1FL9DvXsSYPNoF9wRR//wXLaLqC1iGPX2LvN+ZXLjLy2N0Lln
4qtt0vRV6crednyfzAxCP3s6UcAiCAR5TufT8Q+q4KuzZyG6gkybpjdcgQhsUdlThQGEfaT07I54
+O4l7zgm2ugHRRN/aX31rzIzLlzY8DPumWgopIGaIjFz+x5yiVnSXyx4InGKxUTemKdRa0gSDbpi
9+SExOmjxAhhH/toLv4f+t4fXcNwo/F/uM60/8/bNM0sonth9SZzqd8A/slCrNhxE5JwR2vSOkj7
FW7zBkllR/xhMoJqPTRssA8N3RRFXYlBlJqqvNQoGlZfJsOchUhkbg9zkaoCCJA4rW36i5Pm8RK4
BLBeFFgtt5723BaELQ3/K2Po3RTpqm51/ccnJi/qeAkMmrbosGOTVNYXJkld7qR28IZUcig8pcNT
P6LqQ8Pg+alPu49l5Tkr1G0nmWp16u0ZZ3r+L2o4dvQddFqLhqY1+uxCfUdu400S0zu//XbAnzhN
NoIE3ZWA2XztI9FVupEFIJg0m6qwgkl0mizy1A4SkGkci3N9nbpKhwuz7lqMpfMj8CZaHHg/7S7G
mWWe96/DTIuTLmp7i3oPXXUYUdPqygazj0/feLwvjf3qQ8SuOdMTOneoka+AyCh6z5jvCwweysjX
haXrZNc/hrlEYbrrBSkTO5oY8/RMcT6nJHpgjq/Sz2GFTNRGTUF5HfGsFkc1MnMaCgmyoVZ8QJ34
DSdzsLQa57FPeb2qkz5hgqdDchIHc+7Hzb3ZIFGtophHyDJF/qUpaeCfVhE1AFxd6+LPcWZw8Pet
1bPOpsK3+R7bDJGwKc+O5FKZTDnROUxCQQlw3IIEKdyzXBKVuankyyFoQZ8tWvxNVMld/uV3fCic
uEkOIVSAeQqiJISRRehzBFGhOqMIiGmq0QMt312xSOL0+rCVDLiadZSHCaWNilTZMbvBpJMVOMfz
K7LGOTLtCq/GJycnbSqrb+HFMzw7WvfUylehHc9c/QBN0j8iL1mbybekBqU4pq7mUFJZY+hppP6O
eT6LP5Y+xgUsOtXoFAPSmICfkjWCpiMtS6lKC4OPJqanJaprkQRKAshlyDOiSrlF8gG7dJklemw1
2Dfjs3N8Me4zQvm9KjPqYWpaWGS6QgehvrcyZhoIt1VYoucgF6knVN0kangf9rdgV4rddkBNB2aX
FqzOrt3nxe1KBJ+qmdtRJ7Gw1Ti0oAuzTDeg9woNnSp4rlLTL9Xe5LVf1Hj97J1wrcQZip+11cXJ
kRRoN3YoEynJN4EmqgY/MWMm/svpwcyaN1UGJ7Slac0eeMhccPuOIhRRXFvqN1aRrK4UBYQjOVl9
E8PgFfZ6/hYH9oIoxJ8tA0PXKAzP+5wu0qxoZ1Qn2EC9Fh2eAV4br3xITPgBfGn4X3GfivQz/XA5
o/bHCprFtcRoIV1uhSRyrK2uBXzIdx7/O7J06FMcjb4RRvvHKeBSX5/PIZaBg5Mnr0flKQpBMJAt
pYIShyVKIheYcCsPZRcpTgfquTF+bXkBNZXBN7skm8xoMAJeAnU4oHdpYdo14AbST8uVqY1jo1Jn
kjlBXeF4ilnf68jjkUCNUXqe9qemYq3FDCmd+x4fnVcOaQ51IiPqtLDrBstO6nJu1NKkQk8uAZx+
CHkbUB2zhFJW0Hby9GKmRGC5jSp9hNUjg95fbZEFZFIZhZ8Uo8AJdlEj6OI6WYmDHuSaUAktD4wW
DQiIZmznIxsO8lmAcVYDWbFbux6pmHEVMnzUyRAavVqYZtiTYX+4a1yeVNXLfq3qT+sL026Av70X
1vYk6hMArtKArjreWzwAWmdb7CWzYtk8lZ7i0CExZg/IlPYVyMoDPl0IqMZEB9JkFYXyAjMotGeZ
vjQ1TGXk+skSYioHXkIlqALmF7rVsHCQbQ+qFZk6NOQ5pHMgDBmq5C+85vtIkcdxWTjIarN6dddv
bDy2JyqH+wrpQNJFDAe92fJp8dDkn6BBk6NO/JaYIY1WNn5DCwnrCfFK0SxJY9JYliuVTmJ/TuGh
QOq1LWMX26MVQuNUYMdhqfZdC5m/TCWXxvDMnN1K/67YWblHvTZMnrKs1rbzsXN4okqg8oORCccK
kQbPpb9siBQesmHNJIViYnP0FYMNME9JAOrdFLBKlfbHwcJN2jxOzqFwimNvtoPOQHvk6/y/BZ8z
wZITr5izk3iuCreAfxOZGcuS35x+5khFj948SPBS0vCJdRKKPEvh6EG5ZIUZpNeWmC17Byo5Dh/V
GTZgw92DogKtjUASaGUUWwwQRpogeSeo5LDLy/bPG/HRYikrnODYgse56gqFhwhNIdKpMFNtD4xo
cugINqebyzT3HBzr4DreNf4WI8afebNkzDOPcGT2Z+Np0SRwLHQ2oKWSxo8+H26XKuazB6U6Bm7m
Mioig+owYbi4mcnnLy6zb6aZ1LK3vZgZX+u4iZqnsuDtDtLnpN4KHz3rJ2wjNh7vgA8brEsH9jiM
bN6OHhWA7xMg26onK0ZVrhJFbtawFeBn5nbIXtOchepdW7b7to7R79optv2FlXTvk/PtMzoXIhSo
Pd15ibruWRx3k2/2thgcl1WUv9UXpVaKt10fwjOBYA14SKG/ghsViusObC6lyxVMws8wiTHQ8qi7
MC552lo+t14zOBETUGPwhGO8duqh8QIMEwaOkxlonw4THPZ5GXBh+Qd3Y5lMSW9zFkO72mkY6iAr
XKdW6pjeLIzQtoZoqimPwsOT+fbLTLQGr7LyBb6phDWZ/PH+QInc7z6PJJots49wq/w2W7sXTFhz
TvwM+N/jrALqBSJ1fyDn+sP9D8VhyfOeTRe0q6YiEIhR5xXbzsa6u+g8WrCncEDs1tJN8+sPDwP1
fHgRhjOc5pVtfK1uK/yXqSOnGE84bOCwKzDQPEb/WsQ2BtRk8+2b9CLWS21VzU1OqA3M2XDINA+H
OAm0SBtgmF+moRKIWnWNYKYmh0HCNZxvn/eZvkyItmDjtSnr2vvqXqgIiMPUWMJMfV7SVb2PNII0
viWIjvTPRfv8155lu5GexLXegG0n8l5+TxEqD1XE78555meloiJvpKLfl2rrGERVZT/fwEiVKHw2
efE6aiLVbqfGdsBjJX6poM9vpoRAJdQGOCicUZA4iDC6TbvJNzxtHqudhaMiiVlM+QroDNOJ/K/i
63prYWWRHD7VJXLoAzA6eZtRRUN9Hete6MTbgRB7JoED8Jj8WtSF53D+f+gdE86djREVD5LPjs0i
mcNbM2I2a80t8OUdZsKLjedQEdqlKlfFcxcfIOwuOiSYN7IHxzuV6jVBlQkbfLnv+gv9Z4rUHCUX
VsBnx2i850o1fsZgdnbDvwPi5HTnryfmse37F1EQL7WNXyYUcmBKEZnxj21xr6D+ZMnGDgIK8b1b
tIm4NU9QxoWXYpLNUS5SY4w2JvjWY//vWOdqWNzWdgTzXlyYeASULv34S6oVB5GZccYMrvKy30Eo
jl2xqG4m8y+bX1YkvEwGiNZQK+VyXO0V0fIcSC6T+MhUVJWyFjwGjKNS9hnvv/fWFZdCYjaiXBLh
+W8DMlc3JXRRK058ks1xsRv6LHzIXI9Rw2reepV4I6YA3kUx1/hOYwPlaHlMTgqN0CyNVJe0WyqH
qYlsbMHqlk0eWS7Ov0jWnCfDRMFmafeucZGXhbw7IJUH3nFteSGf8e6933n1SM0ukFWrvGWYrsMs
+9mloAr0VKqCy8jfxTiUzooo6GFpzZdFTwafzhaa9zpwqTbWINeFfWf+SO3KH3AMoPM70dEkE/u8
JaD9FrZH1BzmFjj3iww3oHINPNS2GBj2xCFiDh17szLrZuERtZ/CUDkiJCKWXKOj/mMLK1GpA65L
9jhtAH8RdRDakWv1L62JZMuF2KumtKQ49u/+WHSNHYAh1TlmlMU3VAbQVtqhJskwI9aVYVTrMjuM
WOnKCl00FRLpa1WU4lwKocRdLesaWmdAph/dyTWOEZ419zgRn9roGo2YOVP+js3FdZD2KnkDR108
29WSNdR/uwT0R79C5MNTqnmb2rGXBUbn75jPZD+dJgiMBD1cAOsq8BNmkbl9u6WA0+vrV1p699zJ
8X2sJkgRL7NKtC3pwaBgFtL67AoonX57ZOrSuWLMETL2q5oA5VKXQ+ebe2eJqAEoTWWVomKxJgMt
czOxOxz5uX5HeoUKKjabiE2PSWq0eIZ0wUK9A+H6WTp9N5xJK+1Q4l5DcK1wQFByuTMepFo/iwKy
PUZY3cW1891lM+Vd7UtbGZ+QDbhxlEbTni6Dz9xnbn1f+GvUhXUhgfcDChtpiQXcpOzG8/huASD7
w7Y9xMoOg0/YZg9IXnRGd/zOEV69S4pfLHvtLwfdrEcBk2c1bv4mnSf5qSZxixhtBc7ZYlwecZdN
pRe8xl1kThJof95U7+tum0dFK+NbQFr9r80Mclck81Zex7X8DCV82Ht9pBNafHJDvM182/n/ufZV
QWnNjLtrRg7J1/Lr+KyF4ks3uNImElU83KC4jhxsI93DBvh8D9GyfGMgW40wGuM7PmrQO/6k2Qm9
4OAuFM/1Cga+axYkeRFfps+XpMymGf7moBEIamWjJdIbTaX4QrdsJgeDkeqJBcv0ocrHb/xkfRp5
/vtfup2O7rXB6SrkDCfvh50EiKUJQIjFFcVIMpylUrlsvnEKNJ2qrr7VEK2oNiuwqn/sSIkm4TPo
eSMLg2HrxzNzuBt4FTbnO5ObHnssN/Wi5h0AKYVQqe7ZnTuouBkOnNEbJqu9GhSN/FrpAQmySn7l
KJ4iSEprW4Qjwd7ndH5YagkE4pajZg6tbp9dO4sE6FX6rdTx/RYGYnNeHsb5pZwqGB7cTob3dLbz
1RRA8Abhm3UIO8afUfUMnxCG059SbbW4w5qrh4SWYTRD3VnMspKMfZf7dPEtUHZJTrhE8yskmphh
58SWxqrl/yC1FjUbQJqEGrhDi4HIvLlAAJxNrTA+qHlfBf5u5jBp7wBiXWsb0Ezji3aZF+7vDAnw
YjGAb0mHL1fQPDwI31u8i9BmrvCLeGzlwY8qGmD8KC9ECckJ220Yg4nHllYJ4X4VKH/ESSJlccn5
7xuF7e7RaXhZ6WXo30OhvHdAzeEULi8hgruLFJ/cv7uBhOVKj2AWScMQhwQYbLtJvHrMDDiLtxgS
8afuA2wlcLHgvIXYne2r8RECpqCnelAmpeEX6ZvlVtWdU7Bh+l855sHBGyJ3d2Ztd2Oae26OfG3X
3tzMCX44htKecvI5qn9vx90uZsu5tQwxgOn7yKL/7P/ZF11VnW3rswCpg8V+wj2n6NEzuubfaGPH
ZEKB6Y7SNuJtBQtLlb4ZAe7Uuy1O90vZXNyJzM4R/AddeJA2ZAfcGY4uJ1f/dj3rJRstmjOBfnbP
+YTsCk1CKM83w6J0nmkk5NX556003A0QTjLgCBpjuokqVsCJxkcDDvGyRa9D3bHh16rJHgI9KcFk
BJ5kGtrJQlx56eHDNulkWUNMHiQWgL5LAyLS1uEyLUSFzdw2tJQkeIC2cMHD0uw6BMoqbMgjJr4F
EibNyrLZOivgsufJhXe0b8rv5xVKjaFw4wF1GWQ/xHJ7tKv+hDWm7DwzzzeFplBruQCLPBc0seSy
PilXg+MjLWuuMdE7V9ZIK00kjMZ570+M3vcueETBovVDrkPIBwu6mWaHQeKdfG5WfnEQXUpIYkGS
jydDoaYAsv5a5fW9jzcbNBd/5YgpoHnzexphdB8YuEEQP1KCT3XH6QYoGH+wPN4g4yr9wbcoheh1
PzCrIL2U6gCstFp6dPQ0FaF/emjsjYArAFucCStx383PcjU8dvH8yhUlX4S89AzFBhW+deld+0fP
vcUKsW3eJ8m/9sLJ8FoOYWWiqDtR23VQXgK+HhUfKjOLL46jxCm176POwigw9aj6P/TWJyUlRAQT
qBimPmGksVvgr/isaKmU7JoPLdqjk/pgA40Nv4LYxCGauXwbaHZK69kpXKEmorvDiskKeO/Hsvaq
/RuS1Z6rznqRSgkaTQ8XnJOiusFRDueax/MfUKrPwvVQGmvYyWEOLiRN9rQdC87+eznuc3O3Lj4i
nXJ2Tn7tDOEJe+QqJvdNyu9C80Q1lXU9OsD2yAEE3+KsNGtyFP72W5R2+5JgOeMtVlpY3gK2S2YI
uLX2VAaw+m1a6uzSlDBq4ZD6hIUyRfB2SCkfc5/82EcLwxLO1xrzzldmaAJr3v3SXHyFaKz8NcvW
X+XsNAH5+g9It2M/P0BajLpVZEqC0nw0qNZE3HaUADWxz/4wAJPnZG0u5fof+LiUnkWZC3WK2DID
Zh5TjhU/obRLXk1A/4RykjkGhEQys4WzO+6YL3yZBfY8iMlQqISqnYxVbg0atS4CuCvS0zEr6U32
FtTZF4vRFkA8dWet0UyRZquqBYaIskjUF1UMKYCczkMdHk2vqQ7JDyTVrh3/jgETjbU5SYGD7mvG
v5zc+30uI+0yaQXHmQx2CTvN8NALKZnnooiA0NIjInvWcD8lc8j/EmcjUJzSdAK38zLHLLbyseOQ
gxfL6wPAog6PCwZrKe651CwsO7GrCrBKLZqC2daRAwlzABaPmXohNe3pGTdcNvccQ8ui9YbyPxMk
C1WkRIx+jteLEkJBCv1ukA+Xf04nHq0MCwSXm2Ndga7iTf7sEGbybTfTJ7WGKL2O19/iO7wwTc6K
I2Ke1QdYYBEBBvWHvK1vcW257bpHAHgkBEFFQLII3V3WSJLqqHrFIX4z952wgqYSKrp1gGDoZUDg
VRz3JXviC7gQCEKYNPDUY4+FLFTQq0Ww9KM0uI5Yaevju8BMtvSXFYXuqDSiCcTF/ViimIV56A/v
pqKZcqmy9KJB8ua5v7vi01+TujQ3MHjOVQvhj1kq/F0IbvB8/STqpaaWtlwfV85nbodw1ju3rHHU
WtERNxG5TWdnrLyEisUv/WYdGHvT1CJqNVqyiQkpfByukV1z26Bkb3Uer1xo6m0Be1XZpcB3TGUb
5MbChtuUfI/deSnA7iwV3Dm4sxDooKwOrTUoyep4tahmRpAmpKjp528/4UNMAXJYHOHL5xUb3fiY
ME5vMJQDPtwz3xGXkTgjWxi8ZVitY12QTrW89SL/SUQ1kXtGy1XHVouFlgtG8feZHNpnzcI3iqiD
XFvhHTgijYlUIqFLoStDmql1Q7WsQOfMS9sEqTYGKzLTknns7hxDvGWSMCRly04MjnC9ufvqZeLy
oR0O2M/O2K+FJXxzZHqtHDl+3Uc+zkZ5UOly4O+1nXiTI0i6meBRqcpBL/dXvLU7OUAVqsC2AMvw
Kb+AQJMvZe5s+oy3XzW1FdmKrUnxdVTCmqRQPdcFofSBwIIUBi47+0W3/UAU3cFKLMLbNptdeZFX
1cPLPpeUk/DsTjJ90AfsVTojRDBBjDcpDvBaY5RA3zxk4AJYfXpuSxPhULhipc5ux8YWVPblXHoH
RKiHqEIQUpm1NXtHFAigReakg3lz7EIZtdP6H/3tnwC34McmVYtvX6nb8QbkbFvgLbcPBBd9gJJx
2OgrFk4CWkv2qE5lRQOcc6lOATdGaJhRq29HushbjA7TVgGVSrKpJZ7JJuFmZjfURWqu0sbrsJIS
EnxaUcQOBdW2muLMoPB9TSQCu+s1eCuHyjZYGb08nZxz8UL4P6ZCLNjCa7U3yZH9VN86/ppXJnyZ
Rd7692YG0cF7Zplf/MRbCWCM47QjYuAv2PZdfNPPyVS8hpYLGqZOSlu4t2DygiLkMiE4fFxJZ4bz
+8Y+Sx94Y9m46UxR4lir+T4ChjuLElmS9XSn9Z2uCanWfHCOY7VkIVWcejSQmxodsf0qqBR4Ij0L
QTy48U8aqT1HWLy2J3E8WziTm/KJldMbNYFjQGoMHMgNI6/sweLlQOi9QV04H/Ud0ttSU3QYy26o
c2q72lfQvQVBUNMS5YExt7ubLNompD/a4xoseWDkUWfzDDCG37abxm2uVpk3SQR6pD/2ar66eMoF
MeiENchgoonHiGuK4p1eAotxB3nVysmTuAfDe28mXkSfxR3r+ibwjpBcYIIN6loPFnDCs8ktpL75
gCsmUvIK8eQSz2AGB/oiY9CTyPEBvnAFFcjyhS/HBLwtGjSNhvgardGTMgGD5UXVsPOGZvSUnr/p
EKVKFVy2VDPhJrZT29V3pljsPcY90c/tSiVPQi3e+CNlzZcV/SlIkqlQocKQPkFB2GFh38g64gST
POTYD6anmrciBtpiDilc27BiV096RgXIHWPeH/Dq0okd1ZN1wzrAkKrAkkUZ+Str3U0Y9qht+xSL
/iWWyNdiu0Eym8z4QtLUNzTbqvzGtyk6YXv2MOfCxNUwpJdgDjrjIQOeyahDJ1nWz//6pFBw+is6
aUJSQWe04iQt4cGLfQUYODbQRR/JNBs17pGzxA/+8GtPJGCiyauRQop0tIb8Q5DpLMuRVZhTKB0W
buQr5+jjkoFMtSgxbcGiIKrGFThukJ6GdQ8EwUbtmDZEXl+wzQ2CbnMISmtjaAcB+3hTexVSMzm/
B9aCXOzuJG0IsIavUAEN/kNxTGVVR9w6j8fonJ2vGNAFCRRENiFa0Sqfjqu+JCSLEXUCOYuOeZM7
fGBVbzFVvEPjAzAg9Fw9Ak8YcxKgexcsIKj0Plk2uFeD+u4kaEBRRHTIbbBovLphgkADVp33evoM
IFVIKc/EzanIPR/BDKxwUfJmcZIAN0o8TJFJjWplfd5woC0VKdK1EmRSl5LsHLRxs/5szznT8NI8
WxdkwHBTNmENwnfqyInW3ZJSac6pBmhYufHQaX2+VjtbY1qI4ukA9GMdTckGT0mXtMNucHi0NQwl
sp8/r2tXND/R5OLOO2plSz3K5ykmzlqJW1MX7IbccEjYLNFojq8IlD0DF/CBGGnY7rBWcW7L9Gkz
cwE/IDlL3lfegcuIpdOiaHJvDDwKoYTc2EV9NoTjs1hppjUPgcWeZI0T5ebbrPZe6KvdNU8Kc/UU
LkIDvBwKVHhbdwlkGez3gXJ5oChuNqEC8dSpIuLrs5lsqK/kKU1dpR3L6kTfOaYCTHAVPSZjfKHa
0SVu9rspmW8c2J19NCj0Uo1UP1FHwevick6rOc6msKbMfl5ZUKJVjzk9L+AxRo+HiRNa8EbHkSIo
7QXsuhi3ySYkj4qNKDmIB8tM6zc+8MtReZLWjFFAWlxiFF823gV56qte3T1Hf7Ptzca+wK8oeGg2
2RycZOOnGPXjy58AnU+vHYx1B3/EaUvSc6Afy+s30xcmo+06yEd3WpTXH2kG0+virhxV3D+yOcB8
POwLl+XZGnoILz4X9UPA43emlqhZ9p2hGRzbOdKfbZxHSr7GGryI1dK4iTnf5yxx+P64ha7kJrWm
ep2G/BEKpqHi+kJfZULJyxN/++IZ4Wfpw15+RxHN09NmEmq3CYDjIOgAPyGEIXaoUPtAAm30pUbA
VEsIXovw7gUtXmksC8baOPEZ7o0t1qPXEuUs3LvMHgFfZKbF+MqStTszZiFJXzf3wec+/OpeMqHs
0cvbXtZ+wy0A7knyFB2Jz5MHolL/3t5KX+tKDEYj4DMWXExm3ZDlX+PhPZ+ddjLcwzVR8bRc3G+F
hqUPzhQRwAGW5t77Mtrw7eJV+wcpWRGp3c8//02EJHRFz/tFEc4+PJkV1vuoVcVB6VnEjR3P5RiQ
Kl0Ftdak+e1dFcS3Ig7SxnY4WjBAy56SON7IXb5SznFTWhGGdCLC0WKZF0z8M80LCIlEfRd3WwCd
R6KJJ4vjLhC+WVGE+15OXMR9IPcZYjTQP2i7NjPRt4KWlAH04HvIwtFOJG1prXQ4NvEAvF9KGLAP
2wtRsODVnGUNFPKE+3lT8KRSaAlGTAiP4hWWslE4CNrjmkM29hx/o0sF9D+rMN6hk0OCzH1xi43Y
MRRuVkoDtXV3wO5eSUSJzIDCqowBcbDB1GKaCM6KcUB7DM8O1fw6aHzkG7QbnzuTC2+QYtRnrSQH
lZRXjzjhR0kOfhygmyWl2sn5o0MfGGNl2/3Ch+1WmB8vWMqhK+KH0fKQkqBpZo1Ia8XKPj0YiVQy
ivS9dKoCY2Oi5Sb31ex5Xl3tLWuPDHgGnikWqwKJYGuEvp4eP/W5EBqbgsOjIiuz5Y7U+IxKjCNG
hKEtPluQASHgAI7f5XuV0RQiYKNQ/0yt2lAUjWis1iNFUvQzSMX99YD9fVnI3WO4LCSBvXF/ykpo
MWdnTZSHK/PIiFA/H7WBu6opeeFx0zvyMM9GtR5NXaGMUSRLHrwYNYnZSHUfYKz4uU+aZabhLOVs
OcxjkDObJlJkJVW/SOFDLOBJdCwdMNpU1Gob2Eyu/OoxIhyuShAAoBNeORwW1NDS2Yx4aWzWs14Z
JJIGMLGQ95gqSRXQZD0agrWkkiKWPcmAwzTmL5YMVq2dyXiLWB6db6Guzqg7ge4pYmf65PIfoWgR
5HDeJFepFXvAClidNeC6aYaj0MMF3kADFxczXPnWST2VIdSMwIN+HW7fQ0MHXKqrIxVEhvCDOjQw
hae7TUo6CFN/LWpR1W8QcCWUXip34w06OvGrwiGmsSg1T3+w6ueDXj8DQ/PD0nnIGW+81A1urP3k
msm3S18E3ltXWpsLiDKZsNYAwnJBJsV8z1GBv4NX5DV8xLOQBxRjmpQeag1VvViCkUgP4HzCSOaF
iULC0Z3WP2eDBC2jPf4+v9f2+k/DC0BXf6A4/UyOD4CqFvU6q5vYsUgwHcVMO/4MOoSJl0D2Lx+N
0V03k4KOPY87Wgtc+0C/ib+iYfHp14V/ee9CcaHr0TcQ9WI2klrvLnYfvY4PzW4K16D/7hCAQCAQ
816RMfaALIGEy7gWrMwBsMWwTBo2ROHXKkIGLGROV8W3qI4U/HwBhNgTc5sbavbtbns7o5ggB2h0
ELaqDdvd4z7aobkM1lYHEUObiMpAPqBHziUraElZu9UAluWfO1E01AHhCisxcv+H8BnWw0vhpbCO
0ymUnfp3paJ9YsjUFnHdOA5NueT1qf7VLe+orEh96PwKXw3tVLSd5blLmNHOmchZ0vvULsgEDTwq
/Zb7bjpcdGq0h+/rCWx2xsPY/yqV1dIhaioHSdLwftXbYSLNCBgOqHRJXCtXSbiQTISRkM1LfaNS
rQMBED4TOa0nx2ORw85OibnAh1N7gc0E0DU3y1nT0RVm3aF5YAz0G/V3wTUi2hVK8Fw1jY/tq4bl
KDJG18cWigh2iGkQO0X+dWqG9/8X2+HZrO/Xn87118ISZZsmSS5kW3Li0PcKB9Xxdm0zob2d2SIN
XJWnLpNjYMpwWNrJ3hHyeJAwC6cgNg39jercJvPokNiHhLxgFscvY6N6XjbjVuU338iY9ZEE6pRP
U6Hcjc0X2n02pKDcQlwP/5ZOK9sQIBSA2tRjd/w9Bj9yXaqx7Cm6iN1l0ZUsf1Vg2S/1MIf87Az7
A31YsUQRZhSpvUZ7GqgNR3exk5w4YvTdb06KVxZJiiQf5UbKHf2ScefFihCS4HyIDE9zw3sK9ggS
aVuJpcVRy0AgujlRkoF3bVrrU+KlaRizQP4WM/dcaVgJHw30fVN3jWx2Y/Pp+1JgLkIIqxnnx/oy
pZ1oSLst/1VBiy3C/cZKf9FVVNByNOEiZu798dJdypNQML45KLD2/Z5/Js8GDdBaBslt6fSggoTL
ojYu2XqiDn+SzioXtOdCHUqONJuwAgq9G9fJNvzrGqPTWKEg4w0ZKL+S+YP0q/XvL6Q62lL5wJch
RmoUp0BOgb4IUru3KBqK1XrbP0YplnBwKn9Cq5yzQijJnqDRN0KWnhDmPxJzvdz5c5EqI4d30xD9
iVO788OYeVtttT+N+ml/ttTAXU1HgOhKwAUwx/eJo78ctq4qo47dkriGkexZ5tJxnht/mPKJVkV7
j9nA+XaMjWi7hcl4aWut7cCNoYT8KilsapBwjYhbhVh2hd1cp0q9oWa04Q12Ir8y9iDwpRJsbhWO
GKSEGNe85n5dizAHfa4ou3jojqCqlculccMIi2KasuQ5Ohui6QO2qxZ0jmye+6E/m5FJ4la4CUEi
pKOcrfq69vW2BxVmhBSYEI1/6K+Bxhuo6wtrI1isVroBzcJheEcuAsoY1VVmqTxzOv0da6iJVG02
4Hb5r4E7biPI0YpZpT/6aRbhUWPcHn7kO1G/V+lzAHZnVbbhvY/Kvq7JHw1MxcAdvojYB2cUQ/DV
oWH17cwfHq4MR0pgfc5O+0idn1y0L+NgdUmtspYTsi1/ZtLKH7Ipkm7oxNembtJi0NcUX15lV4v3
nrulMLGbSsxRFmyrQ6GPFzLYzjaahlJDY7BiyTmmaX5wGL02CGXayL13KoRJ1KAPCNAzuDp+8wXy
YNq8W3+/ZG7o+wK/tGLecBdxPVeCNdgLuNb+Np8z+PundWSWwr2vnvg56NfT7K5MeL2gJLNPx+hu
j4FmHE1usC0EJnRDja8HlD/Ae/YQSjglzDsIGyyiFYs9P+/IVpOyzzWZo70CTWWbOYFQ3fy20dMq
8DULNUOKSJFLds/vy13q2S4qJ1BsxN72twfEmIvQ4ALK2dJIX5i5Tz2n2/KkxzNNRkT5kqLb8n71
/7x/uRHSaaaBwbPVerC1+E7MyQh8f6c8fy2HMIpF8gZr/oElZIYG7pgXkiJRdQiXuSFN6Sh/CT6w
qmU1B5H+r4LUWQWB3vdKsWroXnJ1mgZNcA+RHwIIfRkJeqFFg2oSrWheRkah5qybxtYYoK3HR1uP
NSPuboD9x3q7PbHFHx/si37Ha544lI3LETNlg7hj+yPtUF27c2ylkkhtn+JOxMzvM2gwTPkxLjCq
mgf6wGrD8byvpWONCZQFVohzz0uuoRjS/Ue6BxU6ekT2IAjDV1iLoambDcT3WlXFa8QhEU/1mpyF
F5pKzNdu1DYCOO3SjtNMRioaB8UDRU4IdFIUL1gdRrCpeMS1QhZGWLtxq0VdJqs4/OI5R02nkPLY
jVLw/q9UYZ0TEndpiGPAZT06grJ6Sf631t4iVaAp3qqHw/7v9GxZ041a/cVnnLmQn1L9/pgyJeBI
/yUqrckiE5QKALiPq4xRC7xvDh19Of/ZnMvkGq20QvIYImhU5mzsANsDXA8RuQ880tM5o5sRsCqk
U2zIGTWkmVTjwaycbXjN+XqUDN3/BQR41p5LT6tgxv1lqxVIFhosF+J/GHWor63uWKcJXsfZp79U
AMuCwmJsu01FEGXDz0y8KnxmGdqQBhuN4yYrywcADiqTK/khSFx2jtZPKpE8yEXqvwMPbOUO808p
hjAlqR6L1mHFKm1jM3b/kqH2xKLbvem+HsUECQCnSDn97M8H8XebXN/A26PX/KcW+e/h3J1dc16Q
7Jh9rXh1IrFJNcNlnZAUIdVl0z/U/TYm5gKFZcjW2O0p/9sbbMSZu8XR6uAWA3I1Qhxa61iLpkyP
+T5eB6jbcmEXs9eNTes+8n6iP1NNhXhvdPRkrxwn6lvMI2iCcA6iLEKUsxhnSYziezsfY4lgu+fD
lIK00sfZCFkHEWpefRwWzyZIZT72A9TyDJtGpVnaOd/j9pDMo9hLRTlQ3bQ6jnn01yVxr6Lxkl0n
L9l6d6Dc4E/cnmeUz5aQ+rDDztT8Brr4iynnJdhPTdU8BG2oUER7ArAeQdk4g37dmMSlVm50w2EN
dwAeD/i4t4oYrTHZVW9Hs3wjtK/iwSOE9l1oaEdRt1i3q7WxkvcPExzNmJG7ZRMLARvAhtrIlNWd
xpXrxGDC+wGwN8Yz5VNUJWx0N2C3B79J6VcyFQseWT9mvTkbYQAmuFR6bsq2a97PijutyLNiyyqB
qDOkNshnmVqS7UdWaPZNNsGkyOTc4ebUIKMUi/TauPpBRXZDgFJBmdXgxSh75ss83cSq3V+AE204
pshUWKbpcr3RfpgQf3v3KR5kHv2vu/IixIk/VlkrjYyP4uSt7J9baFawvqlUWPSMc1zDmB5AWzat
VMaem9ZZjaQLrve2KZZM/G1C8meQBHEw878BJMKs2fvAQusNY62moT0HTBf8at6VXPOZxesi2jfe
gh5UhYdkm8LquVsaqHemambIsHe8Vnmyx82IlySw9VWVYsW5Ne0fImd9SS3uIIL3elt/w/ZD09JK
3m8PfBe1TsqrY9VQ1f6zxVNNMfyVNXMFZUu+/hfsVQaEbna06lkLrNhDoZSLEj/rgL8oZdIYXjpC
MJOEZnHxrho5aydIiD5SlG41156PzRRCpsvsIcgv9n5gybskm+j1DQXNoOXGNQ9TI7tMhBWGB0oP
T+Uqt1GrObO9u6ebki098joZyUk/kVqFcCJH2XFqnIxp6cv2FQpxd642/PQjayHXfzWNgiomUTD9
silFubmUapR6pV/gDLGhDrD5bsFbbXTXO2yvEd6Sfo4xs/JataDjFdvgcOreJEPWaDOO9Wg2+ick
sP4SZvX0Wwu/pHhEWY8qg7NZCpLgr2F54IkaiArEQDDZ7L/0AUCz1vSjJHZT0hzG5vnhvlVsX7hm
9lpVicqSx452rhvHzZ/OxKOuRohu29YVmWQoFOrUEqc8bhaAFCH1lRRfCJwaeAOXNctUZRwtzfcc
i9YI3+0da+U5Rx47C2F5h70O1P9rptok3KWK+5Is8hyubQHvyvxGJM+JNAcS7miQXmWcgYGRlQ3z
59ctGFvnC7/V8X0dGN9X7LInTZ1oD9rEOTZZ7in6jikM4cHyxFPX7LMg62wajaZ5xqTDajfwx+Ht
w4QzXNTOERFlMbWvY08TuGkI9AHc0dGob6AoeAQaVmz2qZvIgS6rLssF2Xe19u7lggS3Fu/dZP7m
TVLfH6FKmwhrIeTHsTl28aYDBBGtMfWJLJcV6Y5u8by3nx/LLUlki/a5c9/IRx5wpT23AlJkSyub
mnIC7AGIm9AZgkmC2FsQxghm2qBtC+LgegikQRcTcxEg4OAc7W56FxwLilqODqyhm4XCN5cTyRZV
VBU4GBA3urdNg/+Pdj+zit16N+FqqiQlYzd3XVpwqgWdWbRJ2elyjS2B/xgY+gPPgxL3pCL9xL8S
sQbCoosIqClKAP/vLrbjeZnM8RoMjDR48om+GYv0c+SKT6P9b/ZnRIClfJTaGpv3UC/4CyutQlnL
MRfwtZ7jzjYkMyrVjOnCXNkqDVk8LLxaUDlbXCUasbXs4J1hqZ3ktn4eSEkcV5P3yG4xlnX7BZa6
gWBENNZlcgZ9gqLYiTToyTGrUBfQU8PFNW9NocqF0qZspClYM9EKZy2M3Oo00YLjLGu937m1OJRC
tXvd72QVaQretLjFpbifcRCfyvdM+Zka9r14CwoCij+BVHG1YX42C2NolQeWXt2gCyMiN5RkZ/82
9363vKSzwPSKm7J6ufgj+ToONspq/G/7DnJsEw411lBiTt2IqZ9vP4g+OYVWbOx3RsFD3irU9mOv
/hT2RznuZAU3JKiMJpSXkkxLRu9A5HBVpWumQYnUpEq7iQnjJ7VBAx7kjPL4zZyLV+K71gcPuNWb
tFl+jjTz2bsVRdY2L1H17aqCl4Ax3a3iANXXZkIOgj4sf9fPm0WQf7h/iQ4S4LzQWUCqm6WvRJ+j
pxt27X1ANAFmMXmZScfH9WhrdYpHBxQ41+fDRXFGX3XlFuYv5QXaSB/xxcjf+rjINpgIkGo7Ez+q
8gF9WIbRw6eAUvkiqN8QNJbC7HGwKWEx01h5p/7XzTNvllYPrKcsJfbJ7qgqau5s7jWSoBT1xQ73
c4Jg4AubQUYdIvbg4MNCPMj3FzTtkbEMKDmxiw3FRkeQ6CSeV6+iktKucEuvLWQXYBVXG1tb+K92
lJaiNImv5YJ2uYCsJDJ6ZHVcPYJrMN461+YCIEYs4yhVz76f+VJoPDoIkJT7mobL0+odFzI2tcNY
50zbbubgQun3A75PYQGKqLfooqEPVgSyQW55wdoNFTNNx2Poj8/VtLm7ABlVUkOffSE/9wB78kBr
9//mJJzSbeEMi7GLUe9q6WSb0Ko7QaBGLhWUtp9l9x3RVr8ti6lWIo1u46SRJgQ92B3n4beo/nuz
PLBIApTc7LsdPylQMyZARMrJfFTNbHK/9eB8e7txM7wMIS7Gqp6JjgYomV3Ok+tYRFWVBDdnDl88
xVm3mtLI3Vfbs+xt3DF2p526DeKgG9e6Tc41kMecMaqW5/uRiOIxBr6BXu/hLj6mMpaNJ+jGkQSb
fkTKdn+666P5QtruTaWBt/XlWVmRnTgcZRazHsqeGoFc+s+GCyTpJld/TbTD/8YZUjgRUDm6tNOC
LpHKfPZPo20RGbdxUMuLajOAC2XHn/WbSFqr9pAzwZqOBZ8Irzk0p3tM9+lImisOxE+B6p95+Fga
AXC0jBH97oBzMv3rZP4ou2JrPWiBIFvfBM+piC8VG3CWEvoQNqXOKpCLjA0nfqrcvwnAO/dCucmr
ZflTMrb2XnwKuZ2jxlLJfb7QPwF2REni3rqstM71YZx+xMN3l/Jjl+rH8gqt1hzmNTp3akFc40qL
RdxZsj2J45jaMPv7xqqIs1cj38GzcWnYJpPtkzAyMOzVI4BCH/imgsvvJzlPNwy/3b/5xKbRLEk9
GX+k81lzSdb+DDNmAQuQ/Ej/fohrSrNASfH7xR1ANYZ0JYnsJTVxDI8Dr8vOuyIFCJN7Fo1U6D/0
Lbwd7jWWX1eifQXILKtgnh7wCpMrzIOYtGDP3Toh1/yMMsXmomlN/ISGIhGBNuZXrryE2I/IUqeg
0xRcdK7w9P+ZDJhqOXIeSb7cVtyMEJISLa2Jcu/59hdptE75SObvdWeGYwuZ18Z4M+gDSCP70ZXQ
OSPSKZFj1MCHtzkL6B61MrI+1B+L60B9klgPlfmEVY1FwLvX9bh7KGYC6nzashMQdAe9t6gWXaLi
KO8x4Z1v/7Mc9CFood370aeiBNYHkjyqsQhtdeh2uNd5GxsjXv8KD4nM2rWxQYyUGVnnH4ViOae9
LDbkORwc9B6vuj2GEixa6N/nXENW+3aGsMjjzX4hEk7eQsqzxukimOGnrOIsxfh06KYCbEVevlh0
nsfjhikyeNYeGdZDsRNns5+Xt7uhAK1VL+WdCVHSu8e6pelN1fCvYxS9PtTdHevPnrvNVK+hermq
oox0N7cnfy0p8BYms1UHBeEqDkfl0VrjYQRx2Kf2UZSkoQUgdw03u0TVAwu6TsK9A7gvlE5K0OSC
usYk5y6sGSkLu8UzjxrYOx3/ZNpfQYLOQwjuhezNsTu+s0ga7t36HMXlE9LbnNgjKAJSZBK6h7L8
Izf0oEztqVQhlElYJTkScVVMJrvZRo2KaFJs9icTQJM5v6IDPNewdOzkLOvp4lsXOfwFRJsRP8tb
IId51QQfKGcqZKYL5EBqxUNRoogFtvNpI7wFGBpLVDaGmpUe42WaoJ/SjsnAkdlqIHLzJZLCfZjC
0+rMMEfb7IZdVozwmsxtp0JxxtjK/HI0rQpUS6O5KCYE6ZPhvuFJKBt1BVIjJrOT1DT+0ab42ZIh
yDsgH0mO1P/g2IDqYSaJLL2YeOAoYohTe2XekYboitXZ0uBklimmPM5M2gmjUoUJ31N8hTjLbbJw
HblHZr2L5/ozofPY7nIEX0c0sXGl+AnutikD0TuPzKKjysHmw1aaQclw3H8/a6zrsU4hdgVKXLst
gq7xZqygrDOoR+bklscD6TUoCnMMNgLt9VZaOqfPqC0rUHAi0bgXUOGK3ixiMvszFaBRuu03d9sN
bf1YRaaGb0gCbOdskBgkNqY2ZXjLVLHrtI/0SNc+96+7qzA5yFwiyfLq0Vgi4f0yPj9ud9YdLWtn
qnxfMV8PHhJP+lVgkl/GQGRMbohLiq26AZyPQ7T3k4qKSD2/yfH1necuGQM35PHEkfelcT1RvzmD
uppa9+pHNblmDeLh4DH1l0h+FbGPV/rrc+9mW0Yr0T5qyjPQ3KqSQMb8xYEXRw/pRJ5DgywXI2Vh
+IYpyJYJEc7Y5EsI2aQ8BnJ9Xk4qtOtkT6HPNkaIX9MmuancrLY40c6122namEYHaP1uxmT3DbVG
eAfYeKS67DU02JKN40uQWSivbqAafhC0W8gkmsrunyTh36hymsDAI7tS1Lx7S0ote5EPOW9dqjPA
YKPu1yA0rOLvJBZwNAMLkJAaJ7mqh23tPXGWmeay2srXPoFkAuXlmkyJX9A1ic+w3wNTxhvdVnGl
/4ePM/7vJZ/s4hHaQB5an4tjgLHImcmLkCQcsy8zTnXPRM2RUFp0VTuvD5p4rsfjec2tqn4JsVRc
aM6tqXJmytgtmWJEw7VFFt8uRj2QRfk3IN1628q91HH7w16tUONDxtwx6cDfDCzbjLgp2vNyU/lz
8lCCaGkmC4+IfOXQJviiTy7JdXXRBNc3KawhQ1h+kp6aF+XLyZqgBPGHCnLwme2e3npKkn8JWQgZ
eg+0cjPgiwrICOlAA4z286BPRosVFgRKHVwZoSZOOaK2MBWcbA7kBuyxDcRSXMJOJ1+nWD3NjkQP
fNg6+Yc+Ch01VXf8NapHq4eOREQjMfjY8h+IlYRvtW2mkdJJYab/CtO8QZSdnoNSU2BvKlHljGKT
NIAXYSTOKqmhTP3ub0hQY8SX/P/RVnmsR765T80eI7cLE0bYxljzKt5jpAtvAO13vtLyvly8SG+C
tJIEJAYUZbbK8b0FB+yyGIanhfwaV37eKzzaQl5qAv5GWVey5L4sKynm8GcEBfeYtDUiH+4dVh4H
k2EBiBXUGScBNOD9RYhFQqu4pizWMV0+Xb9rYPg6m3a0jiZtAFtbka2+Q6nk7sT0yiam+6Q5o3C9
FoRGYdvp9HmfS9uxDmUfcc30AG9m1K6Jsv98ujHK3Al6p7C9hvv9ma60hfsvvIBY0m497NwRbtww
m6JSm8cLij5pR+yRqG0xmJN8UypF/g17yrEpywgXjG2dsDYZQg9wZIfwzHL18i5SEA0B4KcTmvXj
Gpiq3BIA6FTlc2FKnjgoTnOjRJdMel+VQ9coJwtZhps3DqCdRLSbnU6T1JAOZ0rZVoCJ3KRNpfa7
WhyD/z5tnWPO7gphIv084cEFZYRM2fxMi7KfcyB2XLMVk5oyEt26cUOKN600o6igEZeOsf7WPs7U
KtnWOHlPCHkjj72bVniOqDjb3tXZHujfpqHIdFbiEh5L2IWFfTEN1BF+9FHbXUIy342YwX4xZIW3
QFoeaTriJt2051mBFUviokNe0VVOy9WIxKQ1zfkGyqc2KDNx8/H6hDe4V6gOmyx/XL/cOKIkuRLa
lEP0kMILdJG9jvarGeKosH29CBM+whvAP5bC1t58XLd3O2Dq4llUPlcYfobHOjrdM7R5zn5f+MXm
LQM7MFPjVZOLy8B3Tgb/wMoP/sGpOKgDA2Kg8QpunQHb433W3jUv55A3ZRl1Cdp8v3BSbGwY616K
N3X5BiNnCSaNm8m/h5VEoyiCk0XEWiACLF+qmbAeCDLok+aPNP5ddFsAfDv635XNAFTxz3dnypdG
w9fq3NEL/ioh5DZqXo8Kz1qH4Dlf5ub1xkzoB2TbI3v5VcnT/aoWJIaBsFXxZbuwOoPmFSyZHVft
iyZ3hWuRD03UNXl2FfPOdLop7t+pGt3qK/aX64PikNpG3XkrY6HinYHYA5yBgDhfSa8xk43hCEGZ
idAoGgohYGKVRi4ANt9/7+t/v2Co45exWDCVJxi/HC4QauLXxwBBSpSlrx19S3Fe0rJYsLhD1Shh
2VO+aXWWkw3WMMRADGURshY5QVhPrNrbvV8TAkOMp68Zn53gMQlu9tjCXWfBAk5s5fYyS8vXNo3o
t4tU1IpWcyMmmVHR5YrrLZom5xVOUZY7P2eftFrTeIiKbJoaMqJXTNN+n9HxXZMownLStTJ56X7k
ikpLCK6az7q0aHN8d6f1Ma60BsrXEvLNVk4T72xzGgfHbpnUCE6XiruNWKIDhCxHJk2474RM6ibC
G875gyJJLqtdP77035+ZzsVjfMKJ3XQ2Cjv4gjtWvCmaTgQsqm0Mj3sHNa9WDKl29mOd+IAU7ydf
8CuEciuS6xyG4siggnm9Olc+ROd/8Ctw4YWhV10DCUDUehE+RkjckmrlwmZwQx6Y2cFp6QyZLhrG
mrZ4Jn53qO1rSLaWwedRaOrLLVE18+vT+zULsdLNS/eSdDN0kwVVKdKd0eFJ2aZQi2XC/o1yPAqD
RMmyF3eOTfrqTuI51yG7O0fuclReZOZ8iqggntiUqPOMlzCGbEAfhNu2Eg6mvLOJM1ei7g2d43Cp
Gsm7r7hdz1lmVOA5KKVUrPCbmb7l2RjIJhQN1X6dKaAWuKur9rVFUdGxwmWJpAv8LsJQXDZUaaEU
MeOIEGUkSIEat7e4M2SasBdYIqj0a20L3HbPe2a7JpxH/Qdit12sO/gyNCiK6hoOscn6s+Z+AMXT
JQxUOKeGSbtS//jyg9+C2KgMFvTlz47ztZOzP1av1sM4vsxuf8zpsBW8kG/w3fnqiJM+k4Sv1D51
eoWZIM2MuGwptYdTnKcA5xvLO/PYo7wIjmQ2l0t7DVsoiAwYrrLPjJoP0LAfuJH8+FFLuO8Af4Bc
Ys0puzl3Dk1FexOtqUKhxx/kcBjijmdvGbJOFR8WdrGJ+tFpl2TbxjolN9Bb6NUgPhjXT+NArn1C
Ky79TLMv6xSPHxEn7eOVDeM+b4sN9N2I6wUCWFzMfTCTkD9rOc7g4YSJQrHRa8BNYtYSAoNC5Mxi
AaY1xXjWDSH/axfMuirRBVnv0h5ivT7ugF4PojMMO6VTHaQoOaUaYDSUGwiBmDsCRJ/0e8Xjwla5
u966KKfwXtF/hlKJ0N3KOSThU8FunuTCkPVb2Ad2tuLwOKg0dW1qT+HHIDVvoBlcQEXORWJ0CWA8
yEly1tIp4yUiEsxaOBYYyVlxni9yr++UCmuayIPrM1Z7NGN+cqSK9N49GKC7b7YEqPGy4aZVD2Mm
0+UWRklGdmDIh4EWFTbWcRR9JK9pa+lTul/2Vu1JFCDXj7gMc55uyCqb09nleBYUURRxcXygKa97
Ey7atVHsMn3Imx/X+PrpmGrEDopCQF/HOudKiR+qiSHy/Pqf6isWkH7XrlDEJjwuiN6c3vXLb5Lw
8K5ko18fYACXm04r6qTLTZPaazNcf70pcCk1tukV9G52SBLqz+NFK/4QZnqmC/dbB1mullsFMgsc
CbJz53UsWCyS49cEpT8dOroRDdlvq3CH/U0qTWssszvg+2FnkLDZBQhOmixPfenhHWnINmZhzJw5
fWSeq0QPGVo4fS23ljyZcVxuc0UeyL+10BymDjl11I0gNjZ9bGulwddxtGW8L/oEZZuRjREaY57t
oJkgP5UHT1Fe+RLWzTp2pzbK2ir7IGzN5MBUfV79MgPyiGqYa2MIwLkBSR7+4NqamnsMSZF9sIMF
nRL1pEBzLnZXMaIhpoBo7WEtzX/GduERkohvygkxYwdalO+VLGRlQ4LQ4pPfIh15kAvhbIzEZft7
dJlt8+FIU9K7HMYb01T0QNBfhNucYmqMehM5NTCiczhVgm5xWwF//Ep8NQ65woxgmfDkS8L1uM/o
OFHhr9x/8NOWIWPNyH6uoFb27gKYfNogtkDKICkyx4SL23eCRxXWybE9+PsZy/UidzPTeNIynTs2
fWWCwcmNeaPZHHaQgqjnZYxA+E4YRHI6/J4qAuCRuN0oegOzPAGauRJFS4+7O+BdV41XYsXAQtZy
HP1PrqW5q6QkYHQMv/+mduql1deNmyK4d6prtHm4b+ZHm5+L2X2+lIMkIAuixi3MUo+HrdDm6z+C
OQQ4NJRbSSVJiKgYCaOUPDAhjy5kTvA5edk6+Zq3uBiMsoQe1/vi4+r1nki+7zD+GNI5LVAPBXJj
Vj1NZbQkO2xOGQP9YP8H9o6BJCBVQ8kTFJZNjB4zfXfcr7b2nVV8DiaLIuiQeRsCM4mMSwitw7F3
kvcgmVk+6UrWwDcTRTkVjx7VMsUP2nLcpDpEVceLM1rtZZG3oAi9L84OL8r8gYmiEFLR+H04aGvj
irPMeufbW6pQIcIoV9wnIlhT16OZXLzLtzD5Y8200In0BJlHZKdq7xBsgMhkUz/QOlyDDIfTWb9G
LVroj3nSLWQ5vYs0iPk30z2/57fGgtoPIIVs2xqeyTMzSZdF4lExDB2SCfsLoGTCfEDl+QXJT1rB
HoAD3c3Mk0nN88vL31GFziY7sqadxeIKJlIPMD+Lv4kEonmB/+ZNr2/6a+65CJFEpMIDc2S1qDca
0VP+XpUufvsX0hem0e145R5pIEXGZKbo8Lzu/1XAd2odTJQEWk0woSrrIL6ePTVW1LR+M8JxoWqk
LCak0tP14TUNXU4talqNmkhO4r+m14YppUI0wjnT/EQrISNbSH4pDmrGO4ye2HBpaP6y0MjN1bXP
+6w/k5UdNUdGKWhgYiYy4rwtwBiQTIg+RDFkSqpLgCP5BWJoWoCUCIwvbXjMy9A8mOzqcoSwUyK8
s/vXgOhLMFenGtujj3I89tBkxRG88VmJrguLDxwl9nreiRICEv1fHj6soROheQpx6tCWvZQINMqD
PPLPUgP5I2Au4lRZp/3vZGTrMMkX+kSNGcSwSzlvTbgLWZKw2LVJfm/o7/7O3jBwP+cVCC6X6nj0
S37s/DsoCHdkVR6DWuOF0IYTBgLhTzvdn376iNR7xtxJ2tyr/GkwsUH/FNpmgVWCVqPd1p0uJnT6
Gv9+huEsPjvWyu6inubMtsNxbOpgfwAWivhmx2TwgWpv9TrxYaa2T781YLLThHGnk9YuoNeJW1k8
iq1ZoFQOdTXuWkBH8aGWqIV7JN/NWBxvxNVBZB0DXj6EHib9O4SIned0bY0cqSIrWsd4P0VVv4zH
/tDVSvk15/tgpFAEx3dZDsXgEbn6gJXgiIfmX7pyjkMHws5Jru0N4NUJKWMTVrhZyK/ESRnekUJh
F2zO11HsnC/jgMB2f4OWnpj8OV+AWdH8zqJ+4eCL/NUigmCvaLtLittU93lLPAGVcHmYvMgNTUl+
GK3VQpd1kU7LtnJR0Lc+HZIoVGpGHImp2Og6QczernOWUNAGwtDb/IOxOcVpVr7TrPkuJO6R8cdT
h+QhWf5v9jXOCUwbdPZFcU1reWpNS/fmX1fJiIZjTTDarAdGw1+kKLjj4U67SP5MHu8oYKPjW/zZ
Pe2YQYEepJ1aMFSWsMVoA842OrHlW/MGFLqsVJnifGG+4NJu7j1L+172mBPN0vR3A2P2HP9PfzwZ
3tRpxGVgLRvDo8zhFjQosef8jxZbd/NF3bp+rCsJHx/2PHmnWf4GPnxs4ygTsevglsaqYD9oWrm7
MM1S7aIpD3DhnCDBI2QTQXdwVtCqAW/ujjyMM1FirPhmvperRsof4UuW2qs9Z7RC0gIpTnoVgJaG
7eJDSzd8BSLmnAQjV4Y22gRRZjj4wEYa5rykxKYFHlX4NSws3Q9GselaYAmqBgdbcNKggJL0vEAR
jYPF2XbiZinvCviagYByLWOQPCBXMh0/HD8SvPz+t42B0S904mkc1Z00R8tXYmAr/Uo1PI0r7f0n
6j9hCniqn9gss3TxNZXEMoYfo1Hmo1hAh3wIDPy73Fzp78J8t21ZfE6PLXv7GWeSy6sVIwbrUmtW
DA/nsk5lO9BMfvOnI6GZyDrNnf0tc3IKq8uXX3z9FiF28+FlIyaDxcs1+UqTyMkZoclcj94msudB
rVUvX6QhBXdJm1rLyG1NEoZq3Ib+MrQZYAHDs/0qUBC00fQNux/B6UIEghhiHc7C75f2GpMINOuf
5P+ULjodWA93JgFN2upg458SIl/m+wsPg1OYGkdvaxftm6Cyoz/IlLc2bZja+nOjDVYS224rxtBI
lsQ7pbhzQxj89NUwLsBGc11yBUxKK85PBs9fmzkN5J2edSPm0QtCFKanWWE3Vh6oYfssL6VanvLP
/pZmO++JcoVusiogVTyfwyvwJlBiXWR5YUbfTeng6zE23GilhC2sMJbsKolSXzCcrSzj1hHeiKbA
VEPjnOzupUGl5PjtbQoGD7rVVvHD3te1JSHX91rWoE1+bV6a5yG8nlVPHHBC1/AniCI06D2g75/Z
jINwthKa3lS9OceiFcfZzOAyG41nSf95ukuWYzVpx6EMJLJObw/iyl7hJKuCzg9zEVMLdT/3P/Lh
DgMhwvAJ7G5GijDMwMNfzFe49gLQKQjMxb/YD4B9ZVJwI1PScAOJNDcV8xIhibzr7HTMqO7RXX3P
yEgA5tGiwsOwzMj7Ha30AsTeXlePD/d9PZHmcywWWh65DbCRyqMUnuYj330HvBS07cDr1n7CvaH0
sIIxovj+Ts7G4Ge/IFA8vULX/oT+GuqyzUXSGe6vidWUty1AaoBoSmox/2B1WgakVtoHNJLr8h7o
lHzoJIfOpuhiKdzpUo9JBNasTrS33f1pDiaV1h79UeqtPl7lCrYD2ijOGgLbxyX973HJM/xtEs21
b0APt4EzAOdMN5OsFy+E9wT4pIAz5PYNSWX8PjfId9OvxabqmPRX6MG93TjsKLrOS73EfKV7dgmb
SUMlJsM/HX2tnjbqCd5Lyo3LPg0tJJAVaXmvswAFhJZod7XDV0c4po70y1Fyx9+JcjDmoCqB3oOV
nbzj+Yy0CzIOJfV59SSA3XkYFYEA/4Hdek8BZTiKKOE8gXxe7+15AxUdLaZyhQAMkcg+OQHDVe7V
me3QM6laWvKwHgpMvQselrklaDIHj8J57H1KN+mSFFoAn+U2vb4BLMcOml7chhwjyMglXFGk58Mj
J+WhVTDytmEei5/Jhdmm7bTKuWdgha0WOOavAlLEYnXhFms4coHtQ3K8Bn85Lp4fkawXhQZX5zlq
lEudpqPDqhgk1NJ535hmPBqANIdUow+AWb9nX5vQaJznN60/1BzuH3nYIQjG+pvahPdms/UwYvrO
nw+hdfRut5WqflOp+2ntOuqn7JYOIObExCsT+l9HZpXEpLcXRFA0qvuv9D+aPyKPOo7aPHpu7rXy
5cPFekIVqAbrJ84KONd5V6pvtVj4w4iVF6My3FvMIrPWDXfKD4lYRcFCFPA3mQYsdKOM9tXQa2cV
RsKwMnQ7YW/padfrPsyEVdPPkYK3TGeSBWjCISTiBlPzs3hoZKznNUY8lM+t05GIRIzs3lqyGtmI
LmZ4FGepD7PWqUUyttz6UHRIDhJlyDYf1lXNOvmj5SvMsyBLUKXNHHuILZ3yU/jU61yb7UvftJJ0
kt59rMitNEygNMcdmHfY0L76PoUEop4uVebTmZda4vH7WtVxUkZcKWNq4HGhx0lqqhqbNYuteHD8
J3E4wpjcOzkmZJdBadfxamtKbk0orfEex/K/LGEn9UfK7DCROnp0+mTKXlgwgGtYEmgT4tWOdBTo
svg2SohZ02Qe5tZQuT4NEYEP0OXtML7d/W4Su8xvuLll07bk5cD93Vr3ImR1RA9N2r2R4JKwSEtB
HeRqSp0UHoBbTW+j9dPXFYtoans8zW3rwu6XwBQya5LUWdOy8OA0fxsNhXHgvJIsAQ/YZmZ5oZxY
cX+zw2plpbRzzL9XTMVbqCKIIvADFBn/0NjyAaZYmnhHzt/IArsUMBgDOsBkmA4oPdQclM2VIoOs
UoRHCrUVQyrQIPEenCpaykCDXf45xczAUI5y01LEreHz8j8RPcRwyhRvExE9zfx9qNeIWmoDJ0G3
MwDG/OYSGjvHrEVhDMwA3UzDq4MzkczcjPnq7kfhc+xkbSP+LP+alDFn69zSjG+wlZv7NywipL5+
mLC85aohIZC8UuIPMAYrvOQrdY6K8BQ4nw8tpVN/k3dxYwbTn/BjjwSzqQPxYOC+65hXWFILjgNe
iYgAutmT+E4O6DPIuW88agQpLTqkavPL0fxdV1nAoDgJmcBbLGokV+APAMMTQxXeBkClP4hXxvdr
aSgRGh+FGAdbRmB62jP3dcQs7UYrp9gOLPeCOHvP7Ro10YpMm0p9KO6cwRI7c2OBJQ6DjakEG5A1
EULtitoM3Va+HmF1wv448GEqP6+9yWdMFZ85gJERO7ItYbbEuh5833kAbrk6oxFlYvCNlWGJbUaL
+xxQklZr2cTvfrl/hO6How4Imts2FxZGxae0yZhsj4BnInCWnIBbMQDUnN843EAtJtEDswnrtDqn
almLF8bCe6lypDufPTNTZ63ikYzskg38A0bGaoLKxALLhMMiAcplW7CPKNXVEaTNwCE9S6g8YH/G
EOHqkAmauNkE3vH1MOgaAXL7w/PzhScoK6MNIVf/PjubLGsyOC+dlazsxkLmrS2I5QJ7YqvA2DE1
yqDVaZlUOdaIB4Ov4Trfqsf+hnVGoL91wKsyrlZRlrwzD+Fi33A6/eNIvXbG5AqbwHOlWUuiQhPn
/D0K3BOgwarnrUbQS7ZG5gAS2k2YVvt4pfOkLceUhfmprxBma/sMBz+4X/4hFAi1SGlGzTPL5LIa
FX1DZ1P7SRsmGO+w4vkmCGIG08jDFxVPWxyj49iKSsQWFITvQXuLOD9IAgUCGaX4H/zuV05qJqUW
1qTpFq9ZmbS5vaHzgpQwp3bEuhdmH30xjydUYtUdDptKa37E2t/8hBw09tcbgdWgEZR2Cf0h6qLr
NSCTNYBZSDW+GzbBuZCEi8stv61y8AEdk7Tli2iL35mjj2Raalw2OF1WVewMhPhgSOECHArXswFO
+7rdqNZeVxuqHoPmrR2h/Otco1OR6VvGzQwAQcCveFMDpmYvSwYnHC2gZgj67vnWZgQYUcls5kwj
DyHWaNaCzdHXhDYHCvMJQSu9yy+WPx49LB+On1uCNFMGozQ71lfpz6SwcK5D89UhwCFtMsOWVRsx
mYdxtUna8Nm6Ice6hyV+N4QCS8R3jD1ciQdEzW1gDFvhrDv/Ri4owxF6amBgGqTxsMuH+spreCxF
fEiEi0q0Mxeyvy7aH21jpSSP5Xk41RnxyHECmBWy+z03fyumTo8vZsIQVuWS6lzaZtHa4A6xZ7xT
EfytX81mvkIDMY8v4WWkiegAYrjDh2dKdcb4nHOb+Na9c5AM3IemOfeKY78JOTzRjcfMlj1MDL4Q
HM3PVF/NtCwPVSw90j0bbl1te4IJjFHEfHMHRQh7RIAVipbFmfjh7kXDFnCMkQ0LxPSF5vUaLHtD
rNb1HCOajw9irG2vcb6JcanpiKt/WKyp8+6KA0JslXAe7fGYWucJQG53JPewLkSRoNCM7fzjn4U3
GVp5W19vxzr19ZX0Ih4Dze2HEgiS/xohx4I6G2Oi8njbiQC6bYWRtMFuMpOadZGvbw0By8TfjE0b
5TR+B/aOoaA6PyKHUnEmJqf2Yly3EDRIB/UuHtXgLQ49A90l4YvvlgdfNB3DtPDsDeECWuisjb/o
ptxtnnNs3a5zlzBPN4fCL/CkbCzUl8alcxVD2pPOOkVm8gCbQHNWlEwKmT5NERyFNN196mZgJdbs
SnMqN02S/2xoS2kz/kb1bPzYXxzASSn3WcQPKR6oX8ob8wdKF1rJ9+lEgYIxxao4F4xgqmH0C+i4
p+k0xUQW70pnCVWy8nm9z+Zd14E9FvSladJmffnASmx2BVhDVMbL6reELZFNp7SDpZTbaOJogQml
sOTptljQFmN3pzSmTKRRCqLQVuodXXK75OabfgIQ+3sOT6ZvgQrZwwbM0L0UNyrEwTLVSFYCc6hD
x8CN8qynatDNjR5sh4vIcPL/+yW6sro93RnzwuSiYCMJLaRk0rEtEwNoJx6B7C3vMK9pp9iXLnju
702ucPnNb86K3xPod8NxT7oKgykhT23hFUNE6BqDC3q2M+0OKzbxN6p17D8No1T68RlmzWgA8pKi
SoSAZZafYUNozTCTSYcv/iXuNeS7pCPfLHvFhGPnnQNXo+7hUfVzVD5EVcsQPoAuDG9ertRAHU+7
qNmQRHou6Y9riomopMVqJ4Y+f13Fo8SytPq8tylZhrza2Kataxbvem4e8hqYGUTUr4ybeB1MxTsX
wlPX6Fd+CBypONAqwcL+Vi86MxQWghaCxgljrEXllmRfd4CIRS8YrJFFu7jpqVPkQ9B+BtATOI6Q
LYwDhYKqJhKgWCTh0FUEABCzrYQ0R85NLlBOHED05g+q8G0LKw+Uym6zTyTEzl+F+M8CkjDZ02vK
95nTi16l4d/IiHZTYZxSdJfwPUdCBg4FXiY5rG9bXNwiMrI0tXEp1DVAwJY4EtFzZxm4RLZbfhg9
Vm118kL8pRV0w2ByRhMFI2F/vtbm2KzZUVX3WE6cB4iKzq+Jbo2kJ9edfw9LvibFkusa2mopGf0T
cUnGH6vOW+dH3vypMf4AuZHMhzV3qqmNSjqltuYRv5gGgcyeUraH3ILhzZ+BztyqnvvJO4I+hTbd
P1RqQKuPeQHzDM1S7RnDu+sQsr8rtMsUYeTE8vENMgrhi5vSXVMCu0aJ8zBhbe8PR8BnlQ8Y2Z5k
TFNmejW05skcU27MIVrqKZEAbpkx4EkQrj+ODkKl867jIb6Rbi2gGseTB5pCJdcUp+/05Z+it1L1
f4yJRwymTqAWWhd+/dYoEiZUgjmW5kClctGUu8sXNoF6zDLTF3XKioI3Q2uehgAwqQb+e8IMUM9t
hdG1DnxbyGLyM74CbJvjU1mvsDCT6xtC/C2+6fxXoDIbb0itJ5NB4i5mAQZ7tyWAIc5RlGMl9mTp
5rzyxgATdFqIJKVv5h675XfeRAHIi2pKOpV4KpX6rS0HtXC4eoP8DMhokfnk61r1kLUQMu4QPFYF
uJ5zLYTa4yp2CR5OTyIlidREzWRyPF4IatM9I6m738yyCk5+XDPJ8vveQ9Sdqt/KhLNXKPgbwUqT
vOVTD7sppuaweJIx2GwP5m8Fg5JUlP9u2awcq8rpG8oap3l09TmLtBAj5EapoLAmmtDjSGLBcF25
cpjUNKVBvBBsMrzgYt/gnhqaEsB5yuNSm1fNmVe8aXR8tPejHCsOj1ewv0Yzgh30J+Rn8FmJQKAo
jrpeO/4uQO6H6aGc0IdyGVT+Z7SojTGmjYPFdHomPB6RwrqEi/G6Zotj+VdjSCqzGWUVDNZdvIoV
E0oj8Mts6ippOItF3A4DVt05ZNnBfzqBf3Q3/ohIMQvGsvH0zHagwOEhK0fL1Wbv7seIQLOkaLhS
uLf/KS2bVsAV3VR9Zvlau7U/hXpqfI4SbCM3vW3rP8dtrd/HZKLMprogFK5SiafEdnrLoe1qHZMf
n6LJzyLdndvRqA3eBJ9ay4lGaymXg7LJ4O7gX0oudSk/HTBqgADB2sTLyUv+QWD/Gkk5v69ygR9o
VSmXQplzHnsh1vWSnQYoS0zmFHxE9t5xkqr1SsHoKLjBQNergJzWZ9g1e2ewZg72PPJJrfxAgkam
/oY1oo5d6waVVveTWr7rhEiDSWUc7/eRJ66DqXPl4ngKBpT712AqD6HOf723cEuOxvES5ik9MyxP
vq8rf4QBc/+fBIDzwHy42h/vmwfI+VptF4Bk+GfGpjcsgfh1e38XAYH2m7+T9UI7fiwneR40xC0Q
ulC7OEqBdxvef1uDSHc0ojrzKxNckhxUDtTUD/ncLF2w+xFHGw4ge39QX6wJLgkPj77UaGWwA1Q/
0pgaUae/WGOj3oGICg1EqHvWJSgjsV7JtgaanZQiVvL833KeVAsMSpkoPP4us9oC+/cHnZZLQBRU
p2szeHIzFzG4LfRNI5g73RzIy1wXw0+kCPU54b8SdVwOLkYGbP2iNbrvypfvuY/L1P6QOyxQXGFO
LlI+hCxwYhkZ5/jf5MeRmRZOHY61DK/2G/UuOwGGowZXRlltJ2LxHZLAdYHnWvWD8G2/TESARsC2
JLERUf4sgXYTU/aZ/mi2gGIpfZYlAzCNraWJxhqnyUoI274vn59pVoUvsDYOWKXfJKF9sVGd4t8z
/dAac0678+tGLkGlReheFchzlfXFKkfLLesS7XiMzpj/6N+3No8gJapI1zbfl12nxXbnC5ZqDhmN
VsUk5tdaeMnhjOlrVtupQltW/U/AJPqPjsMKJwx8DzNY8j4HIJoELIf3jqQGY1SxBoItkjmbGeuM
3HOp2spWHH6TuEvgzURfipQfDRTJLS0uhvkeaS3JJhYNVy/OQDrveiKYTMTBmTlRI849VV22+JAc
FQSRUFDI3yvp5zP8dy5SqrncmQauUJ4TfInltVwekHyox2ADnb7QyP/vr29cwrQa1oeuBioHNlSi
PU6UPFdJL51yNySsXmdL7/1VuGgsJFu5CpFQIPwUsUUphqiVDK6FDgWgBnPBrw0uqMxEDQDlD/xX
irTeHHtNVp/lkqxkZWjRBFTqQ77qoO22W3w5DwdlTI6+7ONYahSx3ESzfz1XSXR/YtZRRryF1igO
w+aVtnw6Lv/MNlLd8Sy77tIOMEQlq0hzK5U+1QItX2G2NvlG3NzsWqhnFllzzrvWDRrH/XqaMCCr
liflWwWkAXvceEZOze5Wsbz8BThMHSQfSqcd29UcX8F5T4oXLnfcJF1oli3RcI2XNhL/YnH39BHM
zF32Yc9CdnBkcMk4fg+e6JDEGZw6uq3/kdUBvhqcPbYOo2m3t7RreCJ2aM2bZ8MrkyVhtmauTZ4J
e3kM6mabz5nRFo5uxwT0wR6wV8E/JSkI6EJbt/ItAvbvIdcZoxj1ioQE36xjwXY2CHre0KeTRhr3
mLZ5MVzypRREvf/4jIxi6TNJ+MN3KmZtRtPTTTsKqhbfqVbx1S3sQugkAFp6QEKgjePCMYMUxyY6
rZT+7ncsd57f5B8690cPGcqDOBe1R1GsaSeBQLESvt85bBd16YeoNr1oJHfb53PWu0eLTlzFxvkC
Y9nKDBGh+YrxbDeJyUwtLe5Fh4H+TKrN2nyTtEW/RKaYEVZo0Y8k+eXsJPvEJZsDaIXI3i9AfCx6
rFp3gb6TvvCXVZSLtCK0lpwdAqoZrD+kfmT/jiLis5AN08HzF8511MBN8kYQr/YVDo6ELgGs77P9
rRY0oGMu+vVduqHk3S9hFdl2Xil9qLiUBo3JWRN2jsy5wk0Yz25+EmMBm7+143NwSayUzamN/OVV
vtu4PlQMr+n/0rBGbR1sQlUDCYLbNRvrVaQZY1gqKWzyNwSGRw+F9lWcoCgBaqxlslbumCe+Nfmv
28ib+g0lxxZpXLfEIXmo/pVjX/0LRUlGQcHNHubvS6ErIrWtnXKuetjG3Qbp/K1X4FF7sSlX9+vm
hVuPCnves2ykszwwTpPnhUVRcoaPbtFJCIqx3QfurLs9CKgd0t+XwD+ySCH2kH9ImcCZeDUYDHoA
kU+xF6rBX3Roh+pRIHH0ZTXyqZxTtfhLT1os3PeYYcej4++cpCAiq2cwiAzIqAxlEugE31i/GGM/
QrGT9v0WM6ZakRviopErU2GGZArXUKJInjzrDjeUTpr0fFneRnvvlDtRCgTlxOqKsY24TmIHRm2P
ZlSWNSV1OU76lShrMd6rsbzLhq+CC55HC1XpUczrgEC6yvd2VzoqlmdLBXhIILRoEMYNRonLNcgi
vtz0CZ1EPzvbrJ9v6tSTj6Ztu5oiTvVtIjuvoPiPS2neTqIwM1DxXyxlapnUwq5LKYH3mH2cGRGQ
L37o3jHlyOvJgogL/CuIlAejV+7yqk2iJcpJ4in7L+D1TYOMe/tEl2YBko+HyW7DhGy3rXYpWkFB
mGzhVTiMjWA5YZuSManOFuydl3sdHCTndphWKnr0tp0XslZSF5i7bLgTCgUNjEQi81BrIvO2LxIe
lE3/1reKi46aeCjMabDYxvNbqXvugRaI2vIcUIhfD9NfBEH2zp+MJhHBWP/TfUKQpNbl/SeTXqFd
a+b5q6TFufZFoTor2sXX/sh0pFj1r/SPo08qNSvkWOOx33Qha7AMw8oV4r/16fG4uM2/UDf0xtnW
DEHAoRA8C2TJGkuDiYTybJ4RX3TGMfkZRdCIn3CUequOeZrH/NhHBCBdNGhQZXKnqWlk2lu9uvlj
4Si/H4Xiy9za0a03bExY0hHXP9cv0b13LW+snMoHaOWKQZFg1fe27EmwA4iFtCBXvI6ZbdpGkC1n
+NK8i3S1lmWpzF8OjjoIIo02GsSJXsgnz0zeplFOM4nW7/4BUbvPjlowEigWu4Nz4VIeiFfK+IBq
UUPHQU4KOi/AJRXtqJKodZr/RXjSi6msKhOWcC7zdXjOn2Fg312Jls0iptZVB8JW5SMrur6dqQJT
vS8nFKJZcmIVa8e/dB5eOSrcTsXUjKVysLHqaOdFyb8wZZysd0h3EqHqoAt8QNsr5JMhMPLEFbHZ
ULHOUEGauZnzx8asXXzarNwNeePSsNE1HGuOIVVM3WCuO+ph4P/boDiW6vms/nXrUe4+FgCYjOCU
t4k93tFGFzcup4YF9KJs1Ke7xcEK3EcYKlXER0pnFltr4eTFSe0xFlUtvVpWf5UlPzPz8+F3m2bH
uDZjZP2WRc688TShKrQJI1JZrwh444AAOSbJYgyTrH1/2cGNYsFVST0GtwZ81KZyue+JkMTzpaci
6fwK12Dgh30cBBCTS+n0f4ots8PgOr3GOVoci1mxSbfv1TIdPqLko1ahUWiY7eBLp3zdEGrF6rzx
s7TVheyFX9JeKh43z6b/ep2GB5HaCh7MxWcEWU5pxQVC92eA4SPXWaL3YCC2TAFDpxrRuf+7ERbH
jqZHw1ihgGsYBXrIgnQ7+u6ikZr2XZ3I5Os5sqNwYUpOvUKbqsFgM1EU4PueEPSZVSHLfur1oGQ0
dtvQzIyhgX9dPEwhNn0G0bPsiJWUi6mCk/HBzZkfXRroKnAQ+GlnBwdBbjG4FyQGy3gSdeMKms1h
C9ybXBm4OSBpXM6Q3i+0157/W3M16FEZdXJInLgMFQk4tCg+3DMt/0tIvyBtLerTwzgJNMI4vS9x
2PulKLbIp0VPLeh/aagLQESYaH5ycyVaChZqvT1us5nKl9wIC5bzb+AWS5Iqfht8VPBdDt0vuH6r
TeAOpqpjcucdXGgH/6kHv+3y8v5Xw9YggRbTCX7yJeB8lHeO18YJO8VtZs7u++h1IVFbJa5S75y9
jmm9qUzHIZrWsDMGncLVWpaS0+x6DV5lAQxIR67yRXnrUhDiZc2gPJdgPTYCVId0L811psflVRcq
NlUgL6pVcbI3r22pUsxu7jHZFRGZDp77IWzukWX72OlYWWHGv3hqu4x4IDRoMPP/KTfWU3jcPGED
erKh4MaWbfkmShxS73r1RkxkiO1yfB3e9hKquDCuE6LAtB4KawfM1XLI963WmM0nMnrGDTI/rT8M
Wr02+9mB/kUIt4ZMF9tl8c9+nMOClT/LO5JbUXxNHIJ7Q0OfoQjydywU+XkAtkcjHWSegRFQif9B
DrbuV2XXoYznQz7ILa0/l6p9lyagUBBJOnlTqqhHT9NJjPQLHzABXq5igPw0F6mmRM+I0o6KSdtT
VJWdlmjJlmJxz5SnXfxRBgIjkNWJLyqyvuHCHXx428e9ABuVSim6S1JXa+XXHqZzZ6BFUcyrSEES
EhjxnF5G+yGNFm772aURJQlfVr6/HWMrntg6pcwpux+jI4hvw65pbfYBv7lhOhzlxyThq+u5DXV/
ALUCz4iLzM8AcTD8VnquKCdi1ILLWNh5gdsD2V5hHAdac+DAFNESi9j6a9ZlR8cjnvF+WM2iRPGI
qUbOrJa5zAAhZ95N3tPXm7sDHDrrfuYWoVy1Tv9g8aBWDjXKMgpz9EhFuIOqOnU4z/+34bzCeeqA
HbwP5H5+awwNMfMB2eAttOn/kS00L6X7ywQdMW5ATPhSSL3jOxtk1h7b0hqxoEbj6lFanA5WzdyI
q3GIOwgqWcoFhsutt13ev0lJCjQkm4rsr9fsHeaCUHRkCAnfsL4FuOm9iFmxY4M0eh2BIZevKenK
xk4Xjms3qGq23SLyaK8xG9dh0VR6PAAo0t8Iz6lXzBmIqk397/DPdvKKUuVlX7HqW9r8iQX0szEi
WaJvCF2VDwZiNA5Df0E+2yK/mpHcEkiR430FIxuXQin4lP9DrGlJnk0x9eNHhS6rBVJ3fkpXoEBh
aQv2Qig800QOKECL1Ski21p8lv6LnctCDCPzDE6h/nO0gbJX+QozqQu/YcvJC+Sq3MVyQwTQ/it0
pwcGKQF0wnMsVPnny2JwjYUJd8UWIkSlOFECB7tA596TgEHdao+DPlFdHSJO0EYmurbU6rKTdqe9
0k5TbvOlmmBLPq8YbCLQwOfa2VOew9FkURd0OSADfmNINhAAwc5xZ7fQbyxOmcUy9O8iiE0U/ci1
Z9dqWaMP1c9fBRMIuG+yzndf0nl/i1+Isw9AWsKwJYIAcsz3Yk3l8ufYY545nz7SPNr1ZjC/VugX
r5FbdObPDuY7WSTjWzz0ZiiFatXnrKxEqYYRzg+Zu9R6n3/2NCvwsPQEVxodNCNka1iXTxv4cPBc
nth3OhOQhlPywebSSXw65byr+wa5pFlgzadjx3JOEDZ3dRjd1ikVKpF9mrqL2fPz6RXIb00V46tv
omZNYhk5rLBhEYcI5A9WjLEczORtPjn0bfEpa+9DJ/HCfIiFLs39PRa1tHD8Rbh64uV5xn/m0JPV
bX8QbIyw2UeA1Ze0mVihmCLcGw8vH/5IgUtprVL0UCryQIH06sqYs8NXDHxlHY0ZPu334rw/Vu/g
Pa7mFi7Cl2KJ21gJbGBK/0RVSTslG+eMuTD34YXjdDaNs7GVjP3VVA+bsSGUJrphLC7en8C33U45
eI1iOg4rWG5cM+INQVIwMgbno5Ls6eqSfQDsW7SS9vt+Z5WRK2k7/HNjGz3mtEX0/V/IdNDGbcwF
NOwhDzuOfHgZXlrLriMJwgzwallpYjkc3Yz2Qdr5v6+EVXFsFr5OQwLDu1U1qofpvOgJUxA6inb2
vBx3u5JSFU/MrAOOcqGybGmT85Y3iegNsZtd+ud9iaEwCk1lmMs3ZHRR4PB7MxA5jEMsR6APHYbe
c9v+jAVHNWtT3XpIjR+ITucyBo7GN2u/xndPgPGtk0q9/484PPliupBreZAar2i8Xxgnh8pVmiE9
jcyRnZZMTHsmp0Vu14Dh3bjLzRPOwGzq5SNZNZ0JvP6sEsqhrhsE6tOPRi3CzDopC7WgqxAfroDq
tijDS14A1aO2EYikxW2uM7d0etSaUJd6jJxr67inxIDFTMoz/Jx2OHwslz6fE5yaqIFYGfYiYwKR
3H1z5eMZDkTuVlNEOqAg9Xm8WMni/LAJyAmjwfUMpUCzO/Mg4talswnYhsAsBVgSZby1SMPtWqqd
MUqnl1aPfZ5JKL0q067OIzWkm0Pos+zIP2fByA9HHzeHwvZxeSn69wIdKVOiy6qwTmL1x1FqsGG3
bsZX1yhpluTYVkz67xhQV+cJw/YMnDc1ks8+bt57I1UZWlKJxwTOLyFxHJOigMrBwLeSnP7o+Qhm
tbRL8sEBtEIajDZQZqlrUQ9Oqu7AxryNhBF10p7Z7tjpObvOTUnqncyVQ+Dg5MVBObq86lyXZE5k
tqbuDA5khf7ryBJio0hABBkY/PB8kVlkx9UDWMlalDsuyqNlmPfjmbWN+5PGJ8Fhceqoe6OqwoAW
JVpdeRdJvZQxiUizq/86kmqZHLb23LPgLWM4qLIc+BnWSC43bBDPCmx44WKahZxUUIKyR542rvz+
G04KvJaoX/OUiLoqGqcpUCi97NsDSk+3oPLFYS6poiI0j3Yqu7Op18t7Gy5IJbBtNkZD/Ltz8zv1
4fjfgwzL/64rY4TuUiUDu83QUHjCejLyvPGwhoht69W6zkGvmQjI+F8eI57V7qzus8XBWs88GNYV
I2di+8zxXQRQA3mr+hV0ePsOPZEd8+bKN49rOvNWu4PJNbS5Bd9JArb+rwRvO1rfxBdVqCCC+F8r
/25/5KUyIeJv5AE8bFOHrCT9ROqbbQ53L8WUyCzZwAVIXt4AM4AgC7UZ71Y4z+UDGYXmLyn0EAR5
RMO+LmN39lV0BtUTnt+JuMwF7Pwxjhsy3+f573p6lQ+WIdGd8lYK2ZLSNfFUhoQCCn0qRrSmNCu1
E6Hw6j1uQdIEIJ6JMAbKr9+8S1uv7Ep1JeIqmqC1liUvpwSb9wey3hHBkHgNrNzYAiqbbzVbQDgf
Go2Ted3ocUK7PjknTErmuhjNPplD5V7yTsBx/tM9BIdHB8UkpG4mZAez0vHZ/eFHBlfQFMdcvAvn
IHQ5Da3kbIvyWSJeiDabIKTupiE+F3vfYYawRl090vmIubwz1Ie1fPPu6Hp3ounG/t+uIxhadfVh
8bNyT8jMWL9MXiifSvnW3FIuyWbrx0390V0CuC2OVpwKdXbNLiA22/0UWeduwQzBLZ0HXOhKxZXI
dIexlC2w5Ov/IarhrVa5O6MwyfOi5d6SM22GM4HbjFoP98VorHCfpR7Bw/QXaX80q06zVkQAtgdU
ZY9CHjXswBhBw/sNYcfJKTAmrFQGpqahsiBw2JVt94BctwJG6DbLYMTa4kabHXzl2LZx11LqoJdk
to7cKfAzUo012GxL8q1j+nDDH9x5NKfRko5LjKkQk7Q0aNcnDz3BiT7GBIrXAPvJP/SzmHS/NlB0
xw1MQiFymsBgaCerUl20IcrAN/MZMYNpgWSHeBaE+904RDi6oG/VKvJOg2EZDII3YvDQUMROyZBq
oxZvndU6hOz+2slQtkm/dRKIZ/fQ41S60HaJyt/Zp4uJHNk3h7LkZQv4A9kfvI55BglWTkrFDJL8
uI21IaTkc3ujRMSM4G0lkSS+rCNcFds13V45Gy6FJ+/QLY37NxJbVrQl+cQUrh0+76BIrBhtU2ao
fI8+UdEWJEVWgPFJ19Qh+JpLj6bPUQq6iPrdKllfjp/CmfFLt3oSyhjI2gSjdU3+pMQeaCqeW/p2
/ffxZRyz5U29B0IPBlrUr2ThHmnzC9O20h4RRvbTvDld2x/t6EUAXDC1s9gvpNvpLrfUc8eghq0S
zdmupxjqptowmZX99OckgesCoc4tqDQ9kDw625N9KfvSIKIMnQv/l9/1i1ytlgAt666GHeuiY6PK
MTE/Uzh7lnTDUPCD/5us1WSHoQ6chHEca9KzpVRfuicvW0ZH7/7enebr7CMRTFbP2OwwkJdd2dUq
UrXQTr20DEBoj/Ncm+rORLODBZnj1CX9XBTh95AkTisCoc5rZcWdjnzRo9UY64NNN/6SjtR17U/Y
EP5rLfebvBUov/KktaqAwH+m/SrA5zBN7RGMcUY99t9qYW42mnFnZgHfgnNWg37C844tufF84B0s
2/TRI+xLgz9UKOaSXORQaj6F8QuqNZkKfpq5Hxqr2klhHmCYxwdVuvzZn8Xz65J84duEFjRzREq6
it8H0myiFsvC+WRtNHUU6SyPRXgXXplLQUpxvfe9na3MkYcfLe5FhsMEHvEjnXpIafwgm0eooCsP
kN80Z34X0k6H9z4htLudAWkm8RA00F09PExqNpfSRoFgU35VXD3DlS05IREjQ1OBC1SOr8MA5WF/
Y3ddkpdKaja0X0/8FmnkH/RXS/C+1T4mC9/QT3YdKdlhOOSUdFAYXRRjLFHamdhU00Y6a/Ps61ul
JH+jDA1Qv6zNAFoFrX3C9Q2LY4tI4Lkw/RKML5ouOtoewYR4d5KFUk0xHALRpO/3JRovJaywMbHO
Ow+X5TEwdbdRfwv+YP2XKm9cFykoia7/sG+uMz6rmDp3gGld5iUIvlrzEMDkcRHuNAzx4q/Wzz4f
w1RYul4ydajbZ6Cz3pqIRSgtMSdJSW3oXzsuHi3xBK5uFHlBOq8vbqvtYgPx4u3iZwh4GDsqjMaS
GJ5Lj0PVNZSjpCc9EP9WthCAv26YFo7xNtJUQuMCgJDpAI9mM44RAFQw8G7Xw6GMY424k2lflB4z
hqTJfo0RFN51s8twWPw7HFiTTcmTpICqZx0IaZJobBOxCi3E12/mUV3+/5zWLoF5Zf8YoLovO9RV
0dSPnSOE3XHPTYd7luOkNCBmiztBgsPBhYKkiBPuVJ7RPrfLOrlZZMMOAs/bs/5IAcv2fSwrC3A2
IxmyNrGgwh5U1J8DuxgvZSJlHtK/xojAWeLT/mx/CZstaFFQ/Lvr/fioLcdpbuHEuZ53PR2gufDW
xYcQpPT7h37gCEbG1E+oOi8NfBWpzpVtWFodDmZJofPGJ8XN+vC4vCiC92tBmr6orZ4n3FP/Fwc8
Pznwcn7gKBSdx3SRMnGKqYi2Lf/333cwCxTgHhGGq8K+4jRU8tVPrXVTXIz8BE7GB5jv/UVJCbO1
EyExIreI7oHpAzQAAZ+u1RP97olKcNT3FN2le5Mjw2eLf8uYUDPPL8ybZ1D0ih3GSRZR4NJJ1Wn+
hCXvegCibyqnriaOhMpDlSiEm9GinqDPhvbN7JJMzq60mqlrxDnEgHDKER9rs66qwXf5RqSvKrVP
YqLd+yMSJ9RZuqV6YBtyyiTWjSXEPBoQLYVx+uTcUmE4NYqfyDTPd7nvOfj6s4y+Hvvntgqxs+HU
hRz/u8HbKGnSuTPLkIdsJ1pmgiWwgo92PcklSbiGjNEqGXMiBbiFbIPUYFiJW3lazPekuJEKpI5l
2DUL91YdS3JR2SwRMQ/D7bSFPX3Twu5ouz+BlpU89bD0LB23FqgcoL2BrMvniysYNWy4LinkSqn8
PyaARdR/+Atp0dBlzWr6RuTzkXoyvsAp3qxawMAB6qzQPVadFUYSiuZIJlp2tCjJunZFqOoOB11E
Fl5aKF+kq70et33tXjgghq/RRjW/VhIVSjqDmN75u0zbGBmnOh7oCP0sxka50x7FMcxmaOjJBLWl
XjnlOAkk74/OnrQlxxAxgjK3faHKXfpudR5y+tb//Ay7Zmz2MuZbQ1sGwVNPQk8sLLxdzNF3wOkR
XW63cneiPsmktkSK6IyzN6b4A/+KwIsKFx/vt5QanX2KVRxKBlHyQiX5Otgj6EpQhc12MgrgNdIv
WiUDZOJwYDnCL4dQCKzgH3Tt5fmb3r8C2kaREkEYHMR9COzjqiwmsMFagG0riXnY7xesqgt02tQ0
V2xl3BGSq+dslLwcFdifJIGbvC8IwGyt9mJqGbx/B3YUs1c6L+EmcTZscKsSrqqgIYtGXugFyZ8u
XbmSbRhDg1/nPO4Xo+pM0yhiIWsvQB6lDRcs//7FSaL4yQF8UdOPgRNYifIESrRQ81+Vvou0qrWa
K6N0MD7E5mpeVCmbgCBEijPIU7O7cYsRrITxzeD5bAvSSCRi5m7aHh53lfi0Oz5p6LiR8uV20IFJ
hTF6kevYeWZqBvP9XzqKF2X1q599YAB+68TsiQMjzOFuuX9SFbqavopvzfcg308HPuT6ifI1OWKS
/hLx0ZhGVfn2U9SMsbke2LvqEOThX2ImTIzd8pnNcFxzsIVW6GrkOrmPNruzGmxqE5ntDXmdQd8S
XfqGEw8xJZ20onWDpv11w1M13CgmnVWfPEpg0xwN/97clptgZWONtAOpbN4f/HVWQd6LakmBtKGV
ahT3p6MP3D5BQavrcAVQjkjuOL0khm3qRXZHSaIHuYztjPCx2fNOeCHn1U+xJvrSf2qm0UHwC+La
GrzSwI6T9m3g+wgKKeKGKvpoYk6lchO3lgKnZ83uxES62VXEtLuaicNPENbCAVQ00wPMvHzl+XJ4
aTLN61yZEa0zwLL7z2vixQk+k+d1L1mmnGQmkzz2Z4+i04Fw3rhC39yXOD185G8v3JBYLsA25GS9
Mim2X4pVZ2VzpySN5lA2DUX2s+uefmlwI3fEJwaBPn8F/jvzj9CDzWW8dxwe5evinx1UwKmdj5l8
Zcpt105zsrWfGR8aIQNJtIP3+Du7XxmK1846R0bVDK8UCT2ihL1Y/AaC8WQi92+H3uLpEzZQ8XyZ
QVkaE19rA8gmUpJWK66M0aWtLjxSvT2hf12pgMJhhwKdkxNBfotHCupGv1Do/chy6GFWZma+4Z4c
/jonBsP3TOVVjlNp+epPqBvZRA0mdjMKyDGne3lxANBRC2a2xxJhOpoqny11FwhBfOUKMAlxDBbb
ikAgXd+bdq3XO4ICUWFo4X1s5rSQJv1NDyNiVw33haffP5fTs2CLmRNyTzXQtRf00wvx3faauM0m
v7f/x5BdQquoxuttPgqKWHDv8xuwQxW/gcuIkQD2E/6r+Yp96NzY83Y2QxI8O38ubjGWqkQ+sKM4
SgfnqKzF9OCS2R449/6B4DLktFb+xAUpQdZBShK+XoEzpn59Lo97AlElG1VTDv41On9KLQrHx14S
Jyp37NIH/W4G2owuSjJL0akzxcUaaQFGiNFe1+r2/cFlMT9lLzGmUh7GN+0SOFxEEpxP1WmoDOiM
TzebdKL+ESeORUgg/QsfJqKDlhbH7/FCbR4t0I3faU9TCz8g0nvYzCodby36F1yCbogVWYujTsjc
rRBojw8tvIfzH4aa+LOMCr3DPZKptWaO8vJr38GjwwsiC/cMn+W+30oOnH4v/1XxEm3pmtiFdKqg
lqjlXnCYuKc5WtfbY6dQnBdBZt67j+a0L4tya+1g6neyQSCrZ7aq0qHabZfGuNdKu/3ucY5reatv
gUiotBRQXNIhyVvlexkoscudhH8+VarOZth8j9pB3WyQDI8A28WBp6TwlCuIQj50MJjjyk66+nT/
Ieub6l+/iVUQZjXiNyFV7Wk1yA+CC4obqeDC4NzTE3A2OUJTMNfAqaiDfKDlgmU/RrQy88U4LmRY
1oVgO/WqHrHblHLl5I2A+Bze92Th4G3zhRcdiyeg//sqE0klKCiQgn+mLiGw39gYH1vCrQyhtkG+
9g8orDShk8GKbapYs4iVvx/zx8+cHl4xPP0Krigc2UVewcicPMRW3J6ph6sZZNr9Ul37Watzbl4g
h2tzXh3aEbvuRMfm7ICWQjk0qQufi3QnPfcUgftXuVcOOLad0HjbZy6TtgZkPodPzvVlA+eFLoRY
FYkS4LEBnzrTDJ1gZiPlQv6nGq43jCUYr3KoCvZQJ0rTlHhIY+tXcJpBy9Psk52BP8p7hjVKFAEy
9Vr6ItIHFDI9H+W40cviFGD69jKOdYd6fZw/UbquntOnOWN9GYGUiLvWvVJ9zgFgC10Dbf1GOmZe
+xE4Hu/u6HIxDQRJzBV2khZ12ZivPo1hDpopFAwdjs8E2VbeOXbo4pSCjNoTZ9wZ4aiXbg1EA5fU
REJRfTeaO0KJ0nf3YIi4t2lifaMbUOOfPCEyXmScID45mRbiBJZAv+hbiAQ2fIxZx/zr5FlpobVi
i9I23VhBi4Y5a144dEDqZlnS9wYCCl1r6PoukkHa8jnddBHH0R6vSm5WULCBHOHoBgYHp5i/2LVD
tWSZxOdP+9R36DpdRIqUUJWr7uPMsJyq+WDidypYlIUAsPs0pV8evKCrK5siJzZXQInY+EisAPHa
aGJ0UKTtfsGfUmmQwzEJmylRxC0XaRHIp0mG8wsTBwjeXbBhzEVKXgKRfFrSwQ1vik7UAsprvWN4
tPCenSAgpev9TEpQONVrSvy4Xq1gAThE+gXxgpfMaVfcC3HnhhVTSkBcY2+GLAcltSVem5gt3z21
34fN/zTNkytqf5d3X/cS2c/Ycf8+KMGdun3vYggxD4ZO88r614QAjhq/+08YHPtt5WHPniw8S4Ke
qub82DfTWy/xh2C6IgzC0XCqaSwMhsAfyaa+XRl4gZuL6uojtMfx3YDoQKWeGX2+sAOFmcuoDyNr
0sfeyDXh1TcTxrgTazo5D8wE8dvB46u6RQ/7ZuJesS0ky1gAM3wxJe5xxfw3eyOrIXp4eJJ5P9eU
Xi30oBxNenLWFCUaT+sCs6+hsfvwmYiSrYkcKO1LiShNVMhnDabEVbfqX8Jy29d4toOzhXsxtLGD
ly7AWc8EQtTvjRfjcVtlTo8ZoWNx7IR+rcV/iS5SsHKHBnf80diCY/Ce1gKH4E+xzhM4/FX512+X
i48HSEJXwhVzEzFvfnsW1te5Gb2D+0yG3KvDWDfVjQYMM06XrMrzUdtUjOt6eOHW7Gxyj3agqBTS
TC2Y+36yBHJRYekFUtzssKZz76BvrNlpnXHNh6xGgNRo0hwhJWxmgnCRuWxncZ0oGm3E6JtIFXnh
CXOEX8FgjjVdDN79xiSPi4WQOUDI74M0xW4hpu2yVXbtHTBBxN+opHoZC0kKHLzfvuNgmlbflus8
MxEUwiazuOMHfl/az2te2iuCyeHCLOdWaj/XCc/D9i9HG9MSa0QY2uMeHBd4HHzbDaVT6cxbzUSu
zgeTKn0CeFfj+dWyYBsYRRIFnXUGGJtsf+G7QcrKQUA9Pfaxsgkkn74IXRXkMa8C18lu2sdoB4zr
2bMIpBx1k3jXOP+LHjJzW9j0CW0LnDuw4Zth43kuRPydDfI+B2XnVeC0RGQARqGRZq3HKR3tFeIC
wUN9faNaM/kJ0GvjegvoOGVnJW580MDNCy0bQo1ThkY5/iG5P9Mw+kFLiJi9gLKdLGgn6fBOQu+z
EEB9IfcMsrAWw7UNkKWGRNBVPLr4FcZ63W9LbMOekFYllOeAbzqN8CmEG+VI6soxtjeF21d5Msel
qHvkST4rfa4tyRyjkhe+2qNYCcUoFTVQ4SjbfWeXqbgfd8r4C4LGNLa3nKLeGMknNStvXZBI6JVw
/iCzVacRTSsLfVX9y3KMjhnIVS5FLox3pRAB+cCnJsqZSCh6Kgi8w0Wr9NZq/2dzHqRlXFvqVZ8f
74epf5oqMrz57XT0muqODEVbFu8EZpWG6Imb48gxJvNFAeKSI14En7QGNDOgqaCCQNB0FfOEbOLA
szeGmQi0p96olcQLQiSnQR9yvfIbe99MnOh6GDvPWHTBf+kDPTEVYJqn0RsU216jhwfqILj+GpD2
7MdNaXPnQxwqcHp25HYozBDab4Ua92tIaZR+SiKgKfpw5yTz4VXhwaLDt+IEx+1Ujq7bqKQHG3lM
8bx3yZUJHn0wo4O4YQBQNJCR7SQ+rdvDPeKdjOFNn+EtbFSFcACtcOjHOFbDTVP5WdLuDL2q8TyV
g3REZNA3v7/u+DGuqetTxMFsbscROc3mvORJvsHZs4I/tNhu9Hcv7qB1KkQNqG7WPAgBmxgjbFVr
yVnEef1gk5WYKNxQ02UqCnqhQ0joOcgkDCbj0ZO0J+tgdpf2GzTsCkSMdI8hoNg1pIy6Ol3AlJTK
ofT7uLB6/XTuqOdcgMDhBMj9PN6+/9a/cf9KUW8lu/qeJ8SbZqkjyR8jlU35/XDXPDzVCgugMJya
B7unxrn9TQCMhj+cn6rCoOAKLgvgXU0CozU7G4oBfB7frzm4OwyyuLW7z0gVJPyKKeijOeP7YdAk
kpPEdJAMnOgXf2ExIXPVuzud9xr7++erA5F4+hCmrvCg5Nw4k5ceAFFy6dlW12McmStdcAcPETeH
s7oH8kpAEa55XoJTICS/n455dUXf9PIVn9xcj3gzHtvq4nhB1B4ZpLEszIIz6XwT/dUbTLhRfdHi
ow5DmHsO7C3nQOC3IrFTi4nfp5DWY2rVzyzVjexnZYZJrenH8QpK0kU3nOIkjvNcmPEj/lxzEs7e
rg5+EEzEJJaDgMhVSMvzdI4tNtZu8NeDg3BPgp+Ixm3dA9hH05EqzRAHA0HxK9uTaKIDZK6cxcR7
s+kB1ZbuUxp4B1M276zXMu2EyOwFWb0vt8rOiHc5bIh16Y3gvJEOjRYMsNWKu1QcmaxGJieyfljE
0pW/HRoi6R4ORJO7grPIniQKCpXwKj7eIVPm4KBPLTnvmird9dymUvSuTLPSsl3DnXdV1YRvxb+t
qSitBFb4gRquIwDT0uIzi58HGAXMQL0bVovBqFXJ0YNI1D0RPQMMznFbJJ0ueVOkmhrz6UQ3kkHR
3OfBNbBuIr2cTnCYCZSy+u2/LZtxm6I2oOMGi0W6E8Q8chCmjOBn8qY6HfjZ5W0aq5SDEVHOHAEG
aSjzINFAsdjxsbwB9/golOgmVo7NGXz3SAvh0ozDrcaLSRACcKkZOdBhb1H3jqIaPXnc9VPCglgY
+yO0RCHJxjHmfewE2tM3S9oEeRvKVojztjvu/ZeKccaKH2NzGmPw5XWOJYprL10AloZkXCyrkf0p
NRHygSyXv1Fn1F+WR0xLhfjbhsTVUcHu452AyzT1EIUFdz4CqZSOJb4lUGaHbNvtpTqI2PsgZYxK
HADGtp5BqsXT2KRijtUfqHWLJarZilcjQPLP066hXjQG4Oa1g7sl9XzAwRijBsDDVbUDd0cHXptT
0c7Lkvk2jH3OioiHzrQFD+ENDAYlUg0ijy0+gRGtTIkMhB+DjJIAR089OHPKU30OAp3o+0uQJJ7u
eIK+wr9HF1m7QaUHAPwUsUrCZfScmM3BeOfVsPjmUXNhQdN8yLI0s+tNLMvgqDI0BWg0mOcE0hLE
GqG2l9utK2yg0RpXzabwMbiriH0YtKt8hHK4Y7nbKEhiCorbg1TIflxJLelREuFYxUNmSzbs1uhm
oHZMCVleOdxraOyhaV86W+cchFWgGtsq63U8mjVOPrAYh7794k8Aw9lEqECCe5fmW50x0cgNnDmo
vx3UFNdsQ0jnfVE9ZBnzLTCIHfAmePI3FvhD571OdsYO89b1Bea0R2fJD+RXIOCkuAnCimtHco9I
r+dN8ZjJpqua4aj6HNoKZel4+GeQLxNMBVLGAuFF1cFcXHZHMtUKthkCzJk2Q4rgWUrAfOLS/NE7
JzqMlVDOhZMVvGib/8R3OStEJWKlNegszhGS1NSFaC/lTWTFwPRYnnfCeWx6Laf+bhxo/2NAecJv
3pmK+ZqBUShNWr1+InlylCae2YjxfpY29PUCt8td0mw9SGgskSrsiuf0/7ZNobULZSE+vkCgEKWB
RUfNusEL4sGfPzG9MIM21tit0FoOG/8Y/k6blcUPeoyQz13vOQSK/CS5eisid8qvLJfX3q3+a4Dm
MxyyGyng3FlgCJW7fTGtWRD+Bdn4iPWVVmqJ8N0weVXUbIbrEcIhpy9FyPk2NFHccUj9gBAhJKq0
Zu0dCGJ8Q6GRgUIgf4p5KiPQymrRb8U3Ty2VDpylu2iWor4ZoiVv5xLQYVWMXDeP6pQFW7Rb/gN4
qfypwVBv3G0V1wMKI7xUSmgToQ97wvugAmndSttrcJZGq8slNHhzbhj3lyX80i0H2BWa7aMbPhUo
rSC5KthgKU/OWfQWNX6ctc/lyLKASsYyEp/YKedjQ6/JF/u+w9UShuOzvHbkIXrgvZZPVdSaUagg
7P3o9nFFhFmEW1TxyEP88zqZ3pYx7yy1txZa8Zk2zVCOuWs8sakXW/+DZ+6EKXzJzmGKP6sfNdYc
G1G7qoJV94F4guEEUVxIbpBHu2OFb6eDu+ACb4z9kbApAVcKc8B3uF04smhB7fYi0lk65uYv5yNV
xClyKmJiB57Y4wY7PRu7e7sR0aBE7DHi2295YZAesXk3AOrzFZfi9QRvPKl9Mc9pQmwOjy82pmPE
XaeWz0aVs3deTfBDsqKBcI79XxLyrT5uaXJsw4RXQPMtdFelvlgBElRttMmVOrWeZcmnmZ70jWNL
zZi+FATAOvUQ2+4H9e5amJtoZyHCgBf5Ymxcm6L9WT0ioK2QaxEYo83Z2mb+1yI1bDrQV2Ym28DE
NFVZw0rl/q66cNsYACF+Vvzusi5Vyplh/uMr2Tr0fpUUNd2ezfuWfNLJ0UIHyHtRSAjLcmUQBBZj
oPe8r/cRLVlQqAOx9v4A9kPslsxsuYt+319t5NV2JWdmUcmxZhcaSeU/WCeFq9waOo9SJxlmmoDW
a67uv2wtc6IiNYrKsoOacl5LEKIDWcULJ85Crsr5U1oTkWxG6UoZnemziGQ6uFeX8T2SxHDne4VZ
hBPc9WLamiwkQGXQCLXdcS3pj6uoO3L8IniVjCBag3QGyJ6FleuwWCsEeeAIwQyI1UXW5/YSSyjU
qMtD/GzPKQyiYg/wTeli0ho24/zY1E9gFMwi7eSZFkmzd//JwAwIKa912RDyiNVkzD5j01rdbb5k
TVPiqzmQEnXuIqSqfFCm1j1P4EQzZ6J/B9lk6Tkm/qqFPARMNDQoygdwRSKri0Fl3YmrDRaJVftk
wSsVS+9p5zrRNS5M7g3PV6rerXYH+z1M2D+3uCZ/rTNrT3/Fc7auiozdni1JxxnkiaqwNwTbgMcs
Ntc2akm0+kIA2xW7p57xuXA51DCpxLerZ/7/e8+k78cC1l9GucZMfMHzfpJtOyKAdnsywruRmFDy
5SQnf4Vdk4tGoMn+JseyY3uIlK0/wSrZnQEMwtgM4HwiNjXa2xvP3+2ruBMP76Uxx9Kd83WHnHEO
e/NYT6N1Op8spQygFTeqXnuQKzs40IP1tKe4gLIrPv8m10BMPxLzAhHp7i93jekm9LR5ah0qLjsA
r+JBkO4LBYTUE0T0gQVwjAqgAc9vmygxMHzcdxZFI2PEQLLDHml/JgnyDj33cCbbxa4UzfdGrD8m
P6ate5wr9Jfb22TZlC2tUu2Qhcq7CJBSjVY02YVL0asiXXpWvTdsoGaHP5b6dcjFN6cEhOYaq1Ak
/fba99xX/PAWO8sHgtfobN13F3IvRmdcTd8vzlFx3eeahcYm0qzPApdGMfZQHwxBhdKPzmdum7WB
N0w23MzqveENYuGozD7pbwMBEhtlNVqHfOVyFoAkoV748O8qmj/Pi6PQWyIOAYTecQuy94cHFV+r
qEE+vahQbIvRw5nOHzUePE0Db0ETWhIqSBTcU0GCU4gv/4XQnWlgXtjkWkDN5HsAmqPG1cgWVtAL
RYcY+sxHY5m/PgDnfdnfdiBuKZwExWwhxxoV4ErCe/H75R5M1/YiIVqEEQvL44D0+0AFtwjK+V9e
b1DgPDEB1R8Z630oPC7qlDCRaebTpEyzmXQw365F35+rHZyvckmKfxO2BpovtPj/D3h8N+6Lf2Np
G7HmxtlAVmdkE0Fg1liJdWciQ7e8TTtDqBGhvoH6FPtdZg/yr9wPMgNNvNPLPjYwzM8S8oJ7Jdqw
vtAMeC6eXJ5QVZabVP4LVq30AOPf7AjCTZIggr06DurlWqIAv9NiUylryV7ji/V5xqlMTtvMMizj
yvoWaxPNNC+tBMj6+hk5iTDmy7VqqHAUWtMRvvjAg9vkVPyibdzKa4PEd5KAGNGSF8+le9y+Ar65
UR5XESr6kNp5Zf6WvlimThdFel7QJ32vK4YAKsg782QxC1cc4Vo3B1LZz9+5++Seipj88UJpquDR
zYzpv0T9dZEqGLbKVQqJU22/g6HhKeDX07S/3oRgPwUnNYTkR3yAuZqGbZjtg8ow/gwTRnPFTmob
D9tW8h54oqPW22CRv7dz0jS916yNKfl44R99EQOay7eY88pSAzf7LgUh+IxcxA4LwLMXW0zni/j3
qUnMh5zXecPJoFCx0dmD6J+jCk/i3pZWIa54UJ9Oa6x8gaJhHHwXIBuUjzn8mScfU2FJNKJnOd6K
aDTRAhYqPckpSoUjn9juIlURPoXW0/PuS1iSig9PJhRUyJY/7rphNLBezRCTe8XSgxFf1sXkmJBO
ctnYH/8GygsBZuNL7F9XX1VbiPGGu9EUEcGopPh2YW1l7Mv1B19lUn052ZrGVesSOdUkCweeQHEx
Wq0ZzBy4rgltSX2ccmzv9fhEv402IsNqW4Qmt3gV/jN/+OcQHSrWoa0AO4IILMegwpXnfyGZpgWU
fsRJx2myxpC8DOFxSV9yEZAAjsGy+n39Z3vDMzT8xR1gL0Bug9qCJ6GNVYUS054ujgSWAvEnGab3
69zT2yh3b6vCIUGcYBCkCiHeu8StkE/Cs08ghh9hWGXhLkwar/1Q/aeY9py0MsjbxB2R7uOoJYM7
jpaKBZO0nBgjXZQfnmrCuVjHKgalXhyE41RrwX+j72Iof6In0Wjdcd4GNY2qxmoRYM40J2koIBtY
oenvGtD6zjodTYO3mLH9jol9X/qsrkyZtjpfcubVgu3ZI873vpbvTIeWoUUWjNcumuCr3C2rbj/m
cd3dpmBrPIci0HEMx7C7gQ1k8C9PEmW97VWdUaPDWoh6CS5XW5Moy/SfxbElK+vsuGcRajA8rPTC
hwGkgw9XLLB+d5AisUeXdqIkR5WCelCZTmvyyiNziBbB/OISsQvcUOK2vFSZ/D3IDA21AHoiuXB2
lHMRCmOuH5C4+WqROr9M9pSg9q1u6QChLIVebqETLXx6FUmdYfDDjvrIujRBqk5evv9dK+OSirvK
/tc/MdeEl12Tzxf9QbzfmtDSHq94C1+wmY2/A2h0QoB9tfTZ5BYvoFwXL2UPzD4R5MOsX7cNvWW9
f4SkibExtKbd8ie3V3yPdkd3b85T+agmHK4LTIxozBkzDxiS5I7bMl3yAUStQHucu2/20OE7cvBe
RFxr5Fcd1OzqQNgLDQErtiyOd7y93rYaWXHZ8DPeQwoMZoa0jzokBp6+L+nWR5OuhY5sk0Nkghm9
ZbAO0vf64iVulH33z0I+Md+KYHoGOGwpmGT5kzHkmlkqFkh8+XkjIx/5TOPGQCtyFcEBp0ArEdzK
q0ssGvEFpOrvLMVnDxUBGACGgb5ms7pUxZPYxXBFJBv4toy7L1NZpJ2ZfZy2A2Y7gcIksNLQNosB
73Vq1kNsA0qKhdEU/17cqBC45JiEBCQyxev5g198nluksIFDsZ1rXDw/FqE7e8nr8AjxCYXVRDS2
El1dMMKCLXawK1zSLAzpt3lBEL6dshDz8rU71M2PFujLiClWRAN8qGen3tzDSusAzdHbgdTubPBK
7AtGUjncAp/v/7UPZDNvRQZugTB7uAytXSrFQUEM2vmhvumHvgYi5zyzNPTapP0bhDjw+aodNqrK
Iolmh1MRHRT4G/ei+qy0i5SuaTrEMqzswEeWO5WvjM7vhJ6PFF/w0tpmWZyfXLoZKUwHAiwlNsBF
6x6QNPi4HTzluBM6+fTIL9K5cr/zj/cYWg2SmVFVcj6DAAB87Amyrq9zn+u1QOnpVXD/N+kBvyg6
W9sfddDInk+CQ+2QNLJyEb/7pa1SNZL7D7TN2DoYZEZGoFNYsfDdHvC71W0Yajs7xbPF8pdeb7L8
rctPI7j5+LnxKt9y15rP0bKihff1KTzi8t5FqMrwFCgKcmhrID+Qn+b1iUp2ASBnXVN0l2euQbAL
sTiETyLH2gtiu2EAPB2o8NTzRomyg5lrigcO4nXALc3J+K7sd0xBeQNzoo6dDEg7MeFacCdYZuO5
1E5jci8j6zr/op8yXl/N2rRt2jzXqelVytc12YU/Dn8onegFL5mHIAE9bO2HpSa4bTr7EZ7WMHIR
R6DSdq9bPxGnYNmcwoibYFLx9e3ib7gi3vXdi+OsRHKxHJpLdhjVsvj2GQxwNLC/6mWr9R1xD9o1
fOQMori8LjDAIaxXMkxrS17MJA6WeWk1hucJj3AhlHIMbSLbJ7pDnbbgAynod4/enAiyk0niq/r7
AYgwIkcbDLa/g4vh5kxLUnujGfNRnuveG4dqBY/YajQeCz+FbcB91NcrtiUDVqTeH7anN21asfZL
4KCNm0zDy1L2IK9RQqMoCWFkAW8TP59BWtMA3yD/P244ET5gYhxpaKoz5ujYrGGjSCYeabjzS5kb
5KzPL1vp6Yrl1Ox2115HCB0SPFKAXKQGiAP9p2V62a1slo5vGx98++m+TNnFrXloMRhOVVhFiCJP
BjqlpBl/NzCOEiuT+eKVj4nR4FNTbMZAG5p6gd8DYZDMnjvGJKPBuoWuA/nEl6jtDPVquDQ7M/jn
qhoBqARjmLsxlu7r6hYCnMV42GlxWAiF6TNFkzmuBeoIDwDVR9YMndexAeV6MRgOrieRU9UyimxG
6L0GI9yRmH8T+DXjhHuTON7z7h7tBptdnC7Q7K+eliiVPpq0ik85EQbhuEgX9aY+rdfq7oSnyqsD
XpqmBa7jD/JAqWBZZFwgLaPi2T5/dL8r8o1mapB+cLgauRfPvDPyzZXGWs6MsaIZGAqO1+80I47W
ebOQORiSqFoubQIafooKXSdfdZECkgg4JX04l4MSg/mdOODAA07fZLLJpRo8nKKTE/ti8/C+EBXZ
2w/B9Jgo6EJ9UAYm/Pen8gLBadxdxYp574bPg/yWccAGAQTyiTNsH/SR3NQuOn4RDvd+UnpYZRwG
8Li8IGcWdHymlmL2BzRYQLR4NdxhN/1unoH4V1I8ml3Doof3oR1AUnuSXL1ovAkY/clnRRjhDcD6
sb3L24AR1Hr6hBEL8dgS4HBwhONQQCRu9nTji6S1T7sNadh8nRKHJkBFDULiLRI+/8NaPlVFd8mj
ADfwfQxE8j5I6p9RJx4DBvisfULZSgdZFX8VxJw4DZYUq7+mreIivcTSbGFrRHZi8Ge+YblpLaWJ
2HYBZyOKYKK/9/5b0NFu08oYJAUiPYADnap7l7Hm/90+VUnXHiMb9xQaiv+Cn5I3jAq/+S/9iQd/
4PDogD1J4zqwz9CZxLKPBTpLBEjfc59t4ls+lc95Zgpyeo2HWKBi+H7GjNHbNheSlUylByCoq1CR
TfJuzQVD+RX3fw/jr4OV5w3sgzwO405qk11nTH3TuvC2WQ6HJrz3nih5kj1Mic8uH6pWgkvU5AQt
fWB8KLFkTwApI12toLjv6lX7ssC4tAp0bOiK2cGLOzlAfk3dW+5ATq5dd45AWW1rNWgPeagXOxGB
lXCHUGbUkVvuPB4jyRlguMxGztYHn5UzcTi0ypgbX5luw71G0gU3mjhLrLtn4fRKwRXFiUT1gecn
jqXDw609azS3v37Wdda8ytguqP6GJBUfE4l+Q1ZQTYtQ+2UTjxqBASMhPZr5d+GdfuhWnSOy1W2J
rOIdLCxC8adVRu5RwIIPt6eKnevKjUcl2hFDoK5C25GSUm1KTFtKq5DKYS+fs3wJyjxivRrmKprS
jgtObsXmE3K1xdrSMSz4Al0surZtKD67oOUvwXh978/Ealo4OHpPwTsvTZBYk0JcX8/mmGbO0if1
n+UqB9tYKsN/HE4nRWCauQbm0Ef7ob+ZhImLIzuOi2h/WjbOaFrzKIyNPxwpxMp6BqlhUEv094dE
+cTiyqGiKAvwMmazxSxEmzWxELBGJotrZyxqxW5RMhjPjg6Wr35FYGmFHxgKDIuFSfT0SMp/ADy1
5nqRy3btNsq0lv2dlO16/OecPmYEG/BU53Lw7grzExZeADmWCf5Nbbrvp8rrkwAS655aoG6TrLua
hBKe93P+5bSMKLrDU3xyfKmhquni/1BRdVVZGcZMCjOvW2fiRLczWYDUq+VIfx7TFKZm1hGfYopT
9zsAg5ilbr2n6On4lzbGGLunc/Lq1ZRfnO4Vc7om+hgG0bdbsFxAclEmBaDhEgx1JQD5zX/g7MRq
jna4CNblSbDSKadUBQcEnp/T/zMt+m4ntnnQYxKjgFgTWeli1jE9OFCvaDDpD+AaEI5rBQUTDkay
RQ+2lyxDbIiCM+Tp/eF8D30fP23oTS7EMY2XVu0We9Ivp/P3coTjVAG6CL6tc5H3wJ2/GsarjbC1
+bdr/lprMMn7af4ID1M3jI/AfZfiW5/9tM6Csa/zH0jqXxbCAkCTyO7rdO7iA1dE+vcrq5AfqaDO
t1pkgFGsQ71MVAwGM1OqEv1lNu3SftwVgWnxplv8oOB09jViSjCxdVhTZaKuy3wy3UdSDRBw+SwF
4XDM76qt8LVRrMIN37JiJOP5K4V+hOx7ddJ4mClL91uHARlemmmTox/sB+fjr2w7+tNkz6+T5gWM
wJYUaZufdGTOatMgVPlH2v8WLLnJ5TTHuYTXTQZVfOZu3MALRddl3lMfIb59ORlgrUMOJAnDG7v1
XeVWNvhoRnhncYEJu4imYf7JhWEs80nGuSQjqnBXFC5fUNdnB9Y00LUf4sxKMhMb/uCuHfdS4Qne
aDxVrFeXppi52r/Ae7ln5MXq+y3MNDOR6OZAIMfr0nxwYi4mNHGxn5kI8n2n0KGzJfzJT+8+gmlP
olpmDRLIepl4xW6/tCLJZEYSEftFsifkaVz19vEy5jjAeb2LIB7Bty0oOVZuAqhNetUrhvAeR/FH
I+DKynibDAFamXUbM3Ewwemvq8d9naP5SeJKvCwaZ7IpKkl+a/SZtp0kjBxKGN0KWsil2wZftO52
/CuSpZmZAppozMQPzFCR0e9zFmLJNsLVgACcUCWzB4hqxIWtp9hpvQATuvlsCjeO2WuBoRgOj3xS
Kt0zpLErH5hJjDCSmbNSnhfnFkwji8Uy+zuLgf5yax1y+1eP+KB5CNbpfGxthirNbbl2sQH1SCXo
8RVYYweukA+z/O52GolvRTF77dn0e4Lu+9fPGjakJDJrHiyJL2RgTRjKZj8x8+ljOJapF2W/hkm9
aMR7jknqWqEuq8V30VYYAMSHnk3ILaIQ1jx9AhRMxV/iTKf1nbfyEu1dhPBw2suvCuaGUK14yNB/
wgQH2TInIXK2cyfwiSGwR5knF9CsUVYmc3RGFZrx/kOkAIeeiixvsMtoG0/264QnN0Xm9QxQh3cG
2Xv9dTYp4mqF+gvJ43vMYwuCsSKiJZpJlusRsJmZKwhxNE3X5PkxjAK0Q4fElkoxIdBAnBkmaeqB
JWUVti9N65D9xAxl3ip0fuYR5tC3GGeHANSC+5IRGIOtpxH7PJPF0ReLAi4eaonNjmWoaz6gjlNV
sYu5FdIyV00xZBrlXI0kMxFjUJy6tnLgLp0+Lg40UwEukKuC6pNWKpnTLUGjs0P8GwYt4cNVTyMj
+DIOsEwkxEestixVKVHpwJFGWbNB6nLqt73TCU65jiyWu2xsZacR1qzFCDH94CNcGAtKpYiCZb0C
1mcoW10rdBKGf1y5KtO/Sz5PoVhtefZf3pGAGBfditOLNJLtvKwqZq6baOkzLAf5d4Tx+JmaJKhz
bM1vY72miph4X14RJZhXQmljbvb6CDOL5ws64YoG4+MMDDOmx9nGnayPgUpLN6s/yrJQHaJzm9rr
EKl/74IxtPJo2v/96XHNOo0q0djS8qSfPnqoZGZ1Q3bvdrmSTAyI2eqp6zy4U2DY0w79EL7HYHzF
iHUcdwKrqe9y5bN2Ar0y4hbxtDIncpewShWHQj6/IHtpQNT6exKwtvMd22RdsnL2Cb4svl8EKawK
Ive1/p50xwCr2ekNUIjmIzx8/W07FX7oFxH/Y2O6B0ELd00yKEdfMIxfBYMYi+6dc/YZDISsWneF
INL9xnGiIO5ydddXQhZgQAXltQ9DmKjecN9/pk9usBqTNqmStZ5WeeTSEQ9UdOq3G00zegA8hSmE
koTeRGZFvtVuv5vRoaHhZ9WU7qf314fKzirtwhbCNs6wG3wIBrCni12IbSGVfnbr4XXtI7+K8UrI
NVQRQTKeDetVfM1YboYpwLmJYTpu7piyyhAu0VBkMCwK0h80WIq0BgLStmrOofnXewwPVJ9laryC
b4nBGA8/gs4PElpP1sTJXzG5jY+rqdRYGGLkDp00YpFVW62BrZ2zSkfN6YwPNXMIqd+5fRUf7Bft
0114oTKHwGQo0Ucem/lnBpSohD1RQ9YCJm7dU69RoY8vRIC6suUJkS2NTOXZ7h+VjdsVMqy6AXgM
Q1QwuR5rQHZnNjhYcbbp5WCktZunXkqsmln/2/OeVKtSHJqeIDzXa4+LUHp1LvT/T3MP7S6nXBIh
EHx/CGAdiM9CcweL6Opr8yS+JubK3YOwC7VFJzYg+5jd7CN0eeQJ3Or+lc0O8mGhZA2v55wxeREe
TbFRzyFMtGmA18EB4WBgcb81o78ZxMz5W7xYcNiJQpiySyJE490NSd1BKmHCD4/TG/XnLKVYdeoq
HmcVzzf9jZA7R+6WBvvtrCWC426GJ3WH4PbnEk3p6lH8I60SyguKWvCgny0tqgrXTbNDSHH4A/9i
pOtQrksjOdsbQRc0Qkl6663rZ26xvTGtHj4bC3M2+tOEM6xAkgheoLfp4XD1LD7Z8u7C38rDnI+r
opG0FwjwghBooo0LcKFn0APIjQDRC1BvSp/8lk2Y7rXrqU/f6L0zQoB8gCM43jMrYB9j9WnbNjuL
u5hmSsyb8hgeN5OAqOr8UlepmP0AP5nZX8OMNGwCfG7Aj5/V1uPsYtLprZrISobmwCOJMOsg27d3
Ex1W8Uz7bWEWrZn9i+jhHhqPyOMiBluox8W/n6bRjD5es9Z7oVnLpXREAhVcHvRxUFDomTPpBP8y
6Z+5jwF0Xv0BFwT9Nb9QYqNUkcGYGqXGTCWDEBZcpwCQald1rPoRL/THisdrxGIv0VZbcZiBHXHZ
G9l1PnOydrsmQ/VtCYCH6b24bJzaxubSMX01y0vHZoGPJPkUTyIEHYOV9Q4wacYYWtScomoaRE1J
UOs/Vb1sYwCT0DU2ZRLVcWKPgrVCBNMS2yLEzAqhZbHPL1HznrH43v/pAOLbTUeOufuo39qOSuY9
mXl6mhDzPybAdiZ5y7eV8eKvQyu7Wt6c/Pa81lh7Yxb+z/3nzKGaHtLfDwL7wokp5lTTDwsZblR4
ajBuwR+GTKlzglzLv6fY+jjSJBZpyg9QW8u+JFuWYxGxEt8gyAz/6CgQN9o8myCSLYg1c9L2g4Fm
Eijii/KEqkf6OqpqNpAL5vviPylb3Hvr6N0teLZ6dDSoSsH7Omi7egXQrH0fZhksZxw3ozEaAJDm
hPuyPw9Qg2RpNjF6WAxAx6m6xVCxRKxWY7PNTZKCeROCitcbDcL1smfV2m55D5zM7MvrvV+EolfG
OosE3mp+nD8FSsYFfTv/ecmVi8XlfgnAxpIrVpqBGbCwfluFacIQVS3U3cu5Eav2HfJvdXfqQS66
SP4xqpPbSuFTi0FDL+YJkDlx0aIrzsjQ7zNsfO03sjvpc1N1k9zDt/oIBODPkgPYaz3io7MiRBIE
2esr5RjNS7yQYHoRetrqHP/ztDCu3Vgz4uBbbyP/unCe0Ey55mop76JEwvJxadtGKKyyFOwe1GSw
6krPWj/0V7Xaq0MMqeoqwy/2DQM+58SHGE7XTQnjvMJaQa6bV6u+5pdHzjSfHGEziYl43eWnuSLY
PwLY6+lmDJjZBoPd/eYtqLHi1N3TM4NQf3Hkb3d03ReADqX2t/OeQWPmFumcX+RVo+l0N8/jC5jA
xFz66cNCMhi6mDjNUpk4IqiGHOCKONGlLUS7ajzJHjigU5cdiixCdilog65qknklq9a/mKmBECIw
eytQH731Zr7TPoZgXWLDdPYu/vtaEYbvbzdknfamc7xirHB2qosqX+Rn8Xb+3EJMGMOlpNtU80Ki
EIhQEbEX5WF/hM0WpI8/rNgbPMxiWzBxkxfPDqknrCUVGwJlZrEefOoo9tnWF4/mv0iQZdxaMf0i
8aXYF+GF4qbmib56GWXiAz9+tQzWVwKX67pYOwQT3cdPnV80ujqvoYmwfrj0ZNNmFH2hazm64DX5
xWYpNGo2Y979HBrQX6DpOSt91xV2weYXpLuwxWfDtZLsLfunaRBRzdfj2xHioBam/LOahsg3kWJ/
YPHGWXG93Ym20t0mMM+QZecq0ZbnntS9fE3s+yx1AiBgSWa2p3SzhAOjNoskEAAIB5eMi2Ni+aUh
dD3f/0JxJZH718GYJWtghOya0OQAMNeGZ6tGXMQcN5AvKLmsZNx5VKatdyEDcF7zLogSTBmpXJlg
jI63AdAueCtx9RIKtp6JQ1VdERrXU1Zx4o2H8O+1UZzEIhC+lZnN6Zi7w5a3e1vny1KR65QGAdpv
rR6kN6p2Vr74i4RIQRaaeWCr1ym6yXdhK2liZ9zNR8v2n49rSBprsoOMWC4Q6Xxu9Sh+SlD8W8Sh
eq8sbm/xtUuEkXkvy84JeCct7L5D2m8W18o0QzRR3zDNLAQBvnNGH1aDQG7HWbN9/JT+qAaL74Qw
0Y6jaZfa8lLCxMKUlBW5jRqTbwCklBwMocgf5m9fuH8tx4KcqrIYEsO3cgSLMM+OlPfAkEUvLveX
nfDfnK6+V2mJn+PvG0iDlLKONSwJugVvAwO8xq+XrHDt9g9YWBISwkHAFr1jR3hd3008NcWRVp6U
wqS1y3pwqM0LlK4LTdPbq96gUSZzfMJOJMNvBL1TvJYW5CAptKAzEaQfx5+j98froYxk1mP6QGDu
Ac7295S3u91UwsBhkoTNGTwXBjh6r7PE9dikCMOas1ZtttDFF6oiYFFa5b246pmbk4wIcrY/yLR0
20XYJvxHECM4VNsrmLvx3udnp9NnFCgFamGhOp7pdPAkP9FzlNnkhdaIuKSqwGWNGZAuKX6LzTx9
RRk8K6MS9GVmmavKp3mcTGRxXvSuosapBAMhy1F9F2twTUS7n2ply9VwfrmWg6GDJWM5PKC5CQq1
AUSq3Cf/EcZonuKlsxoEQI8Cch0pTw5cIG+R22MXPcErZ2JBCfKf3rnXxXmTarFAWKhrTPTVof9J
eiszabPGKtbZMCk2TKqZSZ9v1A8chZGbsD0gxtxVsOFcpoCjb4pTPjGH+jR66OdnSvmnpVtwrW7v
a0HalH3mjttL6fspobC/rnFDxUQmZYV1vxSwIIfmc/gD8NskqRhWFMlZt0eUJoAFifpUosRJMtuC
QY8CMFh2hs2DfFjU9i4VB/BUD604bBgGAYEJRJnDcCK5d440uIzWqKbcKIeadZeC+SI+AkVB/4UX
HJdDW9OpaJ7t/ha9YJ2pOmmhdPwDUJ8t9akGNFqiQ6xZp9wgV1OJEFeDyr+riicp9eVho4C+hEnc
AoSeRXatOAbSUrGUZcY3jjD8Wzdao9Ze40n3VG3VR5jAy0Sdphbp4kUsKRj3HJgP/01hbX+z3a6M
iUM651g7FFUZ0QwzN1si4qgrSrPv0pa4K50srAmrseLt3g4zzLmvc3WcvF5Dl/BhfGR51V1vmwXm
jJDkr75oUU3cVKJ7DiZUonCLlV4RD9IN1XPrjNqlJuMSZnfuzCGuNm9b8jjb2WbKdejHudaKYTkY
4dxqZ9w6G16J39u8zX4WaN6aZXaC/efwihwKsvb/cZxMBLEQ+2H97AGxJZQYcANWOC6pwQ6iX+F7
8kiHSB3wVHr3CDnpOLb4HUHS5g6DFZ35AuMbBmd07SYsuwe6EeM7oChrIhEZz1E7Qvj68P3+0K9B
TG5GUEVHNYmK0WhBDVipUHsF6LerZVIjFkCBfyjLWTRRL/sNuU2MeEdRcsNL2UAfLWPB+rTFQUV4
UECZYxmob9s4c5KlTD4/p3GAD3eFgw+qdNCqJnKT7iUvWfZN2yRj9v/jz4yvwVjEAHaTN96Agtht
ut62lNJobaqJBjJaef2lQ+QzQY3NOK7v7ZgXTAeXVPkP8mCTU4wT3M2bW//02zeY03h13TfgBzfL
EkQvT+EnEYJ8nKk4Dxcd7jkiB7B/fu2F47YtCFHwmM2Filb261s90K0FQ79XfKwDXWWQV2Z14tO6
G2hAPb7plHSQE4nepDz0xfvZxI9uZPN7xLiMRkBbVSYrmlPMEN+esLnz7tOFhsWwPe5g65eDRjw2
V7c0JuUJ8kDMWhXeAOKkqZagCxQpmqnQsJu79cKfXijXK1qhX89FI+gDLbDVt672WCTu3ElVO2Va
8jZJOdN6Lk5ZNZC7E29xNKvsDoIlvgnbIPnNpDoUTUigMT4yF+1dmMkXGEoP7szwFnVwKo+t7/qs
oN46T25zcO/AtCJEImrG2C7rryqdpXLAOK7DXR0Ug6XFj2zK4Kemko4Q3KERX7ANwI3CBcP5Z6qW
Vf2MLLjQyqs5NBQI9GcboDsdw2Vp4ycEl71anJIoMpzbdFUvRJrmF4+uuRHhNjA3g3gffwfDzqVs
sMUpN6ARXO8htcksYCmqEv6KXN4a1w8sdrQp923bdzC4auHCCX8lDndb0FFUH0wztLHcUSwp3Wyx
SQS7Zc/8hOFuJHpAgBjMcCZTblZRyIPlr0JwPax2dXkjJAearUpYhqqqwu4wiJkbQePMCyyRJJ1s
j+Q+YjWt0QfiF+6rbSX1GR6RSM0d309xCqqVhnxgsNBl+xnHp5YaQjkQXL17Hmg6XCotZXrt2Iiv
8p1vMTkqf9xDNIGzsRUA5AAkOir0yPF8x9NzNUbHGC50Zv2iGAXynRBx+9JVzVAP9i6JQbovWfJj
KYicpaJ4QlIBDWYK+sw4+yJWh5S06vc+oL/z5hS0VYV9bp2KW+Yss/rJNGKZyAbs53P/VBkQ4HAt
yQX3wU1hvsVGxcIzM/LGoRar9iadB1qrWsGvSyLGhXOHbbSUtFUYVvznJv1wat9L4HKMKnqSZidE
6lDg/Jey3F0hKl5Rnev3+R2FjFqo8KQ8lVNJrBe2un0mNIWgkNkQnRHiabTB/8YJxEsSrGpsL4jI
NWmP1u6SJCtAHNZECzvHVuzaGWkL1iDQUVhLQvWfb/pDX+/aCa9OAC7OzHCagNwwOgO7ZCMwaXz4
6cX3LGyRYNTGQCE6KEWEmVIByVIitAHhQcT79r9ZMkCj3CaqaRtK5e/vPWEOU02b0ugzMvvDt3Pg
yTBJaRexUwuLavwmGg1GTQ9KwZzpHz8m4mF+qMpvsBMLwfTBaT3LyiOIjz54zawwGuwOO/5/t2k7
cu98xtjDBvvzCrLqOnoCeG3fSHegy6hm/i8UWZhdcc/ozyR7j6ps3OuY9G5VGN83L3gSMPexCtur
bgOlU4luhrqGvg45See9pbPOfh/fT5J5vIoUxI3MlEk/ITbiz14S5YW9H/F9/YAyK6EyKOf5+9vG
ApgvsY0TvxGlo+mSRy0TrqsWNXWS71EsG6JBFyypyC9WBjj7sl6A67Z1kwKsWXtRWaJcf009cLIX
yTfwpoTCzKHm1XazncQOwYVmyjvwnnhclwHacTXZc3/JngSOT45wb04/THD92Vo2n5uq5Xz58qII
Vln8Dvar4iCfdW0s1fIy2B72EcKueyELaUoG0/WAuAc40izXINGSdts2TQmZVkN92wm0IK13r9vi
OEnduqpptLnWPViG1qYfJwwLYsMvbZc2W/AZlcPJ1DEiuXdwQtcQNO2MBIZ5PKZvCWCHSpynqf9D
jMLPdqMUr3HgBNWv9Lx6V8UBCJIYEckgV00pqXXZ9Nit2y6xP24Iw4JesNd8g33Zd2nljmogeT/u
Y9DzOhdESwf3wPWkh/XVKnV8VHZsFzk79ojXLkE9Zf0NULZj9iMhrxMPjyHh8AXH4fSBKL5eIhpy
ELjEyBJTzStecvXosktkS+lcsyLSI8LFye6SU66y+jYk4LbQ8RuBE8voQaY+9occJlnivrAL9x+9
jdEJdXncVMPBfyXx8hzJw28xwrEIHRB2XCY19koHwbPICF1s42HfAv8JlU7JKnLrhwhU10jpAP5A
3UOraS3r/qItb7gB5MGjNyEAwIywUpiOOAgGeqY5AhH8p8mZN0cEO2H/g7Q90OjuDhcvH44mCMWa
UGM5zrCrwXV2pvxb80scT6Xrqa4JG4QEr1Z8FdqY+4mG0GcWVfHpzM0G45XuWjhCJIKJ1m5ZRKDf
gu5GWmJTFgcRoIRh5yCpRYLhp4WGqCcObxrfK1PCehBNSSlCo94dc1fh3d3Qs0xPg9uwRAmdw4yg
3ZtO4jWrF1YUXUDbm+qWo0wP0RRqWmklrcl/1oLDEqKNQQO8I5+AcQHFGM1eGGy91xn1xOrULUd+
+BAteF6vWF7PeIWkSh3DfU9ANyey9b+c/CbWhudkIGQiEjBdrfYBxXaLRHrllxqzIHu8Y2Hhtebt
fNLMZESVwzMBmu8Rno4ywSbNpe1e9A4dvudTgVbu+5sVEumt5YnATNexF9D4jVxRxskHMLqmij/s
ifJWWlCojNuz/gX4o2ckGEasWSF448/Nvovp/RdaPXVoMgV9NDbtv4KLkwD2bw3hYL50UzKoZe1y
kNyzn7P7wxJt7FMiI5cY+DJeyWAYMcVqD3ofRiVCR8ZF1lUFq1NFS9xWRROlHB0zZGURlBKexrZM
EGhVi49LOhvRRZEA+qPnRFwGsAggnHUj27jnZIZhDZs15Xm5I1R5i49hkxcnndHf9NAWDBekveO6
UWQL7pJDgf4u8r05qgR6PDP/+WoF0c0teR5uBEa76IXtYlsokteaFSDWiFYsCO3hOk8Cd5N2LnH6
s2MntUMt+9uGyEJjwZLJZKZLmV4lQhZrdCRSec6PIvO/hUjrZhp4SxKZaHw8SGGGumjjMHsC8eNq
FW2O2T3o4OjkfLpt+HViEJowWBb1+yheYG+vm+C91PoIEcyqfdCgMwwLhIpxtS22gfNbqgCZp0xG
/wMDeXDGI3DVpOn27Xi01ubPX8A8NhPe7Vkezol+W50YHE7DEr9PQhjGomzhrDKbcWd15IMV9ocZ
eUu3EqaqwNjeelUXAZ6rNFc6+FSgpMmtzQLFQY5Rv2YGtEXPn3qMJM/pFEcH/O3ZqGe/SWsxR/eD
Iqvs8gUn1a63zSdjVE9gR12uNpxGxGRJKueBf4ZR4hUmSSsw46vSYBI55sTmyE9KbrGB9QnOYG96
K+x0fKj2Tv7hP9N3r3UsO4dxdrVsz13mSnmTbFd/X4XBQAs2rxT8vMUnU/arxaOtm3Wki8JZbfnc
UR6KDBmx0F9Td0dEaEq0sFfUZUtM92r7CjlekzFYsviorxcvjbIgtNzE0EPWjHYyT/xJvUzHkxq2
HmwHAjpcv4PkW+byOwvxvxsPEJBh1z8gOeQ04AtHltNiO0UW+GZ5kH/1bFHcGTiUWnDl5HutH4+y
EfdJOTr+NFc/In2TuK8+dlPy8GDjJcOtv3vrqCvtmoYsCYT24XGJStdAeca6PjIPF4w17gsdebbM
Bl1oQ+52rEOz6WWh+7rnlpdYjRGMe8bWb6TPvqy5CB3XDRuMu3QMbIIKMKLuhl1J7P8CfRep8kI7
as5GRZAnZmgOZhdOAsdjyf+P2tnUpEdQS5Hxs9e2HjrMMK86ZRi6+m1BKghthYW9KyVZEHSrOD+X
/y8fVvvnpJcBY9azLv82bJaJxAG//QatLtVFd3m4ywT5tiaf7c/UcExyrwxIPuVFxBLdbpzJXTaz
5OjIOqX1+NSEUYBiuc9C0AlN3rx+Czjyrk/ZdRhokyaBVuY26txh/AjAH71BJrPE8h8ezrN+5ucV
sE9tpcUTNqiyJKV9ZkulT1F2q+qe7RdQVVPKXs6kRFn2m9tieE1guKz5ZAdiftSYPY0dXT9kHwfB
gJAGjpCQMNiBo6Oa0xioIy+uk7pYZofQIG58ST5E1HqkQtw+ENUERgH06SbRKf9lN2tH58o6q2qM
jgyeLbKdiOmiOCM0rbuPjtEu4sw6JBDSEwS4IJ7CQd12WVYfAx4RJW799aMY6LiZeAc0JR2jTHli
DUAYT0yHsnIDGURNrOfvL3F2Nwo/UOq9GHy0kdFWBvDa6UZ9gzfHgldLx/9TnYljtnShps/NKYmY
hIVoLwceNFAsN1VbMwApDqDMYnPcKQ2tcdXAv7yU6QzvFLy1TAK13g7gY2ry9zHPbfxBX1+r8SXH
mdtTi1eAGahzKzv/Ak84BAyqnGin8f2OTZ6tD9EUpKvpCj5CRiceq1F1kkxwcS/zIBhiVM/oi05+
ViUJ7EAySUsD26Kks63i13ia3OFBxbN0sblShDcZvYGF+MGLP/0ndc9qEI2XunjLeQOZupShIpWD
pGRI0jm70a7slzTcWoOgTm9J3qgLOqmsakqppIasuyqvWha6TguKsUqKb+lmXS9vs30iMI5JnREa
r5dHXgCeMNvn0mVrZY73sRgsAScwde/ueqhGj5jKoW9QfRfnfBnhc8GrB7j5wE2OGbaXlbhai1LI
ugQ+t7EeHwMUr0hQk8TXnfqprNtEUMTTkgrtranYWFvbEe99VgVnAbISFMT5z9HXVi0D5Oek3Y4w
VQdyyOeTU/2P2n//+7K5GUdVKp8k4UJuwON/zM7lgDh0ttDmh+lgC/oIEim81Y91Hd1MW98/+QyX
26srk7svvYWKSR/H8HP4VBl82GOPw5vLZXpnaSR9uj9UIdyQdtImeHnhX0YvxsENkYFUPeLitWHX
frGhf7XSCA/BUVK9mWRxZL55VClhDvp8YbcxBdWjNcVdqKGYf9rxcnEFQ3xhnhOi8/uJevF49YuQ
OtDf7fB9Psu5AlaSfVo+WNDeN/3Mpiie2i2f079fmVGL44EIwRLhtwRoBdVGiR7B2hhM2KCkEAVR
r12wmzSAfZN/kFP/+1mV0481dAoczscpnYHNDQBvpaY5JhibMQSKaJRRUPurLfJxRAISCEv3Nlko
yaocvWRL6eSOILQPy31O8gtD1kk0P+aUpcVEvZvweM3YtDJLFNLIfWnNbYKRWRWP6CCENZPXluKO
Utu/Visr/YGsLEzJ251NPDQf8AD0oTOA16mYkjM2rPQ5fH4EovygVCnk7oaIEcMde8WCL7Xma41j
/Shyb4pg5jwIc1TMDfZIWDnR92ZaBAS6lofsw/QGdG27Tzswxo1VgHqkl8dFMewczZVxEbWm372l
d3hXIVeDxggDJv9xZlYxFFxKL6xkzYQzMMP4Z/lzSveZNzoyVNGboDgeEWrxOje+RS5xKdLW5avn
0lA8Yivk/qKIptdtjmEm9qgtWkd1A0ASNYGXVPMIQy7kT6a6M01ivc81XZnfYsbcBa/OkZ/sp/tb
FNURBeWaRVU2oe7KTgQHEd5Rai9U0q3ibCbXpIjm6Nd8YhMeSbnkavCh7+HVVbkSZXhK8ZDSpnnJ
dUMjzwCdrb6UOsKBHgUQyq8Iy+rSA8QWbmjoJ3xenHcGwkJaN3yqhR6DsVRmMY1vqf4rqoT1KyMu
t/IpQr29OMLAOwSafrPMbUKL9klE0AGRJx36CxhRfv9EGdy/dG1b8Gqa4kSvhriSiOcJk0uTZaNM
DFHhkKq9O/3GGgkvZfjF3iMqcJ6ZXFk467k/W4bq9Pb8XeWCEgA3Tavl9ONTNcEZfMPZVKZzm+Tl
A1Qg/JGk0RAQ5r49yuTE4lGX99zDhwd1oMgVvOAasLYJJ1YgZcxZFZbFIyDahGiDKxdK4YE0hoeQ
Dqv+R8Wo2WvVFqDoaB2didH1fcS3VmoOw3Dubtz6gHdDefIG+Lqnrpe4J7wMiU5gAlrXH7HfG6EL
tkXmlAXZRZq9WzU+KZZx/0+AsrFb1PKQacVg2HxR82Kt0oeiapWjsdHrnHlVj0wUQ8uFRvDVqCG9
Uo9NbZNlfKKaPLActJhC4MQIdhUgQJkSPiDo2WC9h5Bp8JkLmxCgqdrAcPjLYvUwZfSZQlkoYrh1
q2fCiPvOWMezFDjjNntQ8ushegl9MXwszgMwBMHuFNni9d08EPMAhGloJ5yYI1d9EuqABvy9x4wx
9L/s1Lh0f2tGzZ0CBk7tXNgHxbUaohu7E6U5813XlACixYu9V9q8qaMmqSFqq+uQ1OcGdjMZrDL+
9yk5g75Q2+dKmCRIT7vpcheSVKIk0E8w372NacXiS8BUjSAETX3sRvHJwFRHh7KAKCO45ZNZTQzR
mdi8ggl+CFaddILzzMOnJIueMf1npHPDSk9PQSXCFqcdUVLto43h+BvyDnGuxBb209BEAxiQFUfK
XyJXpj/tNag6dcEpVxG8XP6L96UrT0Vy535nhEBkB/FvmIEdxKNRqksGnYu7pnz4IvXI8zgmxKgU
Hzc7brueZTh04N6O3/FbJUgEfiFp1ZPDJoXwWD3+A2sKgR7lflBn7Y0hqDAmKe7d0NTOFXLhTK2V
OxRhNGrRzXvfFmi/eTpQDceBY2+BGgJOqjXZm0xzzzaKBVERimvcZj/LuxjZf3mIO3EKZ7cyni73
q+Ht2NnrFFs+tnB/QZU8Mm7dH2KK5aZRZFt/iAnjrz0wD1Pvpx3IDJUOyAhh3J4ZQpjAgcZ3L0dl
+uqaQvGVCQ3RNji1VokddbN/vRWCCpZxgODa7OqPYLEmAxdGRwWJMEuHEkTMYzBDyuzPX0w4yycZ
ZCfo6OxZIt+bvGpJreQ9c5VJmGabiBXrHLHsE5q4Hdi3Utjd0jOFRl1N7g15tWsciq/32mF8Cs3w
huClaRw56ZOZsXbSXwCyZCTNcrtisr4+tBYzF3nfrdHEsfmJxBkBffcWeI07fFmUCOV3O8znwXGn
kRoHKp77j7eJusHuVQYXUFXY/Xgz574E46t3xmyhpSt+wZ394G3eIXgrOu09naR6pi92xD8kqfy0
N6VRYRlxhbplVRr/+HvjHBMLhydsp4ghJJaRc1SdqzZwDTMYfkt/IYZSo6DN+IjDh90efDvJFHt2
HQR46soq9hDZVxfYAKWHAw5TU/oJYG3coKOBi/EfyK9VEca71RyJnhBpOeOG7xOhPK7AIGQUROf/
wP4dvMcfATKPvMmY3oOLoqlnCojJF0bUqPcOtwLvkcmB7+xI1wJiPCoiG6PVqvloSqYAywU6/CUr
pdDnCdxA0Ksm0/fcvNN+Kpi9UltinvRloTyGUgWoOlgGjy6I2mprT2YulTufsjP+m0Qy7PmgamCU
YnMaDgitF+X0h2QZygflMfWWpaRzsw9v85xXscy11xFWOOly/iuYvuu/1aiegg1haLybSPMDchrW
FxUxURYHgo58nqB/+KISkymxdEFkkd+t4HpOtI3tnnKwUNjacd/twAp4JXcVC6UzEUOjuYhtOgxH
UGzjGSFXvOVFhr1K2rdpnVRWJZafoziLIcJYMyCaLfJBQAJhZQRbJT37sQr9o93RqDxijcoZC55d
Z18OMMDfnyKWw98dumNwyFpCN/6lVb0QNTdf2r16CEdp3JV744m/zWLWKN6DMFVwV1+sVSmbIuMq
KKNXNRZV8RBQky09eutBUUf4ravQrghoyt33KK04bGSFfSDnnnZtqeYTsd1QoETxKQovkpIAahUD
mN/geXwHLPBTQJy/y2Y/HllB+fUl25aVngmnaCimhw8D4tLGz8fACbEXlzof0wXv1pCFwNXN0yPb
dgXZNEZIKbQhB+H3UPRRZWyLHyI4fHK3bjRYN2xmrgLG3OqJGNcdjc1kRmrTLsW32x7pkuKjM4kJ
OdqZ/N5jWdKkoqGHmqvvpNH8AbsAt4n4b2cA4Hg3vG19L2ppsyKUoJK7eeDG5I4ulrLOSzCHkEnv
O4Ww/V8ZiQ8Skm6mF3q0Xt0FJdtvXo5zoyLUvO3eByt/K6ISve489OLoagUBxjsnDU/y8Ri5GhLj
hsUMms9frLxZXAVGXcXHWchaumsh+sFz69rgOG72J7awODaz2r5QQRR2A39M0adkuGB1WXDN4XIB
kyyN7lBtuM398e+5Z2hEwXBOTtqTp34HRAhxxO0KecsrJ0Z8xEyItjcC7sR51niH/8V5L1nT1V65
3zCFcRwa8wr31ly9Ns99bKq0mLuQUEKS8GJDUPcfZACjEHEo4zJmdY6ZTH8+k360XoFo+gSWjm94
LJStpqvV11F7eoY8ZK2jU6xYQ/0OL28osWccrF01RmopzYyO36gep9HyxgvORcjquhouphgGcRcP
//PWkJk3YkCCwkblYwPj7/mBeeY7+6sSJu/XW1f/LQxpoAJ8P6aUVmG+uGGRi3Z0XxdksH9bDMRy
b7+GLFCJkOwBExky2lh7g35bTcYxjmdGZvJsnJPdzxU0j5RGFiHCLwdZQcXGwoOTk/In6sgu1GA2
m4ByBsNjSyjnzCX/WX1JLeXQXmU8bUIPKcptLqP2OvlRq2IAw00AeE5bU+FzfbSzeKOs9hFn50w/
XsWksilmePpQHL5cLP2ZSaSeIZVS1CJ5r1I7nbvlz5cf2amRFdqvf57RYcixWV7gqN3MNTimi5lP
q2mpHaMK0DbE2VORPXCnoEX7f99q7Iub1znhuJKBGVlO8PqXgUqOFUXX5pK+0SADoD3R8yvzXtBv
+4+tXYDlUl9orhACxpxFPZuF3Qd7EhVqoE8NQ0lCk7LGgy1r44AiA5G2oncwWg1eQrwD6y8h8Jpj
suRdUrL/C8pEX9+kUrB9ar3nlh5bBfJmCygqqnVh2Vt8mmPIGQFwKMFUl0L2itZpCbXmP5Im2Rpv
fCVPrY+rkRztoXTNaDuXydLkEWuXxG/oL/avFpNTeesmX8+swAoNG+XvHH0gR0w1iqH/MFMJNRow
AyvSOqoL7ryKqqqYOZdI5JV0hZfyJGzRFmsFC5aNg889qwOGjEEvfqtKdKWAMjU2eciP8j44iZMN
SAxub0UTe8xYH3i7kX5M1piMa7yh1E++FiqFK5+k01HkTQkwy2vXw7NINl7XRVE36y93oZ0JkrYb
d+yEoefE8DxRu0aVzj3v/HY3UJqeoBxliu0McdNvseE9TKhZq90wE+Se6QILsBR6wZHeYVrP2RDU
4Jd5cl1Sqetgwg+xyom3+tbqas0BebRS2rirydPYP363yOgtkcTylOdW+S6n5Fhjk3zb7tTfP6mg
74zrKqhNABGsFmBSOS6F8JiFtrQLaSmHkVkv7cUSmMhi2nXNsyjW3l96fmfED26NtiYBsDzEIbJe
eTKn9IhdVoNt3zJjVP0B9g9xmvSj3vf9C27cIVMbk7G8xV//SpAf+R3OpMM+aU0N0FpIS5XXsu2q
pNmKIulh61Nt1MzJPyZ6ZJeWfKBsz894mpPUq+hnxPNoviZydITkP/KOKItT7Wfxxp2afEy+IzU2
5UWy4U2qi0uhHESnEJ5ZTWXiOZw5VE6bkooMTAD4puKTdkw7/04cji+UF1Y6iPxp3VwQkOfbOGoJ
u9do5zmaHo1uGY8/xhUMiY1gIVcOrSNjSje5V1ByAmyHJW9To1yuQK/hwS8E/bvlORkUND3jolpR
QQPIlC6USHX13f/+O3py3ZRR6Ec/IqA4XhzV1Zk2YFlWnK6DieDdExDNdGbtGpd0jxfYwCfNvlBD
6tVhyMCXeId7BjFLRI1V9gJ/uytM9vGoqiEIXQheeQtZZH+dE4qGXnYw68Z6vWONd8b0cVQwfEE3
dKp56JsadoZxc6qU3M30Y0tB9eBgfIS/vVw4Dwnow9axJYiDFMK6UnSEVFRNpOc/g4RWuNLlEr9E
18CPnkhGadgksGxG+Oe6OGshiDKnQb4WI1rZENLn8kC1DtJiepfzjUNDH5YGv7hMCJ3SI5zTuBjd
kXyqkamscu/A4lfwVMhx50/hcdGNNOWaJ04bMeNx2GdYq5HtGlYBO04eiwMrTtkx2fY11ZQ2eAst
dANF4ZjGdG0wfVZjpkxrUcgiAwnKNtpQirZGZdXKbWdprGUozgnfSyGZ/PPJxMsIVFVcMe9DzY/U
eSIO0vGsi08zv7ANuYDIF+aFenmv6Fu7ahpH6hJTfRvoVfLPrR3dlno12HbcqpmMFOGV81/nTKrL
OBpCBBaor+s20csBjW10jiUuuMNnEOFRz67gmNeoiLswdMVx9NNBaOuHK73jx896ZbZEr2BdHnA2
cn57/G7sMn1R2ElgQ7LuRdaOspuLJuq81Yyu4ZHgcx0tYmMOS4L5J8zT7qbkZSk7taF5EL3BAZuY
h4toJ7RsYgZGLHytvjQmJ/W62Yd0UMC14ZdoBUfECk/P5OVkepVMeZs5yVfuw0QKLIv4N0Qoj+fI
ICayxokwOV2r+yES3u2jI/xmYazGyQ7QKDj8thH1sBQcKkP5Iv6dWxYAleqoM1ZgkJ61eJMeRIFU
OC2vPfyL62H6QoiGOUPKFhgosK2PWOmPB5dbazUGlEvJnbrjWCv91CanJZGGei4E0vAQLu3fkzrW
7s70bSttki8sbvQDUvJkc5ZAfG2ERwoCeeuJZqR3oPI/LorCgMXi6R/33MG6fV8dgFapv8o8gEwZ
w4NEhj6aNG6+XX1fmsCfPOBGyXsEo0Ej/tqNjMgijDEYw1Mrpk2HKJ8u/fMupYrUZE9kzaIVF0+/
vky6j2TAubNMhumBNv1M6TWjyZZiDL5aZY/8GW6flO39tcGcrREFwE2DRvjdZ4gchsakqdIW7DiT
FiMyrQnaYZ1jtSxk5Qdw6xcUG3E1rdjLQPHC1GbJsIXljW25BxLvL1RRpsF2jqiaF4iu5ejwz9Ih
4hsIb+1pKYNQtG6Lnv2G6Bc8P253yapgmbb1Vizp6IBjxzGsrbA44aFE7OKzQ3Q1nEjUwZrVfLuW
e8/4HI80QYkpYTVV2bhVheU4A/Fbye+ue7tvuOrZ4W2ny84vt9mwVs2sBKIFD+3XEkUL7PSjm471
59/KhVp+Fr30N6nVtp+yqac5CCFUGzOFlAYPC3WDdzatqr+FmGX/Ha4NKwqmGM4qdQ73NIDDcTqu
JejVXrNX/3VxHsmEPWjHoZJIOUHX7s2sfeLCQ1SpZZeBbDz3Aqg+BGCkjn3Zv5lzjrn1PE/C6yAB
4Z+0Sf+AFN0d0xlCnq1q+ndhCDa4L+XTTNQYOlg/R38VeYmMADaE4LF/XZRRYHOVI99mNhDftioi
VQQ/lJysDI1cEW8OCVxzAFWCb3eQfrTPICq7yIvoqQExi4INmih4UIg3uh0shTp81Nnjl1bEONIE
25viYGHg0lLXmDguXwGxreZoF78TCO+GA3to93MWoC1oHTHFj0V0Y1Ty9J8ZdUH735Wsf5lcUN0s
SsJYzMnk6g/tI7QINlA0RCUwI7PRVFZJk9PGejVqNhHiZxVcMt6Quwukz8AMgeuSnrufExir/E+X
bc4BGWE37gELht1VyQmcRaTd7kCv+ZW6GMarDXs0d3y3Rsj2Y93AwX1VgId2NPahhoQHk8xzRZZI
sVNVNhkaJkRgOfX92A8cwL9K8Iw8a/MY7OEzaIqFgCwmYpO+WInfz62MWFK0I1WoRkpfmik4ocrD
djS4Dd/itPG86UzVcLOVd3lOZud6Y5MSRFk+cJIOptPhiNpiwThr8o1gNsgE6PNvrI0LUAhJ2vH+
ZE9FC15cz4ZpvKuBGcoS6G61vcvEfuETHLGeWJjv/wb+DwNZo9VGInzboA+Dj43PsOfQdEnzyROt
HGY5OPvmRA6Y3HcQHK3hw/Scx2JBB6P/rDIn5SVsP0/O8iARsifQIvEj+LW3Che2LId7M4xjP+mq
CmtxLBbq+g155c7H/4MzlF2cxD5mpTqrKpm6b1IVyL6P5s7SQ7MdJ+9qnhvb/z3CPqir03UxV0aI
yzfKI/H+p65ocQKmx8cP4ObJdow3IFLoHzExcL+aMb+lOG92JVVdU0+zGbK2ywUn0OEXm1xAAI06
8GL0pFvzwroCrI2KhE33lLhq4o2w7xJpgeWycdLfuIzGZTu3Q0hewoTH8mHLly7QoRMXPXd28Rtw
VncnX1mQIASQrRQhdDktcjFxLf/+eUxowZx37GSrEq5wuLq6z/lh/apHcWruChPxwCXHQrmU8OGe
MnFbCSi0avc3WrGnznEJDBv4TxHp3WeqNVSneYpkJdwj1b09COzlNWulZ0/Qhtg+yAZhV2JS7Bma
NESNBtrK64lcXqhF6IoAxxAZ3fR9qcY+VbJL6eVtic99Y9gZAQ2m7f6V7xsjPaUw8DZVFB1X2Sno
Fqzeu0kLbhILSyyn94VNgE9/v3VMNg/74r73ZgUsw8ddZQHYqveJVNVDwCgsDfQAf9sN2YNkWyFn
cStNpLaQ5pTCoX4gtmFjhegJ9Uh3BJU35RhBNHaB5eiSlMY9em7JDnK1DRSGJUEnL/SQAP90lEtZ
lR/bEv5y6ivFymTw6CXsGV5AOzWbq/VU8TvzCkAW3zr/g93N63yGrhJrbEVwrfNG6eQrQJevOLBL
7VxZSv16SGgWzqNL5QRryJJ2xxze+nwnSyZKPTB8++yjAaBnBP/MNhgXyb85r3fwHcRBdT/psHbZ
SVEmPzra4wdCKUWU0+OVJHHmHaSkxXCLttsMHyTmnGPTuzxDZYAZ0CpATIob0xFcT2RuNR03Apru
TSsBN9TY4bxzt+LtkCE9/weo/UBk77nnKdfFbd4HGu0z0BXkoRJZrsWq3Z3m75YRKyjJHMG6T+i+
CMfMwsa2lDDFUulnZfOEqIyXvOdTN0UxvzUr3VSqszd14Alb3g3+lHOLmNl0Dx/DqLGVvOtIhMD1
ZcG5HE6fsvDyzw8ES/Qh4kWguIBlvxpSJs3R3ijPDahy78cy9nY4YqTVZljBsSBWcGApw92JTyF1
IA05Sae+EgeQ+LzJUvl9sgJeNMZSuO353Uq7Efg4LFhJ3IAPAj8RlvMAHVskPsogVXx6yC31zzG1
1E8qBb8ej3wjTTFKtW8nQEt3uIR7oYW+shhkKmOXuZVrcAHindYyN8fgfC74TWuh8WvtLrnUXqN3
0D7Bny/s1M8QeeWsLghDaM+mobt5yRpVNi7P4FMmYfqMc5cPP6LZOKO5209vFpU1gceoZMwy6PE1
5bqvgU0Qj6iLgFzUrzx7Q0vBXXI+2x+GvcWL8V6H6W/H4AFXHX3x/KdN37g44XStEEDOJI1hqSDb
ykW7ciQOoWntk+nX2BU7lfYIUJzB/rh3wAzeqYsIADKKMa0WMqGEdbs2mze53RHfLzXU67la8e86
bWF5knrqvE0oPHD5c1BXTJfpZP7VLdoaOhIpSfAEkY77jjsbnJ9OGyNgYsF1tkvAxEpYwOSgTd5m
7rU0eUAZdnb9EvSw8G+2T+A9IvWTSPvptKXOiIE09ltdkObrUtxFGDqh9sb2IeVKRyMp7xsX8+uD
MlMpdQ+aP9Y4Kn3TYFTHNByrCdAPj+h3KaqNJ7xMi25TwXQ0evLDLBWrMGhSK7ShJaJZ6L2qEIJ4
t+UWYdytYIBVlV9K9h3j5CbvmWC4fnKeWauo5bUgWkg/k5/U+XiqRMT3rtDgAj9p8jUZWcMl3TiL
tUE6AW+D+5T4cOTrdLQJCzSZqTuRIJROcC1Ot0snTvU6jKWWx7QUzuYnVD+Rfjps+doKC/PRP1Wr
q6WvVveUGFqYLWEhYKmpoiVaDiv6jby61ueY3E56vYRnobf77j8GjMiYVW0DmD1Vk+QMHktKVPUO
jep4DY+HHEBYkolWqag8WkUjKIcUegujMVUf/Lz1x0LHAAiiUVorE89MuFOip+i8Z7EqtQHjArVz
tTVTuCBEpGzFWDyQWl8fmUnUZG1HqrCrBQiS2jC/Fyv66Re7VlpRB0Ah3Sudvsl6Gpi12EjwCAew
PQ2jfMlJN4nLhy9lvNXGqm3BCVd7J7Xgw3AQVCynMpbhSJxTMx7VLLSbRw/ikAMscCK+I7xQQtYp
nSckdW+FLhenlEpzA3Fo+9yAe38kmMbwcJeDrX8zcCtVCras93rDTTdzWezWgsRJpQ42kxT/giWQ
gaLy9N/qnOrxyvaCsGUWTu+hvLEtsAUk83lMzBDJLHiKXteNfJ2LhYecDR56g1hA5K4tkzIIKava
Thzd/f9ZY50n22mRzfu1jV3g3rr7nziAllDNtW+UvafNstUCh/D06PYacPj6gjxCprCZQGQi8gnY
k+Bkpt0uHbCgBs0Hx/qyS4tJoPGG6KTsLFQBgsdwHHq0oclX05xtG6YDYveooyaAOVUpjBu7mdpF
QGldK3SlEXMfitcJN2vPw9PExaZ3OzuGj3Z6avm5bGS1ZDgShcG/aZTAj9nnGkBd0h9GPauQG9NJ
vqZ4ST1qlMpPCIiJarz94awnwNmyvgIwDJaNcfXofy7UXstOYHSk694V8DdMzrXK6y3xTvlfqbb3
o0Sp2WiELgryIH80t8WoEK+iD8W9PfKXBtUxCJzHkXYxiZcTDmAqaR26IHwa1nvxobeBrgPGvzQf
gJRJyLHEXOuR75T49HPyShZRL1nvQDFT0qkCCDdiebd9n4KvkCeaWmUqV/mV7Y2Glda5uXG8W7r6
/ljDN/hhhLo5CZze/n7JL63fSbq+v+dtu7PVdyQn1+q84v9Ld/uhKFPgqV+hqlMWRy/FMf8wdBtZ
i6LRQrYxPdpnBTMgAmW4mApuK2tux9vpkcOlsKj2qFxBbquYeEg61p6raD2CjsE1oMOoteOPolR6
CjeCDYljqoHcEOyJ2t0ZHKfDV6V8pAI/Oz/HxY48Y4+o8y5Y3TJrILCzNIm+s5EnYQMTLEjQ4x8v
Yp1bYQcRBS0Xey0ICU6dH5Kx//xDidKZpyWfZwu6yRenrWVZ1K0ops/f0/vRl0w06LpUceCQPC3C
+HibBMW+1k51FEo6PCQHAoVB9IVAP1IfTNRXfMAuIRga3mXPrMbbpJV/Vu8xQGGoCJ+wdZocFP4X
9dCxXgzR8ChTwto73SmLLFidpg2mWt79K+j3WVO80sltkP6EO9YY/1vxRMZvdyaRmAxeuGJEl0+w
ZNUdT0KO7lfAV824OtRtV+XVCV/wT+Ce6vjPENXeXJ76b9CpRPejVxJn24yleSHyiO9Y1PpJBJ+l
eJEiW7Jo/VzaoohbtTRXkttcxshLkBeOEhGMSv14G5Lqg/54cdy2aBO3khHNgPIFKqu2CLk4qsS1
ZQIPiHHr09dC/qgHOAfUU03LDzNSALmBrWjfyyyqc2jMk+TE+N/wibPMu/QtWcJ9fsHLpFpcxOJ8
L7sMun6frgyhy9MzNQbi25xkqZ+WSm5LTI5u+eVa+v5Z1D4Yo0jIxfb9vDNJC+BfdUMKzijmKoFg
GEVwdMn+Y/XY4z20Zb5qleif/E1BxFYqpPBqBm6wCIqHr3UjKsk8kLRgQASReM+1j2WIFCr+Iykn
3kC3k/NtOn/8NxgP7/9T0BODwaFQYWfhjqAAb/caTV7Ohm9mHKehFhSrBRDr6YXEaHi8Z7B6Vsey
Kfk/l4iTTPbOOgtzHMoUY/xM46yhFatK17No2EFbNtZ641i8AM2yO8hYBGMpYHRwFKxJifi0PSND
KCnBCuTU75Cfz168lYNrBdqaOmmiKD9pl5GHUfvs2YRuYJs1yrhN78iQSq25N59hzPfoEO4N5NLD
5jLJVEAPTMLSs5XOqt6QCOoT155PYwuB/EUJIbZnnS/G1isSe9unzevAaCpNMu2EXCWCmFiWCrXv
0MtYzuEOvifIZB8Ex8PvACCRpsLR0rQLAmxgo4tw862qqYQJIAGyWM9zWrkKvkaCal2vezmYp23O
w0zCeFpJQGEcEqeo9KS3EOPqQdspwrCfUjiP1MyKzHqoCRRKThmzTF+e/RkdYtBj1C0o3fEk93+c
7GsAJWTGYaiRd7V7KiidYW12F79ha81DBvHHcHQTuKgVNo/tSYDtFsA4XCTwubEUG73NyvY/ovjg
OpLgwSuv9mhwnJ+xibNY6hSFajTcbNPp46u2kuC9piVv2JzxrEyy3LPVKtomYEF9hiMvYxKlJR+6
iCB3vs4YYdZA2DfGdBT+4d2uvjsuRobHfT94OaAa1BUINFS7/buW2fg7gfJ8gJT7ASMIflgZ90zS
oPG60zByKGv5iXbeX90KDmIIBTRQ9nlioBBzyykz0CiuOf/Oy+GuGapGJ+LmQMdjPl1mUBg8MEv1
SUqX2gkYwE4jA2nZmgVC8znSNcYKCE1xGDXzJQxCyQuojMSUvxFA7NKNamvlLCT5X4hZACn1HyiI
3YR0Fy9l0Ab9n6TpiJa+XVsnJwj2BqdakPfmzNr90Zrukk71nbIjYLrmpdfgKRZ9UbVn0Mp6toBJ
TphooEXXyve3AUWXyFRxCEc87wMarkyieeWFbRAHydFpe3ODOGaLNUh15JtpvNiNERSc6Ta6FSIW
Bq2Bx5VP7LBA+muyLqbr4VYb+cSBjNv0txO2lOjjsvskc+tPGN7TdvdPEbBm4Px1tvynM2Z1lxg+
9NYVSEIjW8i8fG9nABVv0vn5SNVZquXJRoP5ba9IHxZMof0BfC/gcQG4ympgU/cNiYDgoa6DKoPf
b1/b1RDMfL+ei6kYTO5ZjBZBu5/WsTnznYZXjq3UGuAz82l0d7YQsUzJ9bn8t8gFD3CgoOyZplPb
Lz7VTE4qqJvkD/MyMkJt6jjItm58GZteMGkYRzyWQtSkUCRSD/LJgAkrvg1io8ZQYJ1NqMVW0wrk
wRZ4QrLezbRe0+3yEzrm4TTnOI8LxSgAjw75c2PDaFG+Y7NEV2c9z82hIkrCoBHPrTl7FYCsNR5I
xnModFCpuO+txcPfSR2r3fIDHJ6ppbilfL7h+HZFqs+NJQyaNwGIh3RBeencRmH667OeTg69lNU1
xLofilQkoOKjcYa+dV5LfruxTrF7y29H5AvTJqe0yZhNgqS031Ubovg0e0/9L7OVe9nbygiA1nXo
NJODB/NnUs4kQnxIrfLzVahJknUL8oaU6809LtKJdFdYqE55xNlspXIjLKTtfkvWBcaJyyFVFQ7U
tNAL+wyTvl3pRqHdNDlwy9Kn1en4gMC8FN4VVzbIlSe/XSdMUFvpvRc/X7DmKrWNWYODY5VdB8pw
K5DAikg+yIuj5Qqm41UyOObIBqB2YN1BZqj+n3/fnxpwRJWXhf4A5VRuiWud+ijfE7lBuFd03LUM
tDGtK8fbVTDAhORpNnaq47aH70XFZiWAHeXJ9Edrrwv3H8GSEy82zL2rs19tbXgSCew21YVJDImp
RBxEDZhRrH8eHRJbcoFveTFYmhALOeOiDjcTObT6dn5aVAXE6TpikorWbLoh8ARLxgtDY+XnCdwG
e6UfuAtma49ycY1CoHsn4N3i/0B0ZApbCZuet8/gvGpZbwNKJ1IG7iHAftj+imUKipMjsFBKr5KO
P0RdA/yLnA3TNIJW6aDiMnFhxfL9yrZ9+ztkjzcfQFodmn2fDsjN01GblxuuG2V/rhK8fReXclr/
Cii5hGnSebDXH3c+d+ZjIg+JzDEBscM8WW9ggpXx2z9nVQhZCefzECJI5IbVUobKZgRf7VuFR6Xr
dlwTcPcNCVXyKeBQPHxiNTot5hUj5gl2RkBVVWNEiO2ThCpolZ8LtDQoBIJlvM/z4P5o2X6gsrKB
8txHfGTGZQfOPZN5dRRVXr80ozoT+/VN80M541zwQTOacinDc0E4oWdBfpZt8NimKXctKC8/vUK/
4Kvb0EjRLWybvkJQIN6590NZsEFlpyeQzkXzEI/GRqy2UcFG2f4tG+xx/UZcnkivHeCBUwZcdX6v
ZeCEFrLVpU0S5uAbgoB4hU1gGtQkcGf43F8blPHABPrZjEYh2858HeLN8vFwnYvbx2e9cYp7Y4jo
SPqmQ1CKpBYBeZjqCWK4oAy50uacg3PtNug7XyvIsTmYHeQPoVHPNCq2uL5Fff2uPDAg1Ibn5y/9
DZH1ahaw576pVAexT55HK0FJGZyjWdWfR9FqL0gz49kKpeMhcX2dqjUmLs9h0VqM2mMyuKRqyUyH
5HBb8XCbLmdAnHdqpODgaEWWDmCwnUD9NHjlXmIUS6YvAhPLGbmryiod2Nxsz07tdFlcIgQ5iOQY
kgAA0D8B486R2vBlVtR/u5SDp0BP2zfba3Y7uvkeYxor3cY+/xIsWULlswZbxZSelV/k6f4/FXdP
I398Lgbsnpfhz3JX3IfTmiTh1B2EJDSNJrnv0cihxNeaRsnKIhJCazJ08DJPYUFk8l5uzdSSs0Jd
pA3/mqcD2vDQHgvLlLszzpYveIdMe7qPxKqMw4K+HbJEeXsw4Vx+W1/h/U6xG2kiqgRWpHg8ZAv0
dLAlvKXe+tfNTuQla9BIVOzGgdfkMF6vrYI/h7jdYNFkcNOJYizbHiQ/NoMsKbKnqGx6B0qt8vLU
bACPG5EbHfqdCTPZQJEeE8GbfVr4M8LHLnPOyaIaUGLgA5I8ibeCErnBx2i0ZvOMMUBY+70xjavT
N+8z/Fgrp6aqlKNY2R4+lGy9Fswh3M2RcjYjZU6q38wFkA5Z19cVJ+COSxKWDe9yDV4a91qB43Yv
WsJ/UN4GehD6v4uyrUPaYTHDRR8NkKK6RCJDH/TwG9p5x2esAiE/pYPZA0pMZkt45Y9v1wRYxDju
P22EwfKGEz2rsfXnGtJN732WsMdneINblbE/xQHccHLu8F95lRnrtxq4y5L3QkUn/uxon/SIjkm0
xLeKoA11rfS5pAarIcPl/PKSq7YzHTsebImfQn4VQuH1daQEcNdAESoVNqBuvJMyocPnd2ZCb+iU
IrVoz1gI9/w6Kbo4xvVBPq56UGcqWaS/af8c6s4GoxYyjsWEwsQSBoI1tTco9cOoaziohHXs0WQ0
ivdGITJCuGXnLsHOLO0BHtAv8AbZtxQ3nUmH2BQld94bou2tn6sXSd4r5FYvTkeySBfXKo6w3StE
ZvU/3+1qKskigsCpu925sm1PuVfxkIqK/UHCs1MwBX9WeSlVV1NmU1IsPqbQjdkarofezCMNBRP2
BvEdrywlrAJG66qS5dR0khWCKvEcB/bxJIUTDcvVs+PoJVJT5xyulu9II3/kZLoOmiI/x8gwWisP
QtxrIOg7erEWMBFKvenjE7IiwlbM//cJGSxBl+ii060SVLtg2rbK58EIvUV3CmW2cBlnpjYeAy0R
z68tH3p1RarFWxicSyYQYx1L+OPnBgMyOfm9d8NLUEdL5z4anbELQMzDn2sC1IdNRI0G0tezisSE
cMgtTOp2sADJbwtPG6d22xgqt49lWOGokE9NNz3mEs1A6/o3FtdXrR1jig0m7UgxzysiNI+KId8b
BhQWa3s4Z0PeoOWHMAVLhOiV7uoSEE/66QJeMNzDPZmYmLOsBgsppJIDN0a58FbmiV4krKvQ8U4+
wOpeQBOVbIEf1sNe2tJhxWC7Kl7gSDq9D8JbVnIs13bzHl/NexQ5bWyntEAul2Y65p83ZC/JicAB
pAmfYiiGSjEJmkFGD1ocmcD8PrhzfTamVobTfa/M3P5p8ovBizHSY+AcA4XQI+px2hy6n3eKl0Vr
a/7vO1oBVhTVciUgRzgWeKwZP2147H/ABk7t4yTO+3XIEbWWweFitXzmDHCDCWK24fkw5iuK1pjP
vOJrYIPkpeoaNw1pVKGSd4wdudUBTeLjvDizMq0D937BS709wZq0iSNxb9RM5AvqNkdWKEMdi5Hm
wBo8JRFGDdDOGIB6MRrIDE3BT9x2WQzlIIs7VObeAoUo29rrt0SjroRa00VEaOThXm7lqSE7ElMV
3LxgPfinoy65TfKcsVGetl79fnXx+u1kKFarX+nyfz2vI+0YclSAbR66+Fa6DsdbInkBZhLP9Wya
u/KYxvPySlpfCfW8++dCiuPOgFjxffP/3z+vpoHlzrCuXvayo94Bh8pWNHKX9cLgJuJ5RAU0ulzc
mZZeYfxgNkRelSjR8Q4diP1wT6Q1fLtEDK9N70RjmM6fpAoKXJrSrF3MXRoj6TIXDv2DuXwkcFzI
s5hJ+4CyqKpgfiadRciVf0/JRAOz5wD2KieL/pDJFQ2drMM6yMR70N3vrIZoQyEXG2lDeVwx8SGv
iiK+NwB+4awJSTKWxtvzNP/GUaG1ZBwDv0BYeQjgnX+DbpSJS7ifAZyccA2YvYDDvJDP5GT47TId
oKvvv7C/41t+mj9ZVtGlAU89yDd+kMQ7IyAPVl5Xk6u6mStHCngESvYe5uiuZ76nyovLEklQeHNX
ET1iWA9qbA/5L8VT+h+XYFGCBTmNwERgHtjxrOJsnS+75kdOcgApPzKuTsFHJd9d0uRINe3QYZDm
H0a2Y+OyeFWidY5VgP8GNtoViavcvNoiLV7LuftwoPVlPKLkOIEAVE3IK8w6ieAa/+cmaK594oCT
AuFZjdF/KkfTpxviE56mAcXjk7/bLzs3QghtxFoobifrJJOKawHe13bJQ5s4MLhWNh13gXpBWo2N
MQw/8s2/UsVU4sjYZlQryUzMF8JnwJqxivtKLzewQp0XXSAmrHUVMvb68C+MTzT58b4NhR9x0mQ5
XJndPGlc9gPwPLDGyk2IjFo+pAiGRvpj4HdUOh6LBPybr8u+XVp9cvrJXrjUyDwP62qBicFIJp7N
RxNE58iQdorR8ykKYcBok2yiGsOe3czs3uhlKkXU+l+CehbxwVBQQTh/W+HT44nbKm0KbnRO0wHF
2YLzKZTXFQwA5H+PiCrbz6ROt9i6rELCb1zdvM2aTS6B4jPdgH+3gBBo+7altj9VJF6rryrImYv9
GOLN400+PHejuVnezOP+E5sOi7MTqQp7jFDyGdhRFxbq0oPtA/imCa7QvA539xcWEe6nSa6h5ZZM
dormnZd7tmApucBVyMU8N9wD5XNMujGuRjRO8YzJmuDSAmk0aIxAMFeG5ab3tA/pUTmS2di4OB5b
AbKLqJbhddKyWwnY5eDx1wLPTDSdoSgTZrRhy2nc8ngiHk1R7XnbaYmFRj7/OPK59jpYLV9kYue5
9W1uMDvXpePxyBSQka7juwKyy2lL1HE+0rK2Qk6qKrHZvv2gFM9k1FjUR8eiqBJxI0Y1iKK5UcX6
rocWQjqCldUI7d7d8U9wZXAqaJfOANlgpMDqrNqIVRPbMKSJYI+6kQX5pr85WZLPx0jNPqz/o5YS
sFuevNc9ENguRTaYwpxEbNGD7JZyviREEHY3QSY4YaZZnr0BbrEz3LD8AEKnlZTsZlXMjdYbUq1m
pEMZY7rgDqv7/CZvpoMlyhmZ37LNqKvUr21bNihn5w2kOH9FW/7qQzAI4VJZvSr4Bl8UUobm9wjL
jiCkF/P5oEKpLuKSJ11PuOSUnR1QnPPHifztOeisUnopgXTtKnykPNFSs9oAx9if9827CpbCVT1y
l1Imch2wrUVZ6FlTb/oOK76qkdFmiEXAeft4KPujO5wpNx0FyvDXtBCzKraqOUAhpgp+Po43KN3g
/VqRHo3O9ETCkVdb9sTdvRkmm02Smtp5knlKq/wOOa8NQzUe31nM7P/hQCx6D0vVStY/UMn13zMN
loXWztk2/qP6OQvB2+bCq2mWUoygZ/c+ClQIzDd/9Lmetx5/BvPVMlxPxw/K3Y1pp8VT1qWoOQpT
nXNyfIUALurPub+h3ebYKVXARyqC49AZk/dfEKoSncb/ndSSOjbuqjlERvV+L3M2w/uhufYXE2K8
8sS9ykUq/YucyZ+QwOmFjUUr++IDHGoEio4/as9VDS7pvV4hscqzTb0rAeFr8j3dTW5uG062XgWQ
6r6mplF7naRx++Ir/kkiAyIzpQwrVkE+syrs5I+nyRVAs+YhaLE8jd0C6uuhZzVHDcuxrv1iHxSp
kIxMy2sydBNV+D0jbXN8x7TaerFnTTuWjfFkVfyJfMG1UsEajpTkSTVNvBXX9PcITwaIiXwYRzP7
Q7Ii1K2JgWQFYlKsVkPReboo6fmohnDmYw3vlm6JOtgoJZcaytDMtskVegKQWB6b9etESjGr5IiB
nMYXQRIlLlDRdajTwV92IPwOQwWv5WAnMQdPPKfC5e4QhJiYK5M+bBIc1N9Kk/88XSRt/vlaIFS+
mCUw/i4Ql7QK8i5NVjk4sNA8dznDj3XmGMG7k8mucNgKsjR37ZMktsjY1McYjgtAuwO+FCPy5CSz
16d5Vbud5sVXvZ1B0bGy9fVFgNcnsvw9+G4i/L6JoDfb80qABtHuhD3CgP3cCm/9M0jvR6cpKDRL
ZEjWChsvf89Nafmf6qwLLsDlUuVb5P9UE/i4cKcbtxyYSOP2RzIeQaP6gu3kDCDvGDzcUF69loIa
xOsDf1VB5Ahk9qcDaNP0d5EEXdXCoCnMo2flu5AIDCDhN8lXQBawE1S4M0mYc+Usi2jBfCSc2wMA
bdbMlECoHQoXDO5j8YJO3aVgKhZKkQhA7o8RW34fsFA5falL8pJsX7gLV90VVLxaDDuUpxuOa2vF
Xkxr8hWVksVWfsPFACXgcpiyWCa6r5QZzSwzYswJzcdUinjOIfNlQQAuwMe9BZRofqFjt6aSKGdP
gyqLM7NQpMCJ12+wScrOl7uJLZxNh+sJAPR3cmV0Z1eYYGPLK+TQNwfCgCIGlX1ONKMQgvUtAGc4
SP89XRWohyV8dfLW71mHjQFEY2ReBMU3JtrMqf/JFquPPq5V+IFiJGHEVQoTMPahQ4tsp090E0SK
a1sYU18/oNxDHB74nE4XYj8hBq2E/NfCA3cB2wwKQtctRJ1xmo7YV5UOjbNHjtNGG/ztMMhWMyoV
2AAd2v3rCE93sW0Ycv408580e2T1CfMRuENIpW05LkDsx71H0iv+UuZZa+84OkjAy7qsW0XWB5Q8
argQFVJF6xJk6/1QYiyoCs6qGZqTkQNXY+SjP812fwboJw9+LuJagGwJ8ydvaWy9QKVzj7FXeO0N
Z/xv2xrm5Qe1GhxWWHr7CkGjgMlXgJH9uRRPox+mPDpx3D+2XRKodAgXo16fcS1RAiyt+BYtYABy
g2YvSMS+xrlrMYu4XYmKckfOPFO59/T59z+hhqhb15uJCXK2RGzMagGu4g9oaWxQa/irvUTWf8Us
s49nYc53Hgoe3byVOtQ3asaYxbheOLX3BQIt2rAhOshS318KxnXU86M6u4/Z4DK/NWAwfpxeZewH
OFwmFSmWUvGR9mLPb5rjL+k3uLw1dVIOI8EBfGjkzm0imtESstNy27rckN82KHfoRmVQ2mA4Jpv3
OEsiIEDi4uVtvxTs/5guPQEvP2QIxoo0SAs1GWeYyre2i5+GQ8at0TRGHphbB+EZECW9URQCFMcZ
jQKlQ1EPn4X7vAFPirhLdp1cgzNgtEbTGqxhaPku7E0F3oT9DHdBmMgi+iEXlAAim8yBY++dmkwk
yYcv+h5VGBhtdw0gS+Vtq8JWLFfH2F7SzCI/kjGw+pNgM+NuEBS7IOPEIGvZPwkG4buG3IR8Qia3
5WR3ChIQLBYEXlAbK0RbqI4iO+r1+rudqb4MMFSc4fkpnC5VXck9/QoR9VjlE/azOWRx+RqmxYZE
WntZRqICI1ge2eyFVO4vr9h9GEGDXKMfu9iL3j+0h5N5fRRZ/1SytMbzSkBhyUk2YGu4ynYKHfl7
5Pd6idhHNl7VjDdd7aRZGJ7T6qMsb7zNQkTqHtpi693HY3KUpjFlBYmPvl6kjmtxnTdJBy+kFkPt
9klPPucgPl4lCV2/nG6hr9Hm5wxsOXoAS6ModeV99O9vgCgijTjWzBdsr0ac7sy1ez2tVnDi2Q7D
SKEIOaNZwlyK08j9UGwWDt/mxSzJPtC1qj2CPPxnFA5SKsVV8/lN47Mi2Hlw+PkKvEpetTCEDBg2
EL2SsihNX/PT0m6l7Rp10A++xHEdpzMY7szm3cPt4Q5kqnkxSg/sNdibKChlL7UP+gyjYYtmFZtz
QkZftu45CQVwYMG6Up3eLL7Bma+yoPN0RBkomU9lIwQ+YtmSHR+kC0Rk5CUyqaOIhiRg7bn8vYdh
JGkLXpmxLkNP2xa2JXLp9yfJQrQKvUCj1iMoeuv7HZsP/TZWnHHc9iJSyxE+9/NVpVRdMn+HN56k
OucUUn+Zo6ReUqotOXYOkSsfkjaFO2JHoE4ORud4L3pnDgThWu7H4DKpvuuu4/ZbhRsRY381Ors1
G09Rwjy1uQhIgDl8DA2WnZaLaS14XCqemJC+W7jUvqs4wTxN6++5ORZEY/s4fSH+l9u+Yxk6TZID
gQdXFcs70LDtojQzom6thydw+E5HJF/xiiAkuzRw6s8DH+Fbvn4uz1j4csQuOY2dB1l7qvSdANqs
UMQ5tGYVPrJ+Zl39UAdnFsig/NK6LaVNzahokPMVwyAbysOTEFqQRSgMYGNPFeanzhSO4We6ly/B
6i83Ck4w3N0+o2k8RlA7D6jpYxU1QfHX270i3VjJf0gBjEVPbDH2v4ftt2nUxX0hsjeE9Sc3v4w6
SM83JcJML/iqtDIJPljJn+1uILrFhRRrxSuvBWTI2CNHE0wINKpwLFxA4D9nz0ygo8JeSALjkoY4
3o06h8NOMoYq6o9uALc0iXwLWs5+vR3deokbBSlBkC9QZwYnEzrpnsX71D++UyONYQIXUE4Vpd8/
4e7y8Is/AYAgyBtFOymdYwGyfZKLFqOdpNp2GSRpuLiBeqBX/rNWQBOZq7/r+mla3S4GTjMJcAR+
/qYcD828iKML7f82ObKRuqvKbWaDkXin7cYiIsNPDwkWvVfpCUYZh2yvMTg8bd9ngNpGbzX5xqfB
mQkIyT1twjrCBGvX/BeEor8mhpfkmgri2Bf52eD6frp52FhNx5fQDYzisw9IdlTQrXsmCkKYfgWQ
vxHc97TJUHV15uNbWd/FcV9PqMcivae4GSaE9KhUU6+xpL9hm4GnqymSHkPOqzaxdot0Sf1B4CgQ
8dSMF/8EJvviuSGELSV5kf6Lgx/11vuflqUbj+YeRIDLWvO1xlJWg3klleLQbnWe+dTfDjHcTP2o
9VIXLYmQkOcKu0DlAvql5IVJ5kUNv0JCGwtrT79d5UODuk+UqAW2lgADlv+qGRpKnZ2py1z5UiyK
haeDpzluHjAnF7hubJfqHjuTh/3PZckDrVMtsTMk4p/cj4iY1R06MX+apCN274E55rUHP2Ci2CsW
XnN+21Co0OmVIeVgqsai6C12R7NU/lxPO+nR05DDw7dVn4qS1S5knDkdyWitHIX87XdmbPII6a4/
XIEhm97N5ND27TdliU9UtMl5r5tmaOiQn9WSh4U7giOwGpCNaIWiX0x6ZK0mFilRSdqDEfvmSOgR
U6NrJ3BAhf+wJoGBF+JbchkmJqc2vw+qKpXG71N2jviP3n10yn9JZSByDAdUl0NJbCJ84K5sM8vv
raKRD5EFP1uOJa+8ntgt0RUbUKdQYzLeZJ8C0Rv8xyE2juGmseGUefw+sqgrP8wcntig4YIk1wDI
kDUSECJS8ON+IwpaH/QS7KtAunkDzuhMHlE3gEq+zSLs/I5uLjWzroYkfsSy+vBJCPc+Jx91Lt77
JoA3yGxhdxalMoyb8gGybE+LJXeKBbGetyYDa3qH33RiJDyNcgXixz7cYDKZGj6g/lAWCE3xRC4m
ZnJRnHckuy3Cf+NyV7TkUOtMAcTcDKNvaMuIvIbgP9cBb4e3UpPcMJcP5jhrQ/v50JXI34CNg0qR
oqjhfwhum0MEwNBOn4SuhwMmyqtiJAxQ4yaoe+zTAwS982z9mVWPGWkxunmJotplj6U01+r6WNeG
u19by/HYtEATBXTokxjnfl7AljDpkR9S6V7MK8rTBzSECIldNqfXR7Aoec4GPeDGIMcUIEtls6nP
KNtId59c4s/jYBQmNkI39j0cqkFvGCPJnvRlCRwgpmJyaMAT0gpo4WuMve4DCXImX93C0ukwY2cN
B4Saf1dJydPyVbDE5empbxrfXaDKeSB5gmcw0tSmeGf+RLdvBGxpU42Kl0HKNhDgVR/g6+KqLEwt
ckpQBlvvJ4gHwezI6B9WmnchNyFfE7YGJSYxsHXBRgzaXUlZ5DQGzq+KeDerWPRzOeBfqSzDFvuy
fuR0uLwrVIOAbH+Oeb/6GR56iIc3y8N7PB2CK0eLv4w/XlPpGvXAhr47Gengiwg0DoXV9aMMUZeg
GA4aR/+taIOX1FemFuoVIVw0LrLqPOtOWd54zUOZScTJXgA6IBYI2ksBXnivV9j21l5hHf84S2Oa
USDVgDZ9QnlQBmP96XImVf04HRratJgxXS+GTcYxExk8uupO3Q6Cf83pyF3VwgYIIfdjFkK+92Hz
YK1dqcfeXYGK2p/5YIAkuF5AG5WawllKYysxWmWxKqBQQ7sOjNUxawFEVJYhtpL/aP7qvyqxR8EG
vBu02payUGSeK5suhhUHmJtcP1BLcBcfi2WzbfU/z4V71rGL6R2biLGMN5qVMM0kzqcpOpMgMNGe
1PV1Jf+8kL+lLn/jzf6ePDcko5fmcMX6RgMN2Zz/gFMo7CSkbTFOy9S+HNAp5WmZCkwPAH+erST4
hQnSAAvKpOo93+6fCa8S6nhbMvDzNbxYIN8jolxX/nqAtfH8MuTYRwSYE5g4OFnbllIrdsw0Sddo
xQuIyK9RJFP4N251cQO64m2lh3sEOUdrMT7BiAUt3tkIxhPCyZxW0zzNCurnFWD9kgdHYLCzZc0A
qZHOhOSoS0Xr9rCNHIgT4dmkqfTSbNJscNX9fWuKowRtN6vIRMLj+/xu7/YDC1qYzWPnhcmGrBp8
0a2tRUD9+fkJWAolwctJRr8uX321VKEf4Htz+E03SXMa/EQNcPrDaaYt/TSU2mAji+pFYAb8R2uQ
+iOS6dwbwvNn9XqzzzxJpqy3imrdhNtcyjSpf1atpx3xLZ/bcLzcLyYHa2OIgVVJ1MY8G0zz38wE
byI5sJAb8MCJRY51hhnLGvRyCHBSJVOjvd9jYbz/TgGfa3sgRi2YX+9jBFGMvPDRS9oTzZJvrUnL
OvtJIlulLwNsfuS0VnvWyrSQMxXD7/oRqgK2Xi3OCH/q1R01e8cRrQD21Sz/qp5a4szyik4dGIkr
J+ezyxgm0cXE0q2i8V2DyjwMW9zk5qslUHYSy5o6h9Re36p0ja+BPC1CZGVZVEsn2YwUnd/e82m2
bKBIVaRmY99NkD0lWFxPahdwGAIXawgaHf0sA30Tx6c+aQt+IpG6l06D4KcofEay/JMNRJwVe9aB
Du4qvN3W8bbxYfKpm8/K47F4CeDREk4xbSwaSI8YoQv+5VXasNw0DeuBultTmnYqRU8oyZO4E8HN
Eo31YoCobOjRBLo7bldqyyCpeD4Fp6YSwSItf+5wZA4a38ifspnnvBfj3XNMZEI7E0x7zZFg86+R
Zt6ZRXixBdaMKSXxpR70BB+ZZOxLLM6SN3AarP85SRhQJRXV5/XokJDfjjplVK6zwjaUmwj4bh4s
FyuEySyNOt3wXDVCSCiCo/BZmUp+SY6TDJbf/6SwXJK6nSuEPT43tJxQvUTVSJc1iIZAe9SGA6ij
m6CY+Ej8LK6a8TS/qmHEaR2g5PXYCSIu+zwn/f2/hIrGK7Nfm/28FUwsMkwaJGkWhyCPbwokFnIZ
D5ijrefnzN1VyPSQ3YW0MoJKgGOCx+29EaxAcVqwSrJM91fqzlzuVqzI9fbB1btC4dcav+i1A6kL
/ts1tkU1KFS53mDqbAL5dcqYS2yWN0EetHuF+N/TRcAC4Q/K7QHn7sWMq83g2A+SdrYGSyMCEZ8V
f0bsHRhWybZMyXaFrfpNY/URb7ubmu8IRXzb1110v9U41KThI8uyUcuRrx/EuOQsAOQJ8XY/AX0N
6hIgAPdsIj8ZxJNKXlq+lHKihaEMK6KNv6PhXJgpmgGdTvWbAHXFojXarFKJ0hz7Cgpp0g/KKKkX
GRSklA4dlVr4+faFFOoEmq8JgPl8wahNCQvlbt0Uy0CYp0AFToy5H1wiabHClOXmUQJYvOWzWWGG
Dwn9V56tw6z6oMJQCUfTj6SbzBuEPygckIBAveUuenCgaGu+GXgdl3Ez2+A6hvzeJIADqvrDB01c
Zc1IJHPuoGtV1bqWK3aL//Kkatpot8m7FDEkmpc8XYmMdoKiUEz40SMbVdl8quIRo9LfmwwfZs/C
NHduPJijVCyTR7aG3x+OimMkSldbIOR8PqVkouJpMuGytafhvSNMy03YnbWH952ivPflKWFce/wN
m+6F++PANsgGG8Bw/qP/pbdJOM7Jkkk/U6axJhvvOJncKcX2oM3QzJYDAN6R8Co6PaP8yUG+rf8w
ozRBjhjPuxG27RTJQkP7ZB4X1LszLxlIanIUqmpNstw9oUWc4/0B8n589pp55gquCNNG+bmP23zY
7q3qV6x3vQ7msZ25BUh7npwKtdFC06YqE4Swj/U3EZD4Cdw8eXoyRbuzYsuY3RjLd28J7D00Fnsc
8DEUNZzUmlqFM+iHZJzzErPmfrPSF106Ps4zS2UDKzhUG3SNPbV7/M7Tz9uiUbqoM6tF8u4r+DWm
HgEKbXQxnBvp4adboKO/56KOD3KoITSbtLEYMC1yyoz+SkbPao4OElIFjQa8tTeeHn/IcK8Cd2VV
Yfl6NqFyc4ux0sLsE8wKB/5FtZty7/UFWZgeiLBbvmLgajnfpUlhNSsU8tKlrB4zAgLZ/vRHv/KM
bkznDSY9W42PdoqxIkn8WaL28L4QpXNRzKfkXBDrbZU1uY0QhliBVl1aqFg1/eUhxb60lw5WK7w5
9eYhs6R0je9ATObvap960BoFJUGigZKiUHvbQYqQTqkh89I6Gj55xxklYovNRJi7PR5AK/uRehzI
UF0W4oXM13v3rLpMOIHpXibrsAJQca4t698SIFeuZnnPVHzruoAydZaCIhbD1un7+xp2Hred/KaP
IomhUUN4ZYSKrkh1BfWaY4BWkdikmqumEW9IoJOz9pppJ9Moo5G+YU9zo7N20Bw9dp4yccp3I9MM
E7MPyigLPNZx+9NtmTQdx6j5ntx5OR4suGbbJiqwiNxgv0PiJu+tBSYN88D5VLUg2+lUjDDbZf6l
UlTj10199IcDK7ozTuI83v0GXDxfp7Xs42hJ/r56U32eFituxewvN6wo86AvJe3U6454gS0E4FRE
njoj6Ko27d63aM0Sj3ZtRQm9WKftxfUdF3CYfhKWJUUiRS5S23bM8gR8POsVtJ9TU2ApFZwkyLng
hcxAwMzC/am9E3rrZTBK2YASPKG+h+xvgMBnGVZ45UEbidADnKxopWX8aBF1DRVL2F4qt2K8mHFw
COCLKhTSyVPAevuFLHHZQwM/fx2T6kNEs6TTNxrq4xCHb6W/gJLrF2kAS31tiCp36aEjABVYEI2H
vnmzk/OD6H+vHUr53K2cJUu279/JPltTYANOkxabsl5MXD3ArL2OG+BeUw2Gb4hwPyZg0ZnpFCEg
7iElFlzaEO+ihVS5i9i4fG7XpkhFb0VgQDvKvXmzw6E1RC6GJnKcPrnP966CBaYHZZoTaHeKnCCA
XvFaiKu+4h7N8/omKz0PqEXdq4PX6mA6CXhHTj3IPkRM0gfreaU3DR+MTg2ZzbFzyzBpeAbZp5sq
2C8lDzB7nDXA4L9yXevijSvSgyqB6bpsYjPZlO+3jW1SKDhQWi8eYsn5nv2A7HX8bh/h5JNDQ+DO
b2UtVo3ZqGTUu97D6mF9sVeQd2UXxcRESxvaMGr/4HxqE2UefDGhpCRAKq9KQPpN6+6AHHwiVmiJ
hM+Qe1ICfXbOd+nDJQ6gOXC6A+U60RSLLlCfzp8lQN4DmHv8F7+9LmGC5qHAGTma/7eVoIt2YprP
OzmOGAw24tRqI/OLq2zHedPSA04x0+D64xhh2YNMw9ZHhfD1jKBUpcNiesqvbDEqbDAqZvtUC3DY
Y52zCtOFT41PjzM9TT3DBRhUUS/cN/nAcfOd3OQdUZPMmC45qlov/cVp8Plz1dXvWmdrFbn7p5Th
i2FX1E9mYtKs+ETYtuBDWq1vMPVfBhnoG58BG1AfHBNFD8xgn0ky6p4qsCHwubPrWL4rzm9Fo45q
QKBMk82oS5ish8f9bBPjO8U25HO8CuB291FCOoATnDiX0HeQxRQXWksidHsR8ehLuroRh+kfSdWs
I3C1v2jxbQMLswCwo0BZbQWmayQthFemmuZu3DIlmvr88sA51AaKygzrPgLtE3twhXzdoGE7+hXA
VnjOTSc382GI4t//yIFg78/zkag63qQqojJflEjEjs/uaalbqR2KSi6qlCDStRF4khMAejk9yzXf
d/Bk+u6JiywdRk1ASvoLRkNdoNXHZqR+oW+cQXqaE0I6vddJijEcrf2v66l+OHT+QhDZCyXVdh25
mWBdFtDJs4TdsH9r6HvdkHf5GCHLw7/zVz6XtC/8IjZDXiYTCqO5EQQ64Ng8YE8obMT9bamgbGCg
8t8MIcYiyTus6LitQgh3795CDl00VQO6ZBKX3vBHnJ8I46t6ie+ZkzRjFZthvfNLiBxGXzMcbKA7
xHzuj8xPXzbZ+q1orPG96juqQ/AbWMWjF/P/z8Kt+ic3cXLknQH1KEW58qCkvCOrWLQeLtQxR6hr
Aoa8Lp8yEP75SOpdZLiIs0gEv2TId2hpneJLBJtOaON9ke+Clw56IU+Lnw4FpJApUPwghNgqwGGz
xy6lf4Fpjf3U9v3piYA7JmolkoisXbazDZY8twvXlZ8u6sxVKpShw0GI8sXdMneHr33UxB3k7CJx
nhFgDSfeB5e4T30tWTQ3OmjNoYqEOVZSIwPMrJAWjIprZKE3XzOO04iRBt+HpocJnu5iQgYgVY3G
ZcFZHImVnTOA3hUfW4wWoA4wErdUc4MNsLYxj2+i/iBVbvJYa8PWaX5ZRn27n0FS5fk2d1NWMKf6
lhiERfZh6TwwQiQ6PocSsS5qIcjBSDG11jXwZ5YMCVFow0HiBXpcSTxlhTBvJnjGEXCb8z8U1eEj
dbhuDWuy/F2svbnPvuw/LeIKmLMFQ/ocN27MT2LN/sRIPBwHQHeAqfL0AGkYVqcQGk7UIYGILidK
Q8EuNLA6XjBWWTc41ZYMdQ5O6OcJHOou6rzwBg2VNsIjaJL80R81ON/vxL7vRLJtZEuyia7pDVUd
9dsGqCSDrp6qWUZFkJ3sjZ2k+NSgz5I4rhPvwkdbgyh7QIIteVibI/nSrXYstNUm8WDbgSnFgvMR
HF2d/fosWoW7bTN9yeh1jYI+OpSBzCIvR955eTDQElb1unCLu9NZkaTTt+xaq0fZtaWsb/GdtFzN
ZKZN56BVbYo+B9CGqRBTJ1Jc6UOTa8zmQAawCLuj5QPmN9k6wl/mz0Ty44vkx7ago6/w0i4/fF0F
+LIvKWvol3+ZXOJVtklNB6O1S5Of1ROYS60EjDS+gvmKHUJd9sF7KJkDBRpCT3/RrmY/Vjb1N/N1
4V5ARIAE4/2+ji/5OaZEQBrsLJTEQRO/YDVipPgPspnQhoG7olNH2weTFuw39m8PefXXxB1jxlxk
nmJ0ydyg3pc+ZqbjBTEDXmsWTJ2IkKOIgJCnd4TMYaa2R/u/i4RvfrED8kUtKELMZGXdTX3nJYGY
yiLjUfrpAofcrEA79MNxhrOivC30OIOVKiEhZiMkhnqs42kwiPGSTQOnWCVHLTF0OWykdlNbgulv
Gp6JDgaQd2l2fsJrmnXSMnUpTZYjRlgwAsnrUXokqJOQisGBBi5ImX8ChtMsHSxfvUeqb4uVjNYr
sxsB9htoeIjNYvcEe7Nz8Trmi2ekfc9RkhvJEj/BOblLcFW8Yp/xel9P4hGdmxj+nQgj1o+q3V5w
s/Qhbq/BxKTw7+R27+Ex5wUIY9HVFB+pE5Y3U7uPbQO7vwfg+fJSE4EvIqSjY2CScVclnTIXd2io
afIOi7X4Ttyt6rBQD3EnWPHMiziZr9k1T7hKrTESO+3bdugTfPUxnZ2+Ar1SrV1vxIoA4xt6NyqC
s9kHATjTbKzp6HFUJuUkM1pkzFuugJNIMBk4OTkALokpnvx9yiPcKYSw9cEa91X1Lwi3+niR5fKG
uYFto4XhcZ9/lo7ycIHAGs+0c0/xW4wZobc9MO260rVEMeUp7sTO50VG+EhmVl2/deC2pY3xrv0c
y3Lf6ABLDAxiVxdkXgbxH2aYeVLyXZ4pKDaXzU7BxdgDqvQUyg/pbFoxc6hvPNrwzccnRXYsOZrF
bObftK4+pHV+khm+kdSSkkYp10ZcNgchzB+ArutKZMF62llGwAZk3zxDfM/5ESzVYtM7NaJehgsc
TMZ6sS2abdFKSyc97l7f7GvPgDFSBNiSRzrFmn5cZPh6CJA4/zXn3LsCsjYk+1ZfFKzsJhvyKotf
B50vjgdwXqb0SUioXoVMJDiZkJom0PeCQEyhEXf3v7akRAw7MgkL87K5C4kT6vT9LSYd8j66WFPH
LcSZ/H0kwSq+ukttaJZaUnK89k3NBB5UY7vha+bGXedw7zbQCVK61cyS/+xYzF6Ry9KIpeRcBoyw
QZFPnyRKBLB4tJHSxez6zzZ1mrqPGXfER2I6dMzF3W/YZwN8Wa/8JLx5B2Vpr7JHIloNx9yx6asN
2nSH+qX1F9RGLQn1q4LQqwuSFLHQbyM/vBk9t6M2cNoA9PGK3W2PKuHFxIRnnf7haa5PUu1FgvWm
MJ1cnh7PY2WRMAp4OnaSrSLwZ5HA/vlWQPoLR52W9Sr3kBKoeOu3hlRPaUxZJ7+742+L/WjFLg1/
GnvHQvfQgrI74maq9UImTl5+6czHoWJbFQiC3b2lpfz0R1tfgEONeVr3+xMkf6aHSQVOOhHcvnaA
gPpf4EgC3yZ+0VEIGHo5BSvROwg+yOU02E1dY6Pg/ib4Vfg9zZdra95DVeLxiOobT5ZlAs4ZuQW6
kpi87t+bmt0zoQHFtsEB5sH0RA6kjAv7vpBmYBDdPQDpJbdq1F2H9i20AjQWaBTo+iKSWbljSXwP
AaXqcgYW+5w9/Ewim/zKhbzeA9k8Pg3FBID9HQWImk6FNWG20eEbhL0cnWCj2l40rn/KhsuCsuHc
T8jn42sIRJxOXkAI19ZHAF43hLnNRH0QafuOsj0u/9inVn9Vuo2z7hzFMlci3LR+5orK4GcvMgen
/BYzIIai9wvILmzc0gykmYvgC9KiEOLHX8fLu67rvMwl2P6LqK6VQdivUkoT7jvUeDKMlhPCcyJs
RaYftWSSyFapw+4X9/6c38PznDfjDYVnKKkUCza0dPAmdWRJeM8aXOHPc1hzxF6Tib9wasYUQIAb
0eGv1dXHENcIkQnGyzkONHfsFjw8iUY67oXQQ30cuFwz6RWb3IqUr3eDQe8LwxrmPadIv1CPVXtY
yXEfWXJ65exIVSRAXYbpn9xpEohBh6vKFkn7U7rIHz0qEeajxjLKLNrjc9zWo0hEZkD7PpQiTzlL
Hd4TfCW5AhK1x2d2lR/fr0W1NSJvJgDGyxKtX6arJUxm0e1Za8A/tf7qflSnUsPjuuGurXTuhOei
/k1lbfeoE9F+soBT4nAK4/HRocB+ZYYFrWQpQnsxsW9gkPCj/Fy2GVr+ePxDvjPBfqQ1MUiZ7ptf
G4YBeolgmczsZ1stxI8kpEo2zp0b1UTFSBhFgxyLgv43AOURMWbTgIcP8tJxVEbGHeviyDGR0trm
IO/lmC1ktFYxzF0/KdPeLQrfoG5LZ6QaERLuJwhlcMkEHz58f0L7IwSR77hV4xJkCMikEnkbNetK
h+l4PNdnwdJqDY9fLQfq3FI8bdb8H36HPEG+gTRh10sOLuehBLmiiQBWyoXzy9EETJoH4P4gVOqp
Egy/vjC1ZaV1d7cPBd69j8jtWPYGb/9Tsy4dOWoEv3xy2V+VFdLKTcOq8eHFdJ1Em2YM7pOBneGu
X1pd4bKhAeCjSXVaYe/vnc2BRUcm4byeEDBtC58/PqPMEmg2a9D2Si+DTZKVCkWDGQojJxpuH5X3
wzTBtYtI2dDheixfGw30nBA2DMSxgWIAu4iYzOjPB5h4tyDzJyRugrQfkzE3kRigXF8A7cy56rlA
P9JrRvP1BxY4DtCq4iyn92a6lAn0mgypXv54STGpw3xyG9eV1N4Fh/Lgw8zCUTGTDdlxQoTy6ixd
kWfyEMhQ7fTUa6rtaYDIWKPzPfOzHhHwq9+8cZlH3If2kn8MFSxrNQ2bI7gaVhDISTxFi6yn40LQ
W9t6Q9NRE82TxUjBl+874oEXHBhlAMClZSJ5QNKzdXqsbEI/kxwXjw+39myjdTknP97HZkD8MhoN
dyut6FWUrk/02ldU/A5SXfj0TNwsQ7WA2P7xbqt/3DM3e769WPG83tQ2FFgPzofzRMDZoUykxQ7n
C7awPCP1fdywhDStC6gaNHV/kUQ69tEVib9V8LQSINhbxe6OrTxsueIERt7g8M0slLiJ0+MiQBQi
OHE2eXAUE2bt0gmA+d0whHtlNiZHngHUlrINoOUnx1MeuuLXZ/r5lr/jAtalXtXHTA16RpVvKz5E
LyWPfCupbnEgFQVqa/xFYzeDkIiNVIJz34XBvhByBLItYWsqR3spkQRcSwQrtLWycMTe9/gvdoeW
Q/Kro4B4n9bGesdr9Kb3W3vZKHBAxAd36k3eXdXUVfFdQdAoNxupeIuJ2wZKdBsOAHQF7JrPdyal
+IqtlSll59pz/y3V89vCoWRk0GCqA9NvrvOR6NhyBk2NmzYFNUQewGF53dRHzekfM45w8HVLydas
eRgUSlBiK/8an01g3OMDikdstUaVdJhDeJFM/IVULMNlwsIdAsryB6B0+FksfcGWioH93Svmodbu
p7hnmVZFDMJmJ4z3vSNOh3A7B2BzL3uiBQToqUfM1Dca802XJE4UumhabegaaRM7j6qyvggIzX57
crehVEzEE41AWTNDHQ+MFtDIWchapxdKZMEcBgj0doVDRSJAkoXOVSCqdD1dY8BgZzkbcDYXP+YU
aKKWnCZuH+ybvat3uBzt5k4w7EJyg74Eba2S8IHqdb92V3FyTeWJh9bol/kB0V8rZvgqjp8IxGa8
s0NGUnvJAkuIS2XTRtiFM8LfQv5n+m+dwOFzhbLh8g+iioaUbD9iYIGM/+tbW6kMqmHilg3ULjHW
brkkM313qc/UYg9Kdmanw7LvksvXAY2Oqo1nqQoyaDocL4wA0Cvq8GBGq1r65hZu0sNj8nNTMexB
u1GyG5++Tiek+Kp08XrQb2WZC3TsZevwIwi9NyLdl0SQaGn5Kmoyj3qVFiZPWDPLbrXjQ32KbY6c
WSmSonlg0XyAVPPrrnvS21mz63w1Qnnzkw/31GjwgUSkOx5i+L1C21SpfXvfuDyfwgMLCc7iSxhM
dmzH+s+4Q2KM5mfR88dG9Pw+ir3bC9w7DpE+/17qNsZP5UTg7AdkUDLmZ6vDNs11ZphSwztXI6Op
wtrWbfSk5ba2Fz047ABPY8kXntc89uHoDPnduJbq8vVhAYzFoHOaoSYDPomBwjSEDU1iu4P3MsX6
9Vm+FjI3b364rhANE/qFiih9FQOuGmP5jqo4VHFD/+101520zW7WzCpHGlDiWZwdV/dwNFQ+y6NX
TQpI23AFJ86CnJqyFRKGIkI/exATdptjDNqeMAUg0vU72vp9JppW40oqGXMRZaN3AqLfIqxKWhbI
TRXnnTUYDpZr576Ph7uOLyyXijVITwQgDRhmpMJ3x+Fz+HWqHF39YhzdTl3wcYx0KdnPcBry2vaq
2RmbB0QPe7g40f5a/HcJZAq9AB1vBk2k4rg1MhUKCSMP+lpwJ5obhjanUijpRJwKhP/W6zuR5+/p
B/rmApZRSSxs5BhsyhkD0nkVxvgmbr4p+RJhWgL0DCDy3ZFlOgTDA/qUNcJQ+M8dQ8kKYU9wLda+
tC/gktnBVBWcraOtLomKaglyQydzXdM2CkEXXapJVoH8WiyN04fIPwLsn1AKhYhvB8J708zvFkJ1
uogkryKhz3eQcrrGzhCwHioT/IaglT4CCOUoVDYB6ILqkJe5fp2Y2qKKzRsXer51ewIYR1+uerWp
Dsw5s4mrzOQxTNdPFa8dP5keW+m1TQDJBzHF4p0cfRwvQhfCJhDHpAdXzGZzicqPEENfudEdxf2C
5nuVoNoyS4de//Qda/BNHC/2S5If/4Q+dcDLx2gpoewLRwk+rEaFGmz5qwT0m9BWSpW5bDE/CNxL
DvcgK0rNLP5y3PsVwidj1CjZBo8tRMF9I03tcIJ9J3bHygC7jSR0CBM7yoW4otGCVNuYR/nSIEV3
/q2vLHrWuVhs9UZv0aZcg7lJ7eLlWiBGm1Lldij6yBT2m3WcXwEOtbNw8EUmIXUhN4aSG46oS0p0
swa3gSLfBKYlatpjscEnES9yEK4mp6ISuEnXYt6PZDlhEpow8FeWTJb03tsjGlIHarbv2rMPxsF+
3mdQMGpyGkBZ87KkWV2VhdZtiBPHx/g5PWOeeggbnZM6Y41IOqb0cYWwDrDuO+n7qDDuL79D6yqZ
U/loMRsWs+QAG+KlzX2Z/KcrUwQqQp2GdS8jg+VocIogrGXxpC2+P1QFBW3N3gVCQq4mqwes8ycC
NqqKVZpp94M9SwjxBZxZ3gnY3hDdy6F7k2pxg7HUfN03OXUdfk+aQ5bbe6Zy0kE8DTzJX6hDOh/H
ai6LQfjVFtTpQOiemq+vc0CoFFu6Nn9YG3jOdQ6ABas+ckjA9Y2Bp/ButsI4mUxsz0VhVRrpurQ0
Yu0EG65EmjJl4/o5VidvPPka+jOB75i+EPOTfTyXbCoSd8g7n2vXlSIf6aVrUbdC81IbpItGNF35
Owpyoick3BLHJ4umBl6VJ1Z4akn/N0AiF7UAZWei5u7QSN7436CV9U6j2tadACMWJ7eP4t+1Ae1N
1QP6mFgmu9iofUg2j7gtcSFcHub4cTQ+YWI19STa9mHXQaVxRdjUQxXeO7H54a95WaJvjJDbFkX3
3ZAV11TOlRjrn5MFVpiYzrTlz4O/24vTYmAt7DkUrDJ4J4hsb40IVVC61rakdI3r25jV2gDgcEEY
bkBpxp8kgovGe/jTHv2VcFloAdDPEO/Z2c7CAtHhtFhp1lcgnBjeOfmjH6r7QZQnZddXwYndodHi
QwS/3NqJ209BZLZyDR4v+qPS4BZaFiHzVaqYgesIYPZCmfzBwDdxytbDwxetQFxyFahzyiuUwGMp
ufar3VTX78/3vMkSNuOUb5bECqyqeWOSsjyVM8DO1tOgf51I/SRHZg51x66XagSxitkY9P+yBYVy
nPTjbMgz2wbvW90DEDakoAMR8nfznhCBZkJMavEyLsSCb/a5f1ba64Og1RP0hKbcVp5Qv6Xh1WBt
Km0kLrDvys8Udn1kzW7sVJjbUbXxixJ1TuRNX5/7pwl2xfyf4Oxa0bcBJnrr7Y5aRrkC+hi6SyfW
m49Ju+IlNtIQJw4BG9XL4ZBNIn9BLlXlr1g3p73pMg2zYKCyzX7evSbUNIkscJ1O9FoDe8iFv52W
6CwITWXX4PtuJLV0IV5mk8AmeM6rfY3gjCR4HGnyrLuN59b1RcRnUyB8QP+B6ydG3iS79szpjPpt
iW1/oW3zi82wvGuRnguQjh2/DN6D5I1bTH+qJLm2d3jlM7blWoG/gcrybw7wWBGEPH0upR1mwiyK
X8ud9mH5JjwTvLalH+wyFycR5OfodjxTJ+3cRKIuRMm662OICfmSYSYtUVtp7WGkU1Kd3/LKc/pj
bFKQfv4BISPdGMQ5CMcS+etghixdzYIK1E6eOCoVN0TQt0hcA2+mGYwGhhowZHd3GIyTG1K36lXs
yu+pp6PFFOKFR1HJI77sTMq62o82ZDmtSOVR75ddRsD311iHJabLDh3yI9mXdFkIlqn9Cu0A32pt
60tCcN7w4d+mTqErxRiMEGDmc3Z9LofjZonGPEGoy+x+Lz8Ag20Skbhd7m76vUQcfWpKeWfa3ylh
+HjKxBbjW16p0S0sCRIcMB70tT4+iFR9iX5MOY/YlMXNAAp1htq0jSIfyaa0ffRxoB+SDmFYEOqB
DSemJKzg5JJ9cBO6vvjRAtaX7VBnBJgsPzNSP0t9J/O81yTrPzfIWZ2TXPle3EIjn4CHOWn8xjxN
LZqWZElOyw4IA/QCH+TH3nSKYRNpYU5GThyvBtDZvchukQPD7KD5yVbLPiA8CAKgNbiTHe5Lw7vB
QjSOVHqktHiYp8P2H71SpxIEI2s8EPuyeyJk9vwX6xg+apKE2H+ZQYfetKcrZ4v/x2Z3eR3mCCoJ
2Jm+f/DobwjSd+qu32ouZMzBOaC4ONRrFoaKhS+y2YK0a7Gp0N+Qvf3bHsheISPZXjhUKaUbgnhv
DcOcKrljr62ShngnIlDH25yVfNlvNcq+WlMyFjACzVAeHQMfbNRf3swMtexst2BrKN4s06lwENrl
JEEO+EQGUUXmUEhqB2/q4gZ9uokmhtdvdP4fCgLJvjXpECQ3KDQ3kLV/IMCVTjZmEu/yBMgMd+WD
k/1slliidbxUhbsgGkcJuItEpf34ensnDnHpbSyil4HNUSbPEYdpyT2+D3Zd5exNV2ffCV8kCUeq
4BunddhudKw+yPkX6DOYCgo5Clms6tcbM4qtWOhZD6GvLh5siKcUe7n5GuCWhtdDJ8sPqSsZTVEA
UfsmnYwu5rBOYGI99/AfTdDp+dllQ2AKaVkBPncDg6cuCSN6iU2uMeloPdS6UD+LZY9HD14OJgW/
BBJxl5EeeDZEWKZymyIts781CEvYUAUtlINcE1tf+UluceB9FFSVLpwQO1ayT18yc/wqhlDBKs5O
f2bVATFIui3crTqa/siyjjx4sogFX6R8KeP+Zm04raBLQvOsS83sAzaCOyHDw3TfUalhpBTIYNdh
dDPMDZdTCIsKz60TW6SyWlhm3ptN1Bd8eszk/txjqQ8uidvfjQwY/2mnTWi6jUaoQLKgkKWDq2TK
JXjWAJp+u4DQDp9k1ZNVSvMUlQEEFFaTfnYGnRrE3RcJZKtf8M0mHW8X2VtVuOYiN50bi7x8zvAz
cLg3aS494aaoSNURlROt8+Wrx31SutakFlpni5DfGJoBe6jMHHg6y7/LMMysvO73GemMJqv1QmFk
x0JI267BLnS70M1VH1STwWZujkQfulLhOxwwCkV3XKS74RC42c+VGQi+pvKObmR3T/uHapInY75k
Fygoy0TrhizfVj8EG6qLkSPZAdB6/9UnOSfjXP8aqDTGcsRvtrSYbAmvXTSOECKlT118CET0oSJM
DHtWjntHBFZQRsILoxlCSX9oOpZbl7A9aH12Q6hLiORDpnbeuS2e9ECdfkpj4/tfJplkWOUllRum
zFwSo7P+Ro4tmr3pnXOoq0ez+btUo8c8p68q4QMyWY5Np/u5nZ/sGK3N3uXWp/9PIxLpWz//5mlz
0OaH4R5wTs/ceNGqWbRGKFIhLLk38oH000XrXKy3ECsDh+bDfmuXdR4stF4EJgdrHLpgEx2z77jW
uVmZSblnBk3NYJol6sdP73718BP5m+BcGmH2warYjRqmm1B+IjDLYgLkAj/zjngdaAM2BiJK2f5P
GfL/26AyyRAHheky/OfOXJTq1eoxOb49RfQPvy7lB3IQ3B1tfKrwfj0F0ltnkgMK2dS93ZwnHz3v
c62BNSh1+fV1qAdg8TLfHBGDvCmJ5dAmCBSIDg4/+PPZNklFu1q4qH0MXXMjqaXIhYerqmpR0aJr
pBuIWfW2iOuGCpQEY1J3Q5NgvBTXoM3gMYgwApzCRt4E88itDZlM5A2adE26s0iB4nnNh9VLJN6M
pdWf+gqb6QwwNPnK4beXkzkV/U5xw6xlVEJ1uRCTWLf3BqBpFSB0tYSaJiID/wyIsv9tZGuSwec5
cXveF+vzpLynlYokSxrpQRDOKGvQIaIbH/KakXbbYrqb/7mq/PaGoD1q5Qx7YGsUW3MEZfqqN2/y
o13m0XlNeyx1HCaB0M6Y/9bl9Jo+V247dHQ136w+ui0DofBNL0feh18A6PlZQxASGYGuaetXBSKd
5KWfm2m4wGAJ2Ov6e3m569lTxKOvfJIrVQ0cfkHqZ5cFfAnotsO480GeKALGeU8Fio0McNDOztr1
jSer4qdJrBx0ONzZGw1tqBqs41c5CR5Eewczc/Sii/Df03akmrJ56N9ZHGjSj2K1IArGCPAwzsb7
VXUKdiovJEKcjAlDLW4DQ67jq5igisrXIINpeEXlfeZ0c3NLwqO0x9lwQFb0jJDStumFcwubLEwr
va9rYBtCEri1MAAluQ+nAgXC16kL/JUrI8FYDcNoPOcKiz6RBBNZ9fWjTFPVgn3w30BRfjc0TmIv
GAMJOnSBMLujh6v2wwabneGP6p4Rgz4t9QqnzneIK0UvQr4njZT1Rfv8q3o+bNxDPLFQ1OwX8YJ3
FXUtoMBIuaTTd9MPeXfU+Tv/ezicFLVC1R6Sp3xi971Ug4TwRCIyp2154UFfSEqS0UAS2KjCOPuG
cyWEEp1QnlBMXpXTJWzo+IN/jFKnNc0HnvIQ/L5/407g/hW0wdDNaCtA0ytViRjaMiKQBNhzNpQg
ah/X0e8M+iGd0z1US+qrBBoIeXSawoDUxyCWkxeowxika7ezbfssMTTSxTY8CV7jgGdnUAvSOdUu
VvBI8oj9HziXQQWrRaqKVWVGN/myAiwZSFKu+dWnQyCN3OxovDji5GSBzZNZOdV8zm9KENIKdWnd
LhcbdhSunHijZ7mVvWjoTOxfGB/iOx8YkxFs5Dy7Ie34tJTLoK3F6UB7IKvS+pP7nY262+7Fg5FY
PmLkm4/kq0xndrUk7+Z7NFO5D3Q7dBnrxIYwmJsYXILF12DeI9oxB+Yy8BZo0/maWs+1EvjXfC7+
ZNq/zn49O119kI99rRVnGBdcpVP6KYA8kv1IcUJQXzNQDxwk3CJCLDuu/JbalR+5VpyCmi26FYnh
DCGftPJxlmBI33dbp46UrRVMWxYyQZczRCLlWsdXofuP2FuTRgzQEZgFWaTsrxxtsaMOueqZy7fS
gi4zXYlkYk6yrBeMOCMXox9uWvWWnOlgWgP/ShXwgXVihM6NYXpLN5oTuUQjyyAXokVn+8Tble9O
KISFUTIalFo6+tqBmY6iDYxYjRjXQeBiHbBQCi62mCJFUVJEULysWJpI8zGzQUOg2OZITXpC5Hq3
KENvTBCcfoXEW4j4dh4hrzCeIr7KKWfJXCnDLm51hnOhPxHdeLo+9de2V4UMtgnMSwcgF1d1jVmO
u9+ijp9Atw3d/59EW8BDbRRBoT3V8S+81J8DiowsPww9AVU5rHM+azqteEyIpsf2rphSyqXRznvQ
FD60TipEnOTOLQczS0knp/0y1XNQAwXhuCkmAp/NO0sqYZk/bm0zm/iHzKaSwhRQ7Td8saP8g6BK
z7RbnXw4iQ1vMBBcCnDzxryKA4w6WlqxWw1gf0wlglcCE21iwS4MhHtpQ4fm2GCqiO4jFQK8LLb3
4wOcBFZYWxNZGGDc/jwZninD0sqe/tnH1TtR8LSiCPcYsWlUqoXLjahIUSvdE1EG5LMaTSXkCzX6
vOiShIo2S/CbGhz2ZYX7OsZV/GWMqZDUKRTs+fT+L0B2E4qy/bSbJ9+lEAJ1d/egosTn2IGdaicp
zsljdIaJukUK5L5Jln/yjA93zEuOEuQCMrkDWEUqJbeYfy0dsufnOVx5pEkDLIBPWEQE78AlkVx5
MDc1WBzA41Hl2D8i/cpAHraGwAh8yz34sLSDfO9aX+7GiAgC3h5oc6jqE6pZJsOybvWaGo2/Ahdg
e5NaByV5lM82mMIuL7GzMJKxaAjLzbnht2rsz0vMcnqt47i5noSAoP+g0eG2o4dGHsZAkROSfnRm
I7RMBP+ui2BFAwbY43/0PnwIzvcGU1ejwRjDIwIwOIgXVxPXBWXPEI/xa61nY32OYvjc58xQDTsf
j3BLK8wDJ5cM/OFB0yTyAYe8/Zgx5t1CKdGp3k8F97lmmlkOXeQeFVYjXuQJQvl1SFl401IfylXQ
X06sU6HRLmvKtFuilMi7/9IaGmSvl+Xmo4Xkit/NNBe1qxolfP3LXtB9CHxNE/tpw8A9yniRoNh7
FHq51zUGeiaLfaeaAPgIXtK4inNuxnPuJ7p3O7BgepKKUMMOTlJrUPfyucoDZRNr8kf7VF0WDNGu
B6GAFKqUxGXqsotlIwzXb34I9pqIThwPBpSehyh8LoOoDSzrCke2ZUD+OXhqRNaUSsSG4G9G611E
0Ome0grA1fi4lU358N90C3UJyPN1S7zyDPvl6kB8915/3PsN0Q08yE8oMkCrPeYdn0g6AOUB4x30
cL/P+zCuTyApKJ9OZhHmhvGAf+AgUFM5r+D/vd7p1SlQyzRmAcDSuICfrylmTzDCjtzXZvHH2fIL
UT6892u5Mjbh+EKIK4PvY5bUFiAwSCt6D0G0ptqyWaTqdHD8knrxrWnmvwag7q1jx43ty1jDarNM
JCj5hZ91IPU7ell+n6/651WkUHxDVrq5FXu6zc1x+Xs12IzmYvU9bhZSNM0qmxz/e8P8nrxBBwMB
PtY5Mvbsg2MjsbCPOtgOTXBZx65qdNl8hE9Dy4EyZtm6vZWkdw+WjwNs+ATHBL3n1cg02winWs3T
sBYYQx2VYElRuAbclAoNDbdrvgz/oFKgrkvvlSlohYvrKvaGy/maG+hD3trV3znXzhcQatVwUvIZ
N4UqX2o63+IlnWJbDEcNtevUB9GfW65U6Fl6zldcIm805r/MDaCz+dUHGl6W4qDTvV4ZArkS88jT
bJxq5kfs6PsyY7ntUdEub5XmhFaApnRhNsLT8buXRmqmSlcEf7FF+9A33c92Mk3jFD4M3M7YJEeZ
vceXFccNW1bKIESmayY/Py/HVJc+nZGT0ZCW3yEC9tCziWLUX933KsP9VyKzaEnhNKpLNcLcyZRc
PPxmGFCh1nROVGQMphx5n1mk4DzZ85jlFFlhjNTSZhB6Z89IzLyZxH0C9iOyp3vdK6z/0R72P85s
UHS6DCuqt/HbV/dQ6xDn+UTbOz+IRvCUBcRAStKnhv4U9B0uzOmmOVQFLDylqZvgpAMdlK4+Gcl6
agcP8CcfybJuxVtRQnw0eMq9aKEj9xpcyOzUJL+pTNR1LcHPo/FMkUVxPLIoJTIukqEArrd6i4lg
NvhlhiKKSZ/r+8lhpqJ94DiWRgPTHwKaI1RCYKGX/yCdyHtIn+t0Fjv5kSySKkiZr4ZyS3/2I2DE
UZ5aB6Gzd2Ox6C2l0pEWDlPUQdMw5D/eVN4TGPgdAnUg/HZsh3b5eyJlAD82AEapNKinD97ko7HC
+OOmXn7hILEyL5iIStnqQ8I1q+kR6uRW8u7gU234J8+6xPz7Yrg47oQ1lH+cHSex2oVXG0zfdtF1
iWm2vjUfXNhwIT8m0hYlVr/v+w44S1DsA5RoQ6yo+n6CnJIclDX2j9YEUiHJU92Nbd2Tu8SB5uXi
U7wFyorHqmoTc300N77POH5Ps/txsz52MV9IW12iG7pb2dnz4heWhKhvoJ8cG/427etOTv15YJSK
RdK7mx6/EJDUITJnhIMSYCHwwGBd6O3ThjDKz4+EFqT/tBY+FH+tctMf93nNdQgTLmKrZ3QZIunG
t6P4mBAe5C8KPypoxtXpUysyNioylvHsMAfDwUZl9wt18zo6uf7kFbK4TpaOOWl+iLLcUWT+Jg78
GA/yzn8StJvmIv27EXdc8DyQc3pr3OgpuKRbsvAEslS0RTBukCxwG2FS9IlY0btIDeVmLH4sCDR0
rex/fGRUotrDsX+AKNvolP57dVnnrMIOqACg9wHvzy70hNvBIZc9vRRnHWiWgBosH+1cnWmsY6dC
rnutd7dx1x3a0coM6OLPXX2Z2L4D/ssmsU9UI2ICEnD6aTE565ItVJcECuV15wlWU2qm0rP71XTC
Xv7YywNVqCsgl8qP5qmlr27epzuhrRHdAUAMpAJ3FVO1jou8PuP2WPnycN8kwyiG6O/t87NVx9g3
Ff+567w+PuX2zeNbGIgJjf2UjUmvofucCyyOnFLlhi0zGbMP91kgBFPE2N2yKG+eZjAQ7YPLGeoW
sp1v/Ir/x/R9CTj7TiYhFM4QUUEO0zpmqq4D9jiu5H0MDkib4qNUAcy5UESS8tm8hm/208pX0u+q
WiRARviWTDuwEkM+crQBcpvpwEnbFhKArBL6TYi5G0VhSsu7ukpigc2ctbInGPa9ovK3+dyqys9r
VqKYS1RlEThYqUbNf0S/ufsI69qHDiZgyVhluYbwASeJpprxnWgTEBtUOO8Xum6RnIxjC/QPyyKc
Nx3vVL/Lvxb1An/VHci5dunpWJuPGxTtDBMre3CBF1BHKfwHpuhPPPlC7K1aTPY+zanfwWJEA0bO
TVzKQmDO3a41ZAjLMpNRacECr4Uy+m6dNv0FTX75N/5ShHRLyNnbuxeoMUGn1A28G8lyhfF2cn6P
o5ouK0qq6+cvWivOzrwS6y4zGwNubjLre7Q2/FbvaHCjRFNucIVpdnYT6dZljOu3LdO0NoeyDgx/
0+pZQTWvKTpNNz3FnDWVnVaslIBFke1hE+2xo6zMAdrFK08NCFvIjZX1iDz1HG3Q1qG+9IdWgi1S
GN5dWSSRA/esgUWN3t3EPON5mDz+zFt/kWwOFJ6SOj9+znb1rpBb9uQmrEsNCtIe8QcxHK1PkD+v
OcUClNp9OF1laTobEAuMv9vr5AsZCStivUcbc2UhuFFQ9WOpmygSBfxpaA/UYPUdZ6xGYUGBd2ja
VyK2ZFNRqnq3V1QDOKGddsC07ffH2x/ZgqYvux0jTKnvDW3Waw5FhB7QTwurdpEsFkqp5C5mhd34
mmgUm0H9Jy09AnyGmsX/YjSu42APJ+kHHlQ6FOYEz+FTWY1dPrM4wEjKeC1h/g0inzsGZqvmhGil
yY/fJvTrImoGCDMwC6tH2w9c2I9TR4lG5NEJhlP0/UezW4hwaqlB+DuUl32FAKTlIYaY0x80FcTh
PM7cVPYrPHncHJC+Ct221KaE6E9VloFBmX9ku4ktHedb9f0seRRfHT6q1gb8vn4WNwSW/hX/5AHq
3WIH0tZNNZEVAQzsByz+m7m8cu51CM57SPIvrPOotlkIT98qpGws+I7GbdZolgRlyrQG9BGL+mf/
Pxo19iW5FCD/yX9fNmG9pAtqGXNc/qSGwK+ZI+PEnu1LFuru6MoMQoGovEUGJmdFPwUWdAUIeHcP
Z9ss98fHDPu7djPaCxcJhYUNpscv2E6UwQE0CBN0P0jKSNB2XM0FY4hYwCJqYEimfMPQQL9tnW4d
uDxMZPjPaxqjgUprU1ozpFV8epx9NK+r50cYdLGFOlEZ/Q2sqEdTcBdxwi8S18AXI5Bhex6MVtzx
KSwC7WCJFHDk85QQ5GAyXkva6/mKc+ldBlggGRCeyb4Di835yUdFR32FWeXXj0U+fkGBgM7y4pCh
Jh96qzdyHbW/0Lqz05cV+Yj1t0bw9u6+k1mgmfEZI9VXNY4hRL7o9+aQ/essqigDiB75mCcC8IuL
hUxmmPGLOFLJvrYKqLU5S9KnkJpS0iNkLa+dH5YpgACDilPfvtHTIqZ2JIpechamap11VgY6Mwex
PmPZYnwQ670Gm88MJ7ARspGtLHjyxdx6a5OGTG5RFe98J5D7pUIPhuWY2rUUZYaw6UWkVbytpN2t
VRdqGDnGeoPuT11U0KLdq517LeyERHtKA1CJ3iSkOOQAf3OJwMzau6EVH9AbARwCGTCkbBfIA4O0
9U2B+/sbe71DZ0bEVCrZ/zqfdSd+6DTqguRq1Xd6kgPLDjIj0Av6+5Z4KbOqlmNPQOev1Maeimhe
Hhger8+uniEqsadill2Ru/pm4Pyc4nh4uwvB/1V/A39wiJ1/5LWYGjcvZNXN+T8iUbkigAljCZZZ
56SpemxKbjdHhoXzNsfqn7DrkgDp/u6pLzsNj3u23Ae+z3r7E6Pc5Pq9WnrsoBxlbuKNoHd+efRf
/iQvbg2IePDuPkXU9zy8f8q77d/zZWinUReMo0o38KJuBx1LwdankC2fwHYy5R82jycS5+RefV9w
HDwUQGud7E1sA4FaGvvgNSrLgsUppsBlGEZy1AUMUVSK9EoV2/C1vT/NRQ/oCae3pSJC6tVTmKHt
ZwjZvQh5N+7n+HqKnFyKGMDpIfO71XgJeUK9eCfU7LX8Btc+6SEf3DjBGpCCiQlE8gwNu9cY/S79
fLsaPNq00Oc6mdgaHd+Cnzzs5s23yAeQHSgBudJRDhViBy27upLMERoB8bMAYM/Z6NATMPAq2mGB
B1/19yVy+klGbbj4KFqzrYG10ffqKF4oyVh0O/iOc8tUifKiC0Z+6D4hQEFmmINiDfh48b4X1sVX
aI0QxH1x2eMJ+LNdyPdVbPtw1QgFRBIxA0041h/cYo388AatcIi73xr3t4qfQh9SZdJG0Afv8ql1
RD47nJQjC6k83KEIranoexLT5IfHzbdspHXaS7eZscApFvzRPEN7JThVn9DOWAwRDRi2fpsIQdXB
mLs65z04MXnfhF/FvwMq0kxr+l0c7lIyKmYnll9qghzoA3f5Caz+QbhjYoFe9L8Wc/63/de1vJra
T51QyBe0yWWfws7c1lL+kHPkS/cRe501goXtue654x8kWWfOY4CFGJC88rdgXXO+qBS9K6AHrWJI
M8hCHm2A3rVfzjwdepJtklSEz1Q/n9yu28M7vNQ1xVA2jObgr8d517iWOEM9MwkhuozoQM4Z/kKZ
5f+sMTjg6CS+2SpmwWaeqA0Offz90xVbO68N9kcz2EUwQ7o6XaAwR7GZmDl+Rs194n4MMALxV1WR
58hvZ4vxdyBnk26qFGnjV3v+Naxb7oOtGPzDltUXUjtXQoTu6YrbqiXHOpQaY4E3I7P147LmDIeJ
bL6irQA0GEoGKs9uopWIUsfdzfH7ehYXDs9WgBx1NLEDiF81O4Wpr8wv3u3d0oZQyX8dltnBYqQ1
2La4f288FFnO4oXHYdEQGTT7w9F2eCd0laJwt1AI5o1HJQVMnLKzjJc7us8iakVRNa2WiKGuWe+B
bCBEtB9bs44Zdb8xlrv33XwD0ERgHjJBXg41Jw3yGKsW2+0kCJ1IUkf+p/SZpn+SPB48QUyKzdBi
7MEkVuL04F8D6hAlUz9q0FQDf7U8a9VZHVpULwfcoIIUY/IuAWV9ZQLSYeWfbYOnkp6XIDR059nR
nTgDl3jJ6mVbpW9gZtiBYDGYNNO9ylWBLYxoNrDyLl472R7t5GgcGhfw85CQLtDUxFk3pOtKG29B
maUsF/A332mRUcgmMEgS/0/HWjGbIn/CHfgOoVAzxcj3UfDFVFPQrgf0fqeVLBIG5N4/3lK46N7t
TpHMdxKLUefVOVQMRTz1VfX4PdDQb8Q46KiQELM+RtjUkdKRLgOIYiVvbe0FD52H9ECXBHP45eZV
c2sLf06/vSiGP/V/OINkN/JUR5aREpAlj+QCRhyz1jghaYrStSEc2tACClISfCwN+r+7XlhCuLcH
N1NBu49GHOgfRaIRrZ/SyGwVTa4zt42vasXltWiCdfNc+phym/GU0b3rKmOFdW9F0Y2oRTQaWE6j
ZfC66NdflnR3QqBIssCNzT7zyk4KlgorhA5KzAuQ0f+bI4GjNS8bitfobZyCoAl9K6e5+SnXHOjm
rJmyw291qXr/Otrvnb2rPXi/v087too6TmXvU1EyuP6QZXLiybbWrXJZA9O4uoAcOdQWjsW9iEf4
DDkCwrJJ0Tnc52X1PrYs2eGZSmZHkNx6qlGFEO08w0zyhfMlo4uyj00IspM9OavcPfr0QaxsLTrj
sfUf6V9rhTMIdHefcnVWkvoKx1i/OPCbOlWFTreeV+aH+MxYMu3YRE6v69np9W5UfpIzQd8bV1w9
hHcQZftsN8GXMTlNmsRb9GO9qyouVuUSs02zreC3F71m4UBwADBpyxZ9vWQc6Dr3sXgto5vz66Bw
L28+q02VKZr03YBbTtqtlCYNOGxVZLUoyH5tH8YAjqjn/rj398MuJqnyiFld6AjZb5VFXa58DUqS
Dr//X8bf3wq4I6wvf17bYzAX/gZU7aXrxlNxbCTM9Uf4VIz97BpaBlTwg+9CThWpKESao0Ux3J9E
slv9pENtQ6WD15NktySbe8srPc/RVC7XMbfRScMJc56s+Y8NgP7VA4HmYlmNHkjsR80kn4hr1Eot
zfkZg36mP11k7lgJg7hcEZUmD836lS6LZqwPo5MP9Oe0px41oVaYEGueId5iJ5L2IFm06HnyppEH
Vw8VWQGTC3aIbAmCyNMbZmMGbQPx8b+q4tsdBy67YZ011MjBK+YGN0Uql2brbyJx7752I2KqADAU
3qjp71wGUOGamq/bZgt8zTacf4GUhVyl3MIGGwxCM6FPtAhSL/DMFwmpLk80c6MAnBjTyMKlRTzg
ZtB7925cZGx7Tl6maYE4mRUBkre2bMq7FXn0tMKUqEEaaFlj7fPpkC+bLJByRta+Txn+AzOYmmyl
vLYpsd6mO64CO524R27LtY6Z43g95/kc3329mgSe/uy/H+pA5+qQckDDxA4LCKrvBG5ZjlYsIVba
8XWYgz1rKPl+koSW6KV/aLM/obvw3KNdtMlbVOUxgIDQ69TGwZpDPk9hBiBwPwK3IWh0n1L+RAlZ
7ty946AKsULDNNpIHEQZ7D3LjVFdVxRx4j9kT1EbIKZPVjz/wjmk2Efi1df1D7z0miQe/FsR1g4o
u8uRw+nTZ37VeEcMXNpy7qO9zXTQpdFvaLr7ZMgM28TXMrmctlO4z4m17qgIBowU4//9w/VXnSKq
owglvkN/E9gUBDKVpQI0FQNZLuL58ZoZnHV6dDEGyJHFb7ul3gE7DpnlL8YuMKBuPZCVDaNgYFYq
IC03qE2Kk14Jnv26rpyTr3HXDpNL9IAbDCpMXLYDY2DPUAnWTmTINcmpxBMc0Jw1M6H8FHWFz/f+
DCgPbLH2xUQrUGDNUWv6mwJeZd+8aIpLC4ICeD8bAs6tCHCOWK2wojxV33+HPqzAmZRiVG6kFnsb
sWx/+PPEof84iinfhGBlKNBj8La82/ia24+vxV7cYn6jfZO11rQKhaOKhKZeJ0xw9m2R0htsO6Mg
1DaFbjHRI3KIvXMCPThhr8OYfqNdKIoyKEZXOgBx7goDuNNOt9C2odrRRS6iNdAG1VqxHUBlxbMs
NOL5himaLZqQZvb0vURyHlICIlyHFF3wGDlGdb20kYh9f+EZsPOTNrNAz8pINxG7hTsMncsEObGV
Y2Qh1wZmsv2ozIZAH4wKw+OOdQz8/MohcoVvJX0328Bq6LVrLdD32JHUR2h3rDBZRjx0/qpGvdue
nMG7tW52ks2QbaqK7rgDucv9VSDmQSOD7keW7cUlkVpNhOo1lOdbM3UVaLpuV8eATxlcaJ3SwFJb
v2ZV0TWpIAsYqAODCfls8aGB7Lsavx1l6qBZw5mf/Fedt2/y56j+6UPEWS0CDUKKkYjvDuk4OinG
ibMJMG9Ao+jumeOzCQC1gs1MM2JghkcZOcbgGR2DOSfbeOmtLkTN9k/30rPnwro/rxjpq9oQjddQ
onSUXvV53eEjyuiMEjs7J/CvtN4eZ4JAY2MZju4qAbU71gEe2AnSYIy3h1z7EU/3X5Dn6Vjkr7u/
i6RM+igLb1Y02LrRrPqbXkmxvEiAGu3vN5u2ny2yKhVY1GYIDJTHI3NLpihl/tFIWLyRTLuOyfQM
mGNAQNABEirF2sVjhtXDlz/EOB5Fb38rCBmaIDhr3DyIWzoqyNQIioePJMSsssV5U3oPmnmF2SdU
G14b3ILw1jNCIDqvZQvTSy6+RaK+u/qU/kAjjQN4xrc4B8MP+qq8sFpnTU9m4u14xlZyB8hjPeuB
eooEbnGk+DtySkZaDtJzInVBRhxxF2xAk15CYTnLjgNoFhv0ilFMBemirgSt9n8dQfbcuEa+HmZQ
7OWIO7CtEv/v6Z3j8Ke63faU4BYMaC/XJ/xyuBKrJgw/AbxlEvu9F8Rsic7b3DV3Y8EVw2MDykQ3
t3GCUhIc1aYB3gi6M9KDq/CeNjhu5baCRYhaDtxBjhZteOioYpFBK86JXK2cyQws362O8Vwiyz2X
wm+YVv3zTNeuPzNAyY1wt1d3tGEN6TJy0RKHhc4od6baWNZP4Gg4oboiiaCmNbnVvFuRCaSNMS+e
aAuqLlNscmxU8lNBnrEJQjLu1U0QOz8V0KK4PJ1MXbC2lg2/FGhjDj4Yy3ici+/rlbHUVudQ4J+X
xKM00RijxiGzZMhHpX6x8k+hAM3w7zKvjDpdJI95SJMWgyaHqAkPtA1PyltZUBNx0RDCSmsfBeQo
jDiYbmvjqH6xsi4ZBt0lRunaWapmPG/vg/RTJuj9iidmCjCY0dyfZFawUMIHziC2afUXUAIHan2J
k0X2m6u/lRLEd1ggCa/EF4gE5VAvIayCgu6xLdDNUHWH5yY3CGYk6NX1XyYuretJKRnu/c0UgbrN
hD9pFXIeZwdj/ZzTZirQHlUe+8d9mIOkSzVaoWb0yBxD0XX4t2gKzjCkL45r/3rcNdoTBeb6NzIq
fsTknqCDSG5aBOvSCbTEjhlNHj1wSMawCCS5lgDxU9ZlV8D2aH80AQyy6W0ovJ1zSEvu91kDnc5b
IYDBQhSCcqc5wc7uM5hkK5One3qfalYfdnW93vyApIJTzn2hEhRjQ5+YTzFF6djZfezaV7TKcGtm
IVMZ9W0Ls3n/gvarDuzLLIdHJDf8kSzpjpzGq+SAwhN4o70qiCkIVddgpw9n0gvxWBokU9EPMXzr
LqXbnwFxqKX0nT2NVeJ/h4Hu8eqcVrdD8ks9rVDdoWyaGsMe0X45sWJtYDHnh163z4IyKj5cUkD5
FGiLJHBzADPYTAzgw7aTUsqS5B9eo0QN/NaHq185fNyhuvBHLLDpRVpuCBDyaKIC+qKkVNlYyMC0
YysF/e/fZHJfMSglN+ztnxhuQ9ypl7p5qpjcoeqOH+vlGItIozV6jlozRFd8csRTMwRed/L+GcVC
IlTfMYlfMAQJnIhH0kiUaKa4gTajuo1DRXU4Jbzohbs3QqQ9ntirv5wK1e9PLHktJ3oe9bqO1o6a
bZmN2sjejfdnjC4goYVv0P9NRIaxT8COgzI39QVeyunZlTUmGVasrKhBs2BpH3Qe0msKdHxMocS/
SDpGtVD1Gkg6GxS1wQpcay51+LZza9orWusAN2zOh0sRxozhXF1bwz4jRQnRdy8y9Z/Auom3mUb9
FAcAgPs6JxiXTT76zycwaYlwKHXy6GPxS/rEgGbu9ethtZoFdoGXPSVy7rfZEBFkEuaYCDf3QdDj
FOye4d0mJ2+7ZU7quuC/fcaddFBvReF6NyGptHe+QEXJupi74IEB9bBStzAckzh6ppxhbmZMnE/+
ZlR6yfxSP/b5LXsLj84cfWrZkncIFLzDh8aROahLqPJFjIBGgesk6GpPlDF+Sk/EsngeFUKkex4N
zYBF0o4EPH+3upsux7rAxwQQNjUzuVo7l9dTiWIcXCnbRPmnMEhUb7xoUNV6ZHwPhTiIQXwOJpgW
tlLghka7Nje+bPKu47UpNKiLtVOX5fcfAuUXclkyBx52l6ecXv59QlcuboYjgNOImOsmvZ8VbHeY
T9rbz8PEfpdPSxyBblT3vsHLN64J6iJsgWDeOFkgSMjWhoYRWmrzZjFLhDeQTTF7X1Gbz0Nffj7U
MZnVcwXz2kLr7yLSWvxs53BzSSg+1cLEK3DO+mOnwqOR+tEFL7b0bYkZZtyIsIuyUrKzqPicI24w
wMVJuEw7cPN8RQ3QLGLerRso6HSs55XrP88CCHvU4oK6IFg0+SREuT4mqF7kcjzpJw+BiU7prkAI
0Di2CDo4TW8w+YZ1oxanyuiuAUb1/4nC7HyU1qH9JwM8x9AcCfCT0Yg9e4qF3CTmnawt1Akt6xUB
KzDIG+q/skpK+k9j4QfCMDOGvyyxPlFl0XuSCw3+I1VDh6I4E07XSq6KFuzS/leUozkyVm3U4rXH
q8PhvfZup5I3Q1/fU+kUivk1nxPwMOpKRF8y/W9w/h23LoFbFhqbvbrPeC872XDoZDBA45vj/ncw
8WviYfdGbFbCcdf5sVh5Pbu8bMOTAaqnF0rVFO1slAqPxMSb7UzXMcZ4utmRRJ8dD73dxlsGIPlx
Jdvs7q4J4tNQj+p1b6lY1oaCSKTDi5Im+lRMuZ8WDtHA69k8mxi1rmQ/3bYvJkdZsxKQGET5GoBq
PPj6r8u7DcfyUq0SoccZVJXAI3dR+XJB+xbpIqNgc2MFbRFNyfk+2eQDY81IDIfynjwjjIs7bXwc
K/8k4O3Ya33lE1GnjxyxrNhVj+FLb6p2czKrkFg+xZ9Vys2tOvfAumYg7XnowCGsoufJiogrFlWc
73pvDN+6Eh5Bm6bJzax9aCaX97/KlLrUHX8JaKRJdhJ9vJ14hz8bF4ji5XVoscdIu/WSYb3c6mDO
1Yifr7l0hakWoOhbHCJvWZkYv74I0dozxJN44AeRCUagsgjIN2r2OdgcajiMHgUcI5CpD5K9Nd+M
WQVCpAnVDsjMvuoQJ4K7iEcmMfe3b8Z6Y8pZk/LVXk6iVpIo+LwP9Q/D+eNeEFX3swKYcYOAe52e
iwYZwxByB3Lye9t5zQx09iwQArH4+2sUIvO+vDyZXzLxMSfUTu48hRO7TGBQXsWkIVwWKcWKVpxG
dgN6K19jCJq3+uC74lHpKaNIAdK88GiQYwXtmLBHq/ljDwTeX1CErSEOz2DxSEVFA1aQoANDaLqF
4zqJv+XAZS8aqifKmHpj1FJci5wuvuH0EalKrQNv1WzWmjkSl8X+VAa5vLZ0qsBfTLnIh/ZQJvJG
56k/tNvvTYdHxm9Sn6MWgfGL+/1fWWGqeZrIhZcOfYlrxE4UN4XWXH7aJ4a2xerxBfQWwXS9iavX
xSq4MQER2mTwc1wzz63VAfjwz+FvMf+SzmH0K42h4/babcbs0mBHBGgNxhtquOvIwHNpSLxtxlqu
t/vsjFNq5B1OyE5HCUGoKEr+J9thYKe3ALoXq0dYX7GpARIwS7SMPMxkE5OKfmHGlm3L112USJun
z2HLAH8zGxy1pdK26Ow2iNwL/gl39cy0UUYQ+c5xIijdZnFfAmPY4fOeENFPyNT6uSXu7wBaOlkP
fOqfzoaHb+XOmiFF+bcke8R54br0bjjkYkxcvAJD6eixa7gJEWygyzGT5mXoQQ77Tufw2PIQE4wa
qtD4JN93G0RFJW67EiS6ZiSqisji8k3peRmTDiqx9pK4TBgRSyNcs4xqWy/9cnDOZGAxbvluOfNF
gyO0pgh95vRGyln6Q32F6gHbO+/rvC0PyuNOL+uiDPZOQ/RtzJJFzdo0CjfTR1/FPVG9CFYETArA
e+SnZxCuXILLxeM8L9lQ/kzhv/JMvC0/4J2y/2vkcAOUafxXzi+ggqzhFrSW1xrpqOTqt6/VdPvs
X2IBw4k6VZY7+uoD5XwEyvMqPQ0Mjr7Y9Wgk3d3y78rLg6HCsmWZp3VczJd6Ii7XuY1/o3VRZrFI
roDsak/pskhn6pWcpRvKI2GXxWNstsyqwHdeUxHhJZ5oQ7AYh00JYv0g9Bh8ZMjVi0MNyse1YdTo
kl4Qb90Xv+oTqwx52TqplUY4j7+FAg6VqzbO6t/XxH0jIkcL4WJ6/6LWHsn+sOkqKFREKcuL3b9r
QbfX59uctH2zYHTN/YmedQEy9/a/gP61FL++E6VoCxByBLWwsWza1eTBwKIaS5ZyLyDM97z36qpv
6rQ+Sw+OGCmt96HqKc0hRiZw3xTsFsFWIzhE4zex/6CXinfBX8DIFwXqr2aitAPAEtIsxtc/u2WB
d6hVipLjn73JLX+5/cZoHyxckYxM+BOPjDfzTOIxPGeu/+8s/JHU0QLxlR5eTYdPHeHcAcIt/qq7
nkahSEbtbwHAN+0MS0yeLAqCSTWqiuEXs58wuYfq1EWdRs+5NRCfSvSskBpy4MvUpzSMSluf2SIZ
H9iWPYjTKZKWCTIAkVI8U/cnLenuiOJ0EZ9v1l+ri5aUUrhmffXPmWXI1HJOCHXQ60/mwKR/HHdA
zrofpZFwWsROfbKHSeXoZ+HmXBf3BiOAv8wF69vRgSS59MkSDDoDi6XGz+opYMVoIjezmEsG6Nka
efapzlZl36m7UkD47w0zqLUxZistg7PQY7MW48LOWW5sFR7uGRKYrHcSCnK5YNxVuDMKH7V57R3D
woVpT/z5Tm/ncpsUYlTJwMmI17IpxeAikM7/lj9GoG8MWfoGK82U+IKa2VCHbGMae8Xpm7irTIJn
t14KNEqLjmCIQclHyC7xCJaAkau/IuIIWbwHravICPzAMcOXwbsIXwCJO5kIDa4s316m0t1SxmtL
WO4IVkjAwkWHGcop75oxpeqRo1Vsg9pQGbpR6qcbIS3W3qmTZ+aCLSA1jqgxfVbh/69CABXylvE0
UpEvBlziDNvZHRtTNcfDNK38OuU1a4PpbySegsAqSoOiYDF1O7J4oyTkjHCiOGTbhi0WPcxJsgUH
j015GFUYfvXiaEczxtDcGmDmN3nRNJ1IQt2B+jVh1y9+T/bfeSo5eBJWmZrKunbP2ZswNjMd10ix
cs7xYP1kv59BmgKx9W3gf4T4gslVa7+GGrHYZpWXLGAsIAdbRfqP5Fh/ZoRVEfXjkBIwOY1nFZgt
mDtzZUxkH5KVO1PXkY2xoRtD/cvGAgXdo1S07u+Hyl7KDv4drcBmcYy1PxCzneI3XIXTaIm1gK9u
m4F7glQi/u4Jl6KM8vid2QXfY42m4WlBNg3YXSzeDxkYgh9QlPb8mBq9zkhmgkQycw5sF88/7r5Q
jhsIF3uGiqPirzCunes/bOOGFo2S7BVnMa2UGQ7afFEE5luqm7dTZAKIjHfTRI5c70K2yr4R7o3M
GlQoacBV+A1SdSTKY2s4Wn3k8VQZ6q2HKVkBIQOf6xfpvz9IdlCMkl6MUihhUZycNrXJDFlPrGYS
XJGbNa/nLJdSQBGWpRB3DZp0ynB03ApG7U+6+ShMCRHcdyvck/4dA9ZPn3P9Tziibqm13qHEW0/a
Fc8ff3jH9aN7tlMzsTNEFcHA7iF0UtUJ7ui8F1vDEHQKu8oOLUSNXRhlm0jw7vlq/pt8A9rCUz02
DiGTX4K+a4/F6e3b8d8k2O4XOM/sJRIbL06SWB6g5+0u1Y8bQGjV1netJ4PH8rrGKgShAUV/3TZk
xuW/mQRNZDUFR+5agYkCaXA/B0asBoIisKzdWUnrqoJ3brbPfkP3MxA54IwACRrSZbp+orBQ6Wpi
llHUti5u2YhPaqf7WVkE4QlM5Z6HQCFbBJ+rG+/xi6k4iHIk4S25cig1/Dnt+NUIlE7syo5a3O9J
+MOZCbC97c1TW8X0t5ObZ6iZW+YiNoglSTTfBuLo3jwKX/MRHd/HfNLUS3T6ejU1+29Mg6obdFo8
jskf2jhFhxakuuF0h6OMgzudy30et8BNfn6zLnGgHpmIMDauVyhT4rsb3O6Xtd4dNLMkP1Nppq/g
ecoKEEOhki9lpbLIuo2re+Ul0A5G9c7BXDNi+ZaQQWNTn98d+zJCe5kzfllm3bxI4eNKIXHrnVK9
TPlNqBYztZsZU+0dAnJlpU2AwX2sZvwbvw32N7KCx+L2JB08IGrHAnxoO2u/MhZzyYvCz3zruEuW
z96sQo7ha5P15XBQ9vBI9fnVukF6NWsDKtBgxOKkfLA+uwXycpQb/AWsKNlUZYJsW3XCasWjZ78F
+CMjEniFtuN6OxhfBD1veKz+G7r2tZ9Vj/JE0cL1WghHahCQdha/DJqSRJN/Rhc+ukpJUyDENm/x
1SYRVQUmh34Vc4N3rRFhMiMqjZMndFlMPuRkjvKjMhhVZ2gMqFjm4y5Z3uFtB+cZuwH+6TViq+zW
iRKH9xy0jIbJu8gxXKK6Gp6lBn2DIr5l+Vx4EwZyPTPEeQNw8Fp/js7btodaTfNmRQXmJl0ZOIbG
OckRsO1NzL1W+LeiKBOZxY1+VGKkfptHHgp1iHNDJQw4PfUnae+8tzBw+G//LUoeJp40E4IvVT7p
9T4eSA3tmkofv0N3PPMh5wfEwf6sc3rfYWoNv7VR+lDH1XEPT5iERyZcj2zHBdcypOkmcH4vgklr
f4tpAU8HsPI2+++k6Fz8bMEis8YHyMLg+ss8C96GKIS7yoDcdKa2cnqzTosOrwpr1Gq1IouNp64Q
8M6fm//BwXihTLnJNyGBo0dNt35i5Z8R2G/xqMyXDFziPLQUevk3CBn3QUhNJpVymiQwTBnMZwIg
uzUwcxSmk9XgVcy2ft63jWrUgZwyVkB086CjAsKRILr7ICMpftMrL9UQeeij1eaSxfytis0NBjpS
cBzpGAAYyEfILTaFyW4pySgkNQ6RMZtzD1jTaN9IRD5//qbIpj7V8AspC+QQ3bxua16j00NFx69Y
i611Kj8xLr3pjA7KYMNptV0yZE9zp/k4GDyIKdt0nH3yndY1e+bEB4UaxGHJB7vyzawVANveaK0V
GwjGscAGsHpL5nNVZ3TsiM84Ua6KEE6rHJ9xyfLS2Gbasuxtr1dhMo7ZHXNF5WE4po3UApuBjn9t
Jpp1GDLT9SpYFZlapGS1PxJDpMPswJT7uApRXmwxGeROjRN3z9dKVR4HGWARUKgODU/VuhAId2+X
jN+J5QRIdLbGK1qOwb/2mtmtF/MdEJEsd184Pl/anzMJuZ2WAcRuBaa8GQ7G4ANE0nPz+ooSJdVa
TN8cJfv7jbxlZeTlbY1r6QdAaDTwVAu5QKS7TVYRD49zV06rATd66lMZlenWSPylVbAHH5grBk0B
yxmcoOXpyJutDqfy1p43WbiFbGCBzity0S0LUWMWSZiDoL/bcc1D1FZ99PrGczCY9k1U4pGjGEeR
3sZrGBMl0XFA9BouPvdiUdy0xHnPR6pCi3gYguBTM347T+Pr8Y2xkcfjQPYyk01poZoQTmgHEMCb
miG2NvtqDXsww1j0p8CHI7L63dB+3uYj5MlecOVDOekK1GuPU22wbfvM8QcN5yAm9mXQl2UrDa6/
b7+XcLUFa5lnRe4hMJhDHr9qcBQEBxiKLTn2N79eshguoaINNoNpP/nygNfpEe3g8d99IfPH9oXY
HIsjfnx4gFvE9jJnSWKEy7gv7PO1mSTMMJBKonb9ITKn9KHLCUKPZOO4k/u/yiyahT8p2yCGyUe7
NhqVfJmgxHU+a1lh6gdXEgdCUhOiVhep7mQhGzaFFwFCTZgg082nscutSQnyApr+ydCcoMhXn2rz
keKsimQP+L/qEoE0AHFBejCnwSZTmCMRjDlPY9nwwXh/G1b86HoaHFuas4llD6ExdylqI3UHutSB
oJE72fjFBYwpg0f0CHA8Obl0cV6OK9soacwz6oZxzR3bHbS3pRhw8A063x3hqWuuebbCpptrwj53
UpEMx0mMQI7c3PX99ZWjzamyG0m6PRsfaGK5kg60fqRn8CFr6rmPJ6Ug9wgcyn2Q5kiOGsIoH0qs
fcl1WloWiytabEC/1oyTr9C7MNh5DQMF6tth9NvBeJnB4mhm+vt9HEJjFXt5zOvaNnvZOFSk1Ps0
zdRq2BXhzCCdEZ39O7Xz3yEKW6FDV3ceJld1OsZDehUoLUqSFXu9yytHD42GsgjX+UP7g6hMV4wU
71syHQor1lgjSDTVShPY7QhqGPDmrS1vgh5znbxsXfa3lnCv0z7YxKhjqSSyEblezLJHVoVang6j
iXwSYg6S3EOiE65MjHXuaP59oU+FzAbGOzewhy2FBrVSazHNYcTYbhJaWhSHoJOipUQ65E3dDwSy
VLXdknPuyv+75fo5q5XAJBnphSMOoHuPbbK70u2Wa65OSAizylMdRV1bwWIkKY2+gKC/Cc7Z8NAX
O+VZ3TxgAKKs6q4aPXEmMoA19MxSj2wlJMP4RCJ6EynVhwMLiYMU98DUb/c/Z4o5+vQfoa6S7fNc
FMPUQgLkkjT3qn+gurWQUaLP1yaZC/IjSRkTN90IZ7y3nwk2zOzmJlvMzSyuT4hOLTQLDQVCNNgo
JzaUWpYtSoNVx6fvjKivBy2DL4WnEHxccT5WP5JyzBLLy+SeyuIBFTbfgSb8Gk7P5BMj8cyAcflr
oIsF5viW5QdmQdduv4vDZXO0AvcBNb/AGi+ddCAmyi4UTlRdoJdytYUJ8LoRnNxz/dLq74u7j2xJ
2h9YDqEREOPFIzkaa3TBktvffe89W+Fx0oDfQdFXgRpHjXvOUz0vT+ELATX1r/txsgniZ1mppEbc
9kp40fNVRXTTUh6O+DlTJ0Bm+8Fs+qDGUf+NFblkX/dbn8VJJUPtEI9DLHHghofkXc4Xl+/uQeKm
Hf4F/5WEg0p4Dk4thrzpJ6B3zL8MvY6cef7gb2DCjIl68c7ic7BNk4klq6J8kGdG5cp8PathWe2V
3ejFtGNAuoz2snb9FMueY3XogqGcpT3S95z1NhRRa8suCFHBbcAI96OabLvg4ElNY+R7m2EUi2vk
xTk5Cy9HnIWDp/9iVVUZRqsLtXSH0YBdhUVXCexyYYO6ip0VscSnsKQsNPtWztYywW1+kKIsMC/J
upx9MtXapII/3GWRwyLhEuEHfJQgNK04KJ72O4FnAOJPp300x4QwcMwbjHSyRiaC4rXk6JDfosqW
B/M3+TknTs7PW/nEv/IxElDbn3H0iGmKTkRnWhTgAefHzwoy7edsHbG/XvjBVY3KOKjXJQowxqqe
7ySiJpptonI3FZIiFl/yZnQo/SSAGLQtRVOGuzOLtXXf1Swj98IGHqE8UwqoyY7pDMCZux+xGsVE
WZc3pJgWqX/ohmaGfsDCVY+KgOth5GD5WpttVYoKQrqS3KRA2B0QKYeE7ogGpnREYwwrjhQj13Ad
qCRcndt5C0LZU3tOG7+h4mxs3SpNIq6SHo6y3J5XaALjUxPFOwd89wMaXKmjxJZCKxNDMoaKSjrM
6YCOASye63FDYovheqTttx3sU4oHqTw3jBoiC4OhUFjpZkiuwI3VKK0FYjVf6PT4FI0uvASaGzPe
nX9aIXdC8N5XyG4a/wpi/jAfKhtGJh2pchmS7wEtTiQ8Fo6rww8YJRXjxM8y4PNsQZRM/fYB5OB5
iF//m7jqt/XpCSjo7X5XkZzVChkz/hFPm0apDUQ4iut9mzjBhGoMdy2aOtXpvwiFBQJXWIQAAJhX
UDd9Xb7O1xcmUBaTFaO9YJAtAm/E6UsYlV/yKgmkHa8lKfsJQt8MZHm3GdpAaC9/QEcJx0mOazEd
nIpISiAqWnjeABDZCvXJ5gGfG9jax5gMeeWx8pIhKWcnFVEmXNK0XpFit9gnrW5fosbb2YpJKRZH
gMKwbchtIKqAo0njxhXGg+GqRzXfXS7vzuUb5sALCC3zWH3gieUTY/jkzU60av7xQMmKPAHmjuKb
wH1x7YcIDfkad0ejfhKyy2jNKybMQp9XEM1dKFUWwei8AxYb1fwAP/M3P7t5T0VYxqBIKiT+TEIa
L+cbE1kpy0x55zfUlke8meLkNxuox/mpct10CdWccjByts3/qmH/J75LBsmnF0BIAgx8y+taI7qA
s3P7UpFLGMUI2QEyUbI/6JicbjKcb6/C9L9IcKlWPp5qjjwaBv42O/CDMQDr8kPRiLGS5Rloc06H
hBTZbmgA5vvOIh/x8EdRlFxJXLPropHV+H9F5Fmtxt/yKdZVpEHzGpyIsdW3WhQlzGwzha5SU7Zm
NZ0A5JkH4eJSykIsZ3cgqRyZMeDKY7zmVfpLuMs0v/6bhCZd66LpidNQzP1OuARpwPX5EmH5Wf6w
P/PgWszfg+GuazXL2NXfQ1FRyJ5RY2nXdxTRFEaJKCt7oEgtBLeGFdmNi6oAtBQU49hCsJtegXf2
bL1Ef+rv/id5aXBcHT+lSuIL3Nu42qo1OoYgy/DrtzFQcd0h0xF6oOKFQNvGeqS6unWVZtXx78c8
NAOeUHAnpDDG0G3Fu483HGNp5guJJbadgi/PUSn1izQxOfsPeTohnQpKwpTi5S9TwrbXG0lpdZI5
G39JmuG1Zbs8kCkt8HrIZWop5n8QuRYzzgrazMRinYTOGnd2Wx3+pX3lae1loAKxEpT1ZDlKfoQx
wWskNiHYtJ7O4Z7wcx9igJiOX3YRJAjFC2cD+YgYjnVAMpEeoyoLZVQi3f07mIFlwZpXoav0bvWr
++NS/Y/kHBsx6RI1+y64PsABV+HyjwdPcV0bCjgZZohDk/vzPEjrc7mbmn1JoZWZVAkVGMIPGDa5
VIA/W7RWTKAKOXO0REsHOWjTMI3KIzyEVvOIsgPehFnwr8I+GxfmLQAkY7VP19w/tZ5RD37pe8T/
LRr5uKTQeuydlGxMo+tBsEsgXiGgRJ1FotPXMqA/4zii1u3FemQK0my/lsqcj9BrViFyCQv+D3rj
Q4LOJaYeRQlBbfRska6xu9xInBYzWLBSKfaw2BIMrD8Q8JAbd+d0VI4bYNJuXM3rq0a441183bDD
ufxhuNGlzkbZ2SaqRGDXKwhPjU14Y/kgHEzv6+Z4z/rfEWo9um0w8hjCdnx82LBhu3bUMm5Xitfk
qihr9jK7n36jyiGP+zZ+JhK6z4IgeGuNsixUHnnFBeFszNbA89VJDfnMjOqtVO6oTCvJZmkoMiQD
tmE1HXNBNhw5vbhP4Pe5FuDXBaXhSSHcJamo1h9kO+sGLO5CpthHtuSQXRQCtVNW65kJiStPuStF
ZHYuvwlcAmCNUAeFpdj7mg339x+GQBfydEZyvF2qcnopD3QCHLTX0/L3ZfNDi8Gsg7Zq5xnncGWN
Ymo/lEdeTOk038sAad/xFasOY3BDB5FK2WGKP96o6EmA3F0u9uPZfpd/BADzFszQ6ntd5O47xGPT
GmwuwrspHVJKR85p7aTqxOjHGLxVCuGX5BYiHoegfjAG6UpIdA/XsP7FzJ2O+o87dt30IJuwapvc
k1Fn0VcClrqVc9AUE7Neys/B+WvtVeLRxoodJDtOIHX2qOhPAE86f3FkZ5K57WLdLddoXxpb8uIu
F/RXa4yIkVs2oZE0P677gSxU8xYTv4duX1pfgkwcqVifgGoeJVZxTpZrrNx0SO0Tsemj1hDrxXOL
8PdZu6SAVBQWkjJh+3zNz0YCwTFrFNagIg4XlfMDQHs5gKPimmJ98TXQ6cFnYA/9cEPdkOVCPg39
KAG5GH1dZKBcyCb48fEV7k54qVmhxi+auVHdMcdHkZUJiceENuiqAt+pfO55BOQXXIDbB8BqujUr
NRBlq9I7z/KjX1DX5jXO/AJ3waTe3HfR90//oxFpm1GQJRouSoOvTEldcUnYKc7ai0IySWu6dGqG
4/KYHtSqhdHuwQJJnPCZwtc0cwCtot0qLOlKURz2l4LgN5/Rp0dWut93jREqZi1Txk6JILGMsTO4
6IooRUdKn20NmSc1xmgRYgkzjkYXbdL8/ZpwT5JyIrqhnFEb2otMakNtHlDW3Mc7DtZAugSre3Fh
rZctMHpiCXEHy7JhXth8BP5zqdnyUK9rUCh6pq1CRnHXiETw3FHDQZn+Qa8tcLCfFnTNc9e1zUu5
tSaEPo1xOdtjdE0oCgKDakYaEhpzZbwgLpuZOltEar40Nv7ESMLYS1IRE0HwDm0WOKyl6XHvN9aD
xSF4obfnkciq+AyeQcCqhEGc8Nkn3JXH4Ia/jOaS1jvxELdlx2nW48+2VxiBtQOrZ279nMF02Qi5
9vDVAXVXSnvL3qobaLWfb4Oshi6XPdReZoX3dxKyHP8uvl3pQtqCPh6+oDThujKd+KewW+7/5SfL
TNfIb7ZdtHVn7IISbFOeBT8QkMcNlD5iPCMVs0kmUW11eY08I5U7b4dKOrHzqaXeoLE8ZArjRGfM
bbMvosiQGGWY0errVXMBiNFDrMSTcQN/wwjv0S/JoCCt8V+Rebh/Llk2YhoRzEmW56JEt1ezmD0d
quEIFaM/OeLX99QIhJ9xHn211sFrD+oxzgb2ghNir/admn1/Bp8xeUoaVFeLQ1oipwFQpOTGYyUu
rhEaWhI+quqUxTZ42Cb/xNKTHX4dTom/jcKLlemMBg5OBSdw21092A98sZeAkD3Nj8ZQ0bGAieGP
2C/KxqBeQcNUGkpDkKP6imfwnRpjZkarKoWq8DmwKR7imxdA/E0SMDsIQ1/eFE0kL06wq68PpqNU
d/Po5kQhCJ9NGVEDLKpZVT6GFvadbCqmzyy3zDIlzaY8299/TtACWEMwnzQXI7+G172VqhJ6hyFA
N094W5XBWxo8e0lldSBBRm2bowEfL0yjNQ4br7lTz/DJdWtYl/HfZOZ7PcuKrpANm9zapRnGOWVU
Pd8TlLkChYZh4qvC2xs8R+1zkC55mlI7RGuD0FBfA9WNqsin6TzKA8pylT8F6vqc77rTA4uDflvC
o13SaTCcN1A9UpR36NDmteK13AifVxDk+gLZeQYfVyQYaleoc7I5/t9HaNb2N9ZdyVrRCKfhERDr
ej5T2ggH2kRW8rL0oqlGLUoYLraTL69giV3EWRbvPoXQ+fppk/rnnijrGZQgOzGayULXuRoz8H81
C62SnQbD8DWdRgL5KT79aRmIqvRlAqOJaA4XCQ745WIlfOQHjSDoUPWXKMC49RjZOSjhgs1kolfb
5MzercbO5Om7UXbwh4giXipfYoVDNXEX6Euzcogrja5qKAqiFdrTpRUxoGNdYtjkuLDSLP6sHp9i
toI2FZkd3XOGkSbRnZI2+VXNZaQEASNVIfr+XRifVA4PZO/iihTUSQ+rS7YplQosIOC2d6HCp+kK
BS2H3pbEWDsfWLXlORS5YSQ6alv/Wv8nIY09r+ZZZa7bE/geDQIGGATh4iYE2lC3gPlxA//o/slE
MmdRVTJkdlOUrYLyn0Xwv4VVDhk3WxPB/jSJzS/6z03SLBKyKLf+Id5UZkaHY5v5tfeMPA2KdF5s
o21sl2vGTD5Mfy7GU7DsRqo0rRw8ENMSW0fULErVJ/MckZejXJXkUg5IwLhRmrywPcoPXtclKwnL
opQWZGXaARcqCzguUcwjFJkgDlG5S1FdKhuicIGIXeeGeR2WROHQTNp//6zHgvZGEP3tTnYqmDXX
knebrS404Zg5bVsKZ0Wu0rbG/UUcRZK0lpoPm7ugl6ZYhHj+dgup5HirHbHCXIiaKVRVbgJ7FLE+
OxmcWjKFbLe8HujV83Sy6RnFx6fTKHYIxdU7Ej1f28zTdRjftF7q2jBp6uGI9vAs0sR5e084fac6
1KNBPKJTUkyRi/J+7pqBdIWX3p+i/7zP4XqAUigFBqVS8GJWkH9AScAOgQELahbpPv7WFvz+OEJR
VNQMtGpJ60OS2KbZSHrIK+S3PMQ1OnmMaYV3Xbzpwp4xzF4L0jcsGdC0JhkbohwMa8WpOzRQ64Cb
Xf8AasbUy8G8C8s5tGfD7oxk/qRI1iUUlehjnI9efBj7ciJWHmk4ldqphfwrybR1/bwK7txH8sYm
vYyg36zrzi1Wj25ZVlq5uAZERB3bZ4sdo7EfwYYJRGfZpqbR0rl7nZDYGWzUkh361kw90yU63XSt
agV7A7H0XgvXGP6JFdjvHdTkeGRX3MXMxI7KBFPdaj8qDi50K94z2tnRg6MeyKrXFG+w3n0tXLsN
rMaZmKi/Skb/TuTJrI54a9nh1WMhFei9cNAfGhiG2McY/s23Sy6lhHhyblZm7+VEFRt9Fveesw7R
U7MCOs8M+sjlH+f26LfRFiX0VhDgH1HWayOJx6ADPfNHmQe/PsNddcLNh8CF8beFjy14osiV/wWU
Yd4IoybSH2LzisVl7lz7TjslGTdZJY06geQ8vdbLNCq8i6CNBM+da+nPnWo5zeBn0xeaJ6TwHmFM
SCHluVP0fB4Ubdo/9ntNCR2i7+rZJYmyZVnxg0pKDoodiBPvksnu85V6k5xWiIy6hrGG5UXOWRpg
q/3qNQpAGI8obV1awKK+Rbeom5y8qYqOyjh6QVanw0WXdA8beoUoXEXzsBR0qDgtebZ1d73Wm4Co
tugApOWNOFOc0PEKviPzSfLeO7em8L7Le8eWKYVMmJv0RikQQVkjqJUrfSB/nA0h9cBxh3Qsurdo
oO8SlX5T8slaQHdvyB3axpp5te4Qe8P2aFewSNrDuX8dbi0IdCJKris6vL+pSdtXU1uyUe1m2aof
9nQZfOCRJSQ54FY5fYDO3RHcbctyAnDOBv2dLN1Aa9AEy0XaHZN3CddgHAb1qOpX47jMqQGn0oQT
KbRbeYB9gGCuvLWpPytJR+hQkl7SB4zyTDvQ3f3Ot0GHgouHlpbGQhpLWEYh9FSzZvjAJ+i1C6QQ
q2T0hninwo9MXQ9CgB8G2kr03q3VPqsWYMHwm42bkZKQJQN8rZVLaoZPFE0UYNkVHoUg3RJNJDRb
t9JGHi2hmyyOgxsQhjI6n7cN+dltLYtty2PvQ9wWo5cQjABuB+O0FPWwKDBGcgKNjLbALCi5mnLe
PHGzf1cveg/GGDwTuGBP04HfuIDYL/Px7HTWLWuNSaPPXtZIMpgD3nlJGDrXsebEH9ILZpSXbiPu
nrx29XpTR9Yjd3Z8DzTEdIYZq/kt0JpTZqKBbtPDkgTp62anClHZC0l5KHiQwnGGfy+BrHmEpoP2
p706x+kCb9gfWmgWSH7xAP+i5zY2fKr0gEWs7COLyKrYD5pR/hW/cl5PaSQwPa5KccIrm6m9llgn
OwshVUkc80NVdFfOhxHJlTXRUqkEq8Za8PbDws/PKr2XZlE3P/9yxZPIWxL3/DkQnR/pIjvxXrOp
SPWY2F4uaFBILDdrKwY6+jk0R3WHKHxRAdcTGRz2DeNi/vRKQFEZJuifS4gzfFVfK4cGO14XeydO
QQ7x+xJOuAFxYEBoiSMcYIpMRSffFp5dcS+AgZPhOKUmgeBO43uYViEKnhuXWlu6WwQh2GtrcB+g
yJTonv9/LqbJUBr45V3bfwVKEuVr1LixYzYUAyS5TcIst4L0IJ4NPyVPWI924gqKix/NYxKGu+6m
plnfhBTItoy/m9LjOh2xoOiMD2HoQx99BvHYrpZ91XzlaTd7v/LvJDtFMrHXqJosW6FLlRg9msCM
6UkD1oLozRD9LGvOpsU1JcHcrqnsIEtOk5x5OSJ4mOro7blwU+SvViDl2FgiuZwuIuXH4MSqm/yb
GgVHxZKbA2d80w0O4DaKmYohFrPV5pZR4yF1gBb8phKPZGN0HpvzlwLX6Fxq5RJ3SMb9C7GRJsSQ
Dwu3gc6UGLH9z1KwmeZy1AK/Kw8MnOiZD93I/dqjcJop5vpmnLNYWVs9YtVnZnRgQr2LfyF1sBLz
FkLOGNoBhXjdYaSyhly+oD6zSP4JSYs1AGr9YTqpyNq5PLv6XWry4bZBxaa3F5WR+EC3D4oy+Pf5
w2grAeS3dCVsB8oF92r4aqKF5/KRfygtE1nTyLAObCRXB6EeCqwTze2SuHbxqSGnOsF4ATcHD6sP
+13FdvwdsaLMi8YSXqzd+QSBzFMLWamyAVZ2/GQklJk/klis9nJXKm4N+a1DaYrRLsC1LHo6gEjk
zBIaekVMHGMMLuohIZJaS0JpfwmJamdhsPFMUX9T+6eKNf/1LdnznYHYnxkuVcB1U4PEOR724lOs
DAAOLESriJixy9yHjITR4W+YfJQUt4QW+MwsCg/DRTeU5DhYyePFVT5YFQnbX8Yzb81COnfJ+EZF
wcwPsw/WYowmacaW4AvNEUGoRRTZn5nx57bYj7iRoaTjDtlScbd8snM80mXVF68w/qgXMYysJTGj
dAmwkEp+gmuFcJozpPN5xI3TNwoDbrLQkjapo2BhuiAYo5TF/SvXd1VWS124Fo7lqpR1sY+y+PFp
k4gPVZaGxbmEUbv598I9x7QEuIH3PJvWsO4BPiZMJ5x3mxuM0r11wbXzlh3jhEMWe+ZgN2cwuIBi
1vVrO7m+JgxgXWzczZ036IkFmeUsYRXHwyraQmWBrCi9RKjXrPlaMJxyjxlgar+k8zEP5TnXajua
Cm1WIuO128Mzl2ZYByWAv3Rl0pFx9O1sb+1WEhKz/ENvlfBWwAgpxlC4x6kSKPQpmOWnVhJNzNpU
xD1GxCFujX03Q4ckkjwGtxXFGn1c1CnjlDhygaI/JE59zjCJ6KCicZYFfDZVLO6rZI1zhf6lks1c
+e6xKBhyk0d/O89g/3MlNhQIyjzMA3xa63KXGrDrQmQKzfF724kkFq5OzfAcIVGoB8Xa51F1edHV
GOkys6hg3QPew5XyLIu38RMS4YhHZ45lN4u0kcuKSXViaiEJMVB4EB05FeyVn7hN/Jr6n+i2Yok9
2ul+QDSn+tt3FBIh/GT8BcvW2lEMhuUx3GcJjQcv0f1dUwIsHeT+5u+evr4umYmds23q/k3srpjl
ZsmuxldwZpp4Ub3CzG/2AIWcsxYBBQDDZXRipRBXjAmu7UxcCYJ1k2s0j4ImMwoCqYPC0knUFllI
2favr93fEDTrudHT5c2zSi0KD5QZvjXGlynjeXcEJsJtFCU7huHNe6r5R+IROyh/9eh+2GGnwKVt
Pd+IgD621ZIJc+ni1N270qOlD5KSVhwWnZnU8qoncnJYmthqTGMM+iAXOAn3cSbM0n2PULEzvWkf
BtA55NkgMBVf2DC0Qt2ioBNnVzYt3XYLcMPPg4WOlSp5JAjg6dvKdUD1cKp/bHDeTq8jEDRMX8H/
/Mh1THlBU5EZUq3y/OucKrID+TkCqdzN+378kIs0fn0ba59cJNJwCKGstUUbVYpbJBe/xW66hvYT
3YauYT5ykIiYKqMC22u659PeBZUyaixOVvHVYBSsDhmQKDHLWQEdNTYA+z37Q3WVcT70OLaymbIE
nxk9Jtd9JTs5tuGKRPVroEZsbRSGlrGUzXIOmbi/B0ClCekFJ4bg8fGDgpTYEqwoc0I4XT8flaed
ya7oljTGvGSV0jdGUJavi8e4gCr6ZQ/l7qzUsZJZ+MJiZpXifhfE2nOZCMudB2SnVjSg8mSx1d04
E+I6z1qr1a2hpHcZ6yB11bTW6f5feDT14evtT7acm81v8Ft5Gnu4XFeVFWzlm4pE61+3iIpMf+m7
q4jvsujXGyvvvrXcyu/PCZhe+RQw2WMUfVL6eGD8bxaKL4+nmH6ubg7BSARusGzPCjID1Hb9lr2T
1L7Y1DS3E8mgQ0dCrP6yywvSt+a2QUGExzviIS0sDs56bFctinUjUV3I3dQeCEvQRKHGiolbmUlZ
zpu3BpOPItaaKq80jhN89bRjCpvrmZGhcfMt2uK6ysYtOH4X/M3g2FPsJ9TH2O+plVgPm1FvY3NZ
D/vCevhBekz176fpRclwk3tYttRMHEqDTntJQsrt+Wax61TisNYWAT919RcV5GlupouwE3BgIalL
Yl4YwKUIWcr+ly22lxYgmxQ9Ruk0obKqCaqHlAV88X3bXcWECPEYtgeiHlFOqAo7e7LQwkx8KjDl
C0iC23mVJN5TGe5q/9tATQbiYvsIoTSn6qdlcCEG+3LZ6H+NVTXycPN/XzDfxhkp2QQM6fZ8yEBo
aTGNlyysZ/yyM0PXUyJIAbSUovEoKKn2CbM7df9fdMPrMrKm1bVeFDzmKpPEY+p+5WSVclJSTSyy
V7woRT/YveF7MzQ8xnWHp23ZutrdOg3wXV3LCSv5N4LGRWuGGuV9cqC50DlV/UEzKWKMqG2/6iYJ
ojVMLhlfpYhNF4PfluMHSmQ+e5mW3Fl/CchAwJXISLGuI+Hln3ojDKId0MCzgsr/+ulSan4WU5Gn
fZ6NSFhc0CbQTZ5nFMPj8xOehGcYM412udP4QEv+n3HJXxJsgUyWXLuL0J1wm/2KjuTTt+k040RN
UeayUgyNFl8D4gzd3jEKrfWbcVfJbONi4uRbpB+o4g1hrpyI0joK1N0Ib6sIIF0FqQK9YxYko1nK
NYs22Hx/eVjbAoeQGHrM//tErsy+iQfcqophNBSYXtlbw8rI+eX9fbMwm9ovWtR43ikX77ROX5w8
YCmYXMeJFnkFnIrlfNIVxpGrRmqcsvCpjy5AKfOO0xXNAhj7iNYqVfGRs4m3qOOFvfI4hHxoRdih
ZbUFCcfVRcojGWAgW9wCbjBoVlggUJuqRi2ahKcT/sXqMfJTmZ9x9IZb0Oi1W5+PDZBwwk/e8++6
1yVDrCU2m7l8FD/VE7Ei7c/oydejXMXzdpXJVy1UZK0JBIzSg2LyVchGDuO71FnW28/IBiJBE3FK
SSfiP44HSQKDCWtXSnkOeFSOok/1ABjOpNzHBSLBkWWJ082BWmjOrRfoEuYIjaDWYY3TZcRWDZco
xC8hHQj+C1fFiJtHmdj2AYf1QrFUfzwQZ9ToOEXjdMVvAu72VSNIJwyGErHU3biJhX4vN6l6wNPk
WEnAnZ5mK2zqOeP0DSWiHepst3mYXYDOFdUuqACg2lfriIxi8lh1TYftouybCRjCE3AKvB7UZwDU
fJFDblkDSLDGCDCfxsnrH0YyqJlaOT3xL2efhP9BNF8IJ6qwjiQzrssAybi8l+cJhyLxQJUxPudR
m4kS2nHb7+MFfHjN780Zo5LdcY3THLvP/anmuTwAuvi7nRPob0Sr2o+t86SByPwUt8CzC/EliJya
Pd2q9HpxTVzSbr3Eqga3G518me0rBCVJv1UFXfqKEpogwm/Ew+c1NwWC9EVyC+Sm3KDtb+9el0yA
RroCcZ2QFswGtphcFc2rDmjcOPRKrfetzWTcJoaakNLTR5RWaRAKAM+hY2P0a8Ckp4H8s5pVh5Pp
qZ9Sz0ku9A3iUcIq3DOKeYMQwJbUbUzIS6Sb8c68XzMTUNPOfVb4jYTXXh9pEC677od5Fd7lzdjQ
Hzh41UxDO6I9VZ2vOdaAZ3GT5q5mgqleUlY1pm295xNVzKTeFS5p6lA7BemlUC6/DPuCM18wxH81
GuFnPFeJ+QQb09pV/bE/Hv+16yPptwYBffOJUutF05Ugs0aeiAWmiH9LVGZA2Q/9KrAhZpuD23lV
g/lPX1WZVbhv8Kk9e3SUrHzjs+YyEraiAisMsVROLNM4iFOe8hfalP8TDwQjP+XDOdXGw4nvC/3i
Du6hl44YrjQyw3fpfU+85fh9tFmpfOSVMwuc9a7partngcAj0u97uN+fQo5CQkJw/B0+WJCTPM3D
jTLON0+CZEFRtNx8f95jmk3g1q4kIY5ZXcEwVGxd/ypxWvBSmnW/NrRF6og72mD4WmrafCdlMfJ0
Eq0Bs4K6F+PkB10Lua8p55p7Qy270S+eWlp3Bztt9KLuTLtEi5KgaXB2MHQZVuF9QLxp72udiYYj
dN2M04HOBpNb0biNqXoM+RGJ34hfly04YqEn92AqE6vSQImySQ7YLiMs02tYi8xf75Khnt69QPoG
x9YfUN+PPMFBJKhLFx4Kxv42pb9BNMhJu2AbX5Nds0QOmlupS9Vuvv9g2BTl32J9OnJFvVB3zgy/
/lQW8lojwcnyMnxkubADjcXvgdXcJtp6zDEraU414YHS0wliDg9dHQ+2v7k/snIBRp5RNMIZy7tv
xaVLuk9Jte+yYry8Pi37akgJa95xYIfpOhbFnOetPH7CKe1tpE00eZXBWA+QFjlpYuQQ/4dqTFk2
RCP8zVx5btASBEjMXqi9efMayTen9dhD5YhnD9la5wPh98yR8DesIbud5k1kxvFx5gC2YLlxVHPk
3+m4mscMBVuqfyHBywrsdw+8F+kkq5eGbCTla68sxmfISnrNadSqXR/nuWQu7VkeFTeTOnWPJQAq
ORxr0DkRSE+E5BJPWu8hM1anULtNw54SDnrZVmqgSQfYBto7uod8xHegXO5OlGrTBmHjDRCXMd2q
+Hjdhzd0lUBYtPgfhe1mpp3wXhexLilQXZLSkzb/LVSnWvPopr1P7hp1dGP8tA1bohFl6cC3a2f+
Rm7ne9kNJx5l5FhZW/yC+ABQV7BEcxu25rpkLaesbq6hqyN/M9Adw8P4yK79HpPAIlI9xoFPWGGQ
mFo0E5vBnhFxew2+MMKmeEcxg4CAVdsJ+oqoyEC9jltGg6H0MDFDgY6AuwlKqPl29rFAvpG0H189
uSUBm9g5hvwiFhTesxcKou1xHPwm6E3g/b0YNWCT2CIVVoNKjwJArEsGwVB4B1IbqUFaTRUXsV3V
lnX9cJfGXnZBQXo1YsUsdmkXgNMdj/Mqjt4kjFP8BRmp2hndZ8emZy2y1ftRLgVkw+4l1IW9PQKf
k4tz28pvLwhsi1G/hAQnzn8xq57RxQe9cGaSZlPsYIPrpPs4h8UhuQRRBOPYMppPuqbqoKKXgGYa
rOUk/scmKm57ulV7C9wdCqRvMBNm96FPNO0sHbcOBUijIcir2OV8t7jRV+BjHy5WahznWrAN4D5s
Da2xvno9qC73X6Y8K6CfC5lWSTYT11NL60EgAUeHX7U47AaLnbhWh9U0ucizq3oFDBrQ0GJL6M9W
bUvfoNuxJkn5ICehjqK0MVUpiDDte63V8FNKoVUhXwrqgo4Qd3sZt/ozreUd8rN+TPxwfg3wN+YV
f+IOXHd70eF2gISrWwE7JXaHSnkShzm4ILzf24PJfA4Y01JfMa9aP31dkMnL5xHNu9G0KAxQpxXq
eP5yG/KKsBH6VQNcsU6G5TuqgoUhbvUvFlo1DmrzS1qYZ3Qgcy+2MpIfdYqDhErE9rqHRNSFw09C
23QA7nHIykOh65n5my+fNo9jwExYtoccuSM4e7fIaVcmh2B18supIksGGAeXNiOl9jrLH/RpOwWm
rEZ2E/zYrRaKMDXiw9s5Ocou8I+B4pNCLlFaeXKkNSpbRxCLQZ/3LrBfy1xnZyp6+BJE8b+IvC1z
9SD4O6vtR2k+MGMhsXhCvHKyPu7lVJzxAP8dnZBkDLYUJ4mss2nPEy44/RKxaRwNceAlRDiv6OJ9
ZOt0O8QS6NGfxI2NktkShTWXTE7T3vCPTWn9bTJhSjU1ejxOZwvQj4V2Fo5y3v2d0oa44jO+TOB4
oxht2wD8E7e9Fi6oDIC1nYKuYu/YZOakx243ZNL2G9AnVAp7LnLQ6wmE0doanP7EGtr2DLduR9qc
k914XEbg5R7eivAzRNbrlqCNvFLu8Y1WrNM5tt67xtg1sGKkEvq2R74KpzyXNmlfndhVquUM0VA6
RNBH7j+uJGsyFKEVwBs4mEtUVl4VQ+eD+af7dx6/bqFQN1AqekI1jTFNPilcJFhgROCU5FS/5IL1
xxhDMC3r7Sf0u4SRcbJZN+pwaiJb+Mi+4aruvjmutv4Al3n7r7C1UBRinyQ+RGI9aePI1REX1YVr
W7Rwq09FDioHLob5rLOeAf2Rtbul5Rn+4wlMr2BvNxOrIfkkfK62YVVs9tPRPt0cLOgCQwokGmNL
L4cc6KEcnEY0Hep47P/fjfXJdHJAKKF/oVP3ZBFeWvGNkL2xzflDaZ2F+fY6xVEC3g+einGuVWGk
mv6JtrmxNJ0Y7uqhKVEEY+Qmn3z5qnobDHwtQB3Zl7ioe7Y2GVVUgA1ar42KXFLHIYxLciOYByrB
6+FqIXgvpLN+cbPkcJohwq5zZipFjkq1W7WIf2hOAtz9a9lZuFlxdY5RkxTT6wwBBL+SNhKsAioi
drm0bISgE3JTP32aNqs7e/9lOKGltWh215lOjKJSxqL6iYfQKICazXVtdtdY5LR3qETYHHgy2g4C
xZj4zeBSoNj5lMbroxHRo/SiErGjWJUpXaM9iPNXDGAmAdZhuOrGQ0B3mi+GkeMWTMwl0Y1CYzpG
m/ZH12nuJJTGQHt6hc+1OrT1u6kHQZxp17NLblSpof1uLuPobksvo5IJT+vcfoXNhqOtIJ45wq6F
ZtRXI78x1GA4t9p1e12QrBO0SWo54EjGpkeXJX4rRHQsWma2ZbsNh//DH6ndpp8rD3d5b3lRKrHp
adHbJzNqgYEBoYk36eEEC9OJO/FP+pBP9S83UJszAYtbLqdYNPsq0orbzD37IH1PeVKwZk3FF1+o
0u0OHiMDALrdtrtKKAXbcM9obZGpiWLPKbeI6GuvFah4b9p6jIJ3FUZgFMowGuA8Fs+hNqFTgLdn
R/Z0pZLUjLjKF+uT8dytYFOHqOwiAOkSre+4iWJZNWIiY7+p+JqPU42fo5mJOhxGU/yKikVU2z+v
z1KbHd7WSX+k87OA5TVodYI8ly1ZJ2RylLB0Ym9gQTN7UMkj4KHiPi0MqOQGL1X1XzravIy4VzNN
w6rZITXTEENkf36hL10jPLIKIV+MdawEqa3gUT7bRnja5Ndxt4OtPlU1nJizWF2kk8uYicxA6Vn/
SdziVnW97yR0N2vBw9yPLNfsg5hTdwdUwqEt5CNbwpPlxayf5GYwU/iXRYU0NqpDG7/PxdYYcRlZ
BYxdaGi3FEOD0l/QTnvFLcLOvOKhdz05p41wD5Xq1KFeFXJZZTdmebUSqWCJxuSKFX+eq0Bzwh9w
N6XtLUA6UBHnU7ZfIOeS4DH2xOJbSbY5qNZOtySYCUVCMtkLlOo4O8h8qw4lHTlGmLtXVGSkmhc2
u/9gLwcLvBt6z4Uxgww/omNG7oDeKT8HZfXoyK2m1xpPwHKPWPA3MAon2Z4nfZfAGaoOmo0GkySJ
H6wWO8wfSmuG2ThnZYlaqw5kFX2Or7192D1d/mh5vmJBbtoPA+JuITLkat8DyaSwimHFwC8iPfYD
Cgy7uJe14zFkd2j3xOqzKmXQMV3W+pOtlwX03fc3nIgllmSWR9YBycgOnhku7P9CtMilrPGMfmv0
eakcLZ33EWp84zma5LYT91fQnOY4AGar3LybjgBzsecM7Fl0l27kQAL9mFE7uJaKeJmRLSIU/T1s
86J54kx8xBBftVFud/+7hs4++LG7NRDXQgnDMXS7GeeoPxjnZdSHVrtYCTYdNBfImQM7JC574Fik
8CKBNpxph4Lp9ewcd+BbERHIaJ1d7npNCtfCaeQt18bGTJpj9jIw0MIr+eY4RT5BhRcg7O3xfVoX
1zCPMlcK8yugRbcqzYb0Xdn22LdFOizcQ1GaCFOou9i40/aUPsLFymk82SjRuFoMswMqKxk2ePQj
7eEtPf2Ndsetb7vanrCzdkZ7Ogeuph82aGmz0xGE9+wRpwh7ZY5eNM9+8mnn4cSUfAxoTXeygCuD
Kt3POtc5MKJpS7Pcs/O5CrS4/iUtjhXjhX0O3eg1VmXygXJUW8Ml5TMMmY6TvHJv1wQQhd/294Z8
CUOGNvRwQTmeHdDCQsRfOV80awqmt+rqW6kYhsFMwfs7b+uovlyG/j81nzwixPrQQVVwEpisD+OQ
xG/f9SvpdQXHaJnemISSIhCm2bWOWl6Nx+CEr339oheyXY/pjSGvf5jmaDNDcifqQ6qdn4QXDDBj
+oyMOenoIBXknd4L0crlzInp3+0tUOUSq9TEEElfzC14CUUKmeh67cUlCZdkicFh4DHXy3ZuSLrN
/bADeP30m79bIpKKJgOxJEJlCDrk2fM67qYNfierJu2HAZFkYr/u1Ar8BsQ3FJ1wHo6hurwmRNA/
wVJD3KVOtvSe0KshJhNlt91WQ4A9lqcB+svzoABOMZQT0cjOAq8s9EOHw69ZEHEutejg0zbuoinE
YeL96bh/trYgaUVK10nLc5FnRFJvCkamp0b+7huAGVIk/Jx3QdQ8LE0pSA4bzoEaeOh/L2sPfgJi
Lr5U0NdnBcV+FWNTgTYTGDY5zQMa3Jad4VFtB3Hvt8XLgFwwnjAeiF77HeALmPaJGoDtGZW5ynFs
YRf6HSN4B5rudfD6W88NiBZ7Lo8Yh+j/iaB90+PJdVyfcBaQj5Cdf6vJzVyO+w9dLNsMyeSyROF1
DXJtn5rHXOA4eqYYZaYVndUFeVIAkd0OQtH6k2dr/2r/QjnloZuW75KuW5F8xqPNfVf5wuvuuorv
SujiSW/kjX/xzLlZEdk058z50jTgR3XglHnqyxwQXzkpOprDDVS+6rRaGI6Ks4tXjx9VtG7cSBmI
4/Otdm4MR96LCcvQXJRZz4OeDwfuYJ0o9aKPG1gCh+tiSTW6OLQihbmkrR+WcKu/JQ45L2N58hrj
Geq5A+PwCifxi2FrslJMBiLYW6RjpZ/9QTfNDevYbNjdi8zmsmHupEEhf+QhTYO3VY11rghzF4hj
QO+UjTNHlMdbr1B4OL6XHW4qTz/f20BzzShKdk/Uh8Y7BxshaFXXLIaZlhv4B6471wyKFjWL1pwu
yO1FlmUvhWbSOR8r++7qfk+vwAano5lwzbpm+r7eMPk6+jsLzi9cGzQBDBbqpqOsFV/upc2cb1Ms
TDr7vt/mCKmFTySUaPXSzglnrtfl54ATx2idPfxpotBICWfkDpTZ5yDHu9AhhWjM8LjxLFZ177dk
zSVNulOvyEZqDZLlEsDcjhClfes9FqhygTAI0VoJDz1x0pKSg+Tc8Q5brp5SvhIYFg+5ETJqfeVX
cgQkbF7FgGTUxduwWMPS2XSSxeMRkWAwxTFbM1YeWrWbuLEZYEaQ0uTvxqToTjPf6zus0lEyRpyh
nN3n0gQv0trFEf5rrmMfpTht66BPKZWmdqkiaQapX357W1WLJ+6bhAckmC8Yx+QVyiG9/0TTwt3z
kbNYkPTJjVVh1XGrMSXHOFmWhLQEDEY+A2D6GwucM7pshJoz8Q70OL7ppNckIdeZV5bQKnYhvWVu
XRS1j4p/5zkEF0PDJ4fbRu7Z9VZd5wYLvYU8zVkchXv/mfYAbRfR84PVs6+H8ZEsy6Y+hqimpE+8
30QadBRFtOEjsAHPTF0IHClUuLmeQAHvJFidMSVnCEf0UhPY2Po6xyakm2Trlt5Z2b2ghQgkJqR/
pyTmkkfBIKzFPPrl/A0PKTYWjCeQ2TLnO6dt7tYmlK67T/4ZIaebNMtAwAPcnyIPnp2fg+4M8Hx9
Sz7DB8iNgjga7+1V9BN5OPyYeDj5LSx+UDuMHqmibJwlqFDsndgCqPvxRtebUrpGbAXmAcwMhi5F
AVwnmSFeifPrhj7DhdpKzUnB3yzqMhB8DK6lMY1OQUXdgE86s9RNQFlEziuOrPIjregcpBF1GaNC
js/RA7/F2+uPKnZ+7984t2x1A0NPVtQB2sYuTAFy96EHEVMUEJ8moWJyvA5v728ic+C2D4OJDu3N
K6EauGPfubyhlcrMEpl/Pil21NeNh5py93a2XoH4NU7EERD27fiSX/ubNfuP+GkN+d95iO3B9Bas
m1wOzQHL30cpmBSY38rR0NcXj4VcppVASaGCS2U9VGcDlrp/zX33nzpzEOsMEQ5D39/jgz5VkhuX
zIh7mssgOkor/JEHxOC7alTgBn6Ys8X7I+NwNzdLKbKWOORgES5l0Icd37m+sOTFkzi0P1LvLnxM
APbPSEwqVWipZvOgth5ZHhl7dV+G3K+G0syv1nlhX9Qdj4lDATeMnd3ck+kDkC48bVQaBDyxPivO
sFjSxd8o981xOEnP9RO8KT4U0u3KDRfzmZAHXxmjEshhf28Du7A3uJC5AHHvSqf+lhFvT6f54bgE
WDhFIYUf9WCGz3Bh/2ttvVY1wCDriVJ2UuUlMys5cqGu4yF1X1oGtuEZpcd4OLM9OsD6Ufd0ffu6
4C+OpKFHNfLWX8KubPCbRxT3Odal8pS5k/mBEXqQkNwneuihv17fISEwB5pbyHDUEjdBhSPGL37F
YLFXHo/vKPoUnj7KXwlCfm89kdLk70msEicBLkt1mVWdETobhSrgObWlWhn/DOqyqndH5oI85UlM
VCZGYdQ3Ks+HyempS+15/N9r58ux1Qsen8BekCCTkKf4sJO07jjdtBNj4OGbNjo1ER3SA1pAmOBZ
zH9Ir2bo3vP6Ioz+MKOQIhj3dN//2X1XaIUgyc5f3ITxc8eLzlpL5QDNbhY3nvl37ZUFIRt+fz2O
gADntWeq03xfR5Ubkcgs30ncmwlmf1Xj96XUX564eQAAx/inf3PuukCEDLFZFFhMjfnyv8chkGyB
P2+WXw5w9acs+tGe+AAc+cJiA68NWZMPc2rxu9O5RXWCGfPLWYeoxSpZA37a0p4NrPqLB+WS3vrf
cdnEsHyoSbZ2YutzbkVGPuoPFMdv5eEJZBblBxg2sA46fNVmnXB03JnQfiPCEjLOzi+dqX+L9JN+
aHfvpIXDGFlnMSVGGqtlZCr3zr0VDKcr+qxquIHzrzp/55NFBD5Q7gjlX8jBoE72+4OL55J/7r9S
oAlig1qPMPmezvtln2STMphCi/toKpcdGjonr5pZRfdYPtsJWD7pXZ4bQp3Bo9Y9VARPrupnHan1
i+EJ2kGBYxS/EAksCBmJLm0DttRYa9fsc7RFeuLgCtglbslSY03KqEK4U0rjOkMq99FJxMSeSbFx
rF/g6UV2ek2Crdk5AS11zyLysXOxX5iVvzTe24iZXbrHYCZwbP0ubU0ciVnV3sTpfnPFKWSysJEX
eZCELnijGQgp2joLVpRtNOPuts61HQoTvQbsrk8c8jFU/be242GfXamPv0n6siaprq2RuhI/YIrF
pwiCfPziyHyjhT48wQ2Y+ad/UJuVZV7vC8hAKJOwCiShb82pGJY5mtcUve/LrMtchKN7qvyEj9Dr
B/zoWA8OrDbUinMsw3JVUNhCRc0KbEqPd7YL3BAc4B8VfKFeirX5FauO+uFHlIJiCSBgsKyH35M7
iRw2PmOOIOV68W0Q/IcfJUbY8cD5eCMKP1uG+21+eKxh71q/OctEMsCEUzMzTH84k1cja8zWmoQW
Bo1upFXGVpFQcbj2Qch3WOGSeSkVLPT0dOKXaI9dVuQax9hm0s5aspx0zZDMsRciRTgH0HPw4X+f
r5P/jUDh3/JJuXrR1UCS6nciHPHVNCaVNaQ1J2VNzISktw4WqlbmJtEcieD1z3wfFTLjRz09FNwG
OqQlqLg93vD0LJjUgl5nC2ivS+hZ/fX6PgMhIhZ7n+4Z7UuBNM+kE3f5mlO2bFC12Q/ibdaljpDw
Xs7GdJlKny4i7C6Jwba/hxYZn3rZ0WhcIUGyO7UFGlgyej2UwO4osm5jCVFxoMydCm0KSpCBvgWN
Ht02DDNiUWaurFvVCvMEvek3A5ToRslivY/m+4d6TlQFNFcB3HHitL4u7sKQd7T77WlV9q8Au5+v
GNEQw7R+nxxLi0nSSz2IuaCH1PPz/GIw3TEoatBLAoo9blP8tevK0rAM2KBEfTwGFLZbf7uofOz0
fJ6qPbhbvUysP5O/WorinPB28S5huNIKYmGZo1/JAjWnKiCB5UznoAY4jwYisGi3B1EsCKfQ1wHH
okRjrVu8xctCeNTHBk5J2U7BcY8xSv5ajOjG/JtnmT19M6g19Q8Qf7uTqBRAE/ammkf8L+2HuDbl
pY91haqmL1Ux3myC+fTN0Bo2yIcUy2VKc31hXFeEnAiQgq2vrmufhjuq0YmA5ehHRFlxCIGn0go/
S/IskkVU45VDyh3kWtY55adMDLnCt0AHEZRbVrteQYuJOt+Bn8XFUWVDbdTNJMmxhDF5uhcqYvFp
kmGWJhSs8UyRrVxnTfCxB0O2M6JwzQDjRnjYmDQYfA6fn8lUfvYU7jI0l7tZCwGZRBA8qB12mLTi
HKOo30Ty34u/quSs4ZpYEzOU1I14vp+XDkCC1W/XChDZ6xXn7crFPv5T3moqvT0QVrIdL9ywEnZu
lnM10fnuiw/QXOoGmH+soxqPLy0mmmLWpzVRCDydCfDg6MXS/jO1oq3jnrgDl6HpOfzZ7I2Ylds0
iH6cthnLVnckbvWXYXUozmtTlnUuBX/eKuFHva9w4WArtuRjjQrCQDyqd5nJCFTQGXL7Lfl8SoWk
BGKLrNBnJf+gMni5PaP3KH2UNUevHzgdUVfMktD4X3nu9I489xBLjDTpJSu3MCZMtCxrMvMFTPf0
j2a90S/yvxwE1oRiTiKXAmR27zr+aQnjsFFb9pE6+Gjr32j1k5gweGJjgzKv0wqiBINCmxxqlw2C
Omg1WXmoXKO6GTpM5HiAgkbBPjfykm1dvtgMXG1CQ8qaP5Fjb8P/V/T8BVfbzcZn2f5s+IRJyS3d
E+77ecmuywAqupI++5t2X/SEBbH/Z3CHYxQQ7MDMCvSeVLN8sIvwXTOxYARHoia7pW1fpslehzbw
jUuEcGrqmKq4kbf5y9nWtw1EdBi1Hvmsy0acOHKsM7d0fl4Ia7aTo2ZoCvKw6wPs1CGKmqrmyS2T
5w6TbE4Y/Nlh0qYDdh39YOGBVRAScpanwmCero+BqJbbBqdu5+00sQqmZUEEsJSehuMjhJOUyK3s
3mBeCfajgGjXofRL5k+A7HAcUNQKJnEeeLxBp8nsyTGwmKl1yvfbq4q80heDvTlZ5akfwhsTYtMu
KMI9vfHz7bVgvJ5srbbOlLpY/Ke2PM4X6a3Y+Yd1f+7kAd8t8WLj0+X8AKeg73ZYoG06GrZFeHms
5q21WvDRIV9HsiElR38xuEIhN6LnifkW/FLrurPrHaw02KGDOiLglcF/D7ap7UWIXgrniuzSN+GV
zRSPyqWzAB1jyi7iJYlryn7sw4h4US08dOJ7OWi1si0iL47bq6WCFcMquq1Q8rCynuEEfCgb055e
FYZ/Dqa0IW1FgjvW9UGdDtDEAoSRvrIbcYej7cibVsRmk7wahSs+FrLsff5oPPa34noraiz70kpG
NeRgo7dAiAnbFpd0A4ZLSN4WVm/THmRn0GbBmOXYN3NjyiNZ3sjKiFJTxJv0e89zzwFlj4pdGPXl
yWdlRB9z9zn+3tv7gnG4ltbFjjUzZDXRHAOslyi7lQSXk5QQxSDZ6IfmOpvdctywju5rU54wZ6j0
MICOGixmkFF+XzHnAspYQStZ8qSEYx1Hh37qaHOVHyth9u/VJPqjC+gqMVbG71fpaq7eu+Een3fj
cjVFbVVOElt8An0uN8qgxOENl6YdE1uPBNJZXIiUkZhesuIKmjyTZBqB17IecmQfmkb0gT8fkLnT
GXWcOt6xbsjHf34sUcj0+o22+hY1XBKSGESK/q5KK8sR+oi0urECw/0ajHZ8qWIO5viRTbwHR5Rf
0yTz3CvpzV5RmQM0mEFkrkN8xs4lrq7fIbUYvC+up2qNG2yweRtuzv8IneCW9+aObeXCJhE6iGPp
ut7b4rBei0ar3RiSmDwqDkbVM9Eb3GlGWOfmuXY+eQsSKZBKlA6iKstJUri/Rai8C18esKRx1Y2I
upE8bbvBI9Me6njW8otKTtSuqffriCkmSt5/GvvJ9h1dEnOwrPe7NJ8sTsDz3EJl+PvrCR2poiNH
bVV8ELjNlFnUdIJqebkYYrKmd6fCfHJnRWhM+JflJ06hMx1LO7FuscVj3U53Iw+I6ewRkJ18NsHF
4jnwr01LmoGu3u0KEk+39Vifa/zdSl/+kJS4vJhiWa6/HCYmEF6k4Q+b+S9M957eRioA7FtR52Pe
qoZD1rtjH6KlAAwmtnn2vDIeW+xr2qSCIKD4HJAo0oBwRZuZL1iPCiCWw1SOH7JUIo2RaoOo0BC4
HL33y2kPjrrc6XYCsmZtt3pgYDSToDk4L/y+k1m0ZiOfTIetC+frz14Q9YkxAL6unkU0pPNNG6PV
7YQ9gC0KiPBkBEJsGUXc5G0mAbX+/1s2n7EmZ6+kmfUftMuAu/JwFNDP0Y52H1hxOBA3unvtxsOI
phqdiMc3YyfNkE7N3bsTtZC/bwOZsXk8gCwZaw7FxG5miedWAU39HJrMpRP4Zf8RJdsgxP53/jB3
0/DRrwO7fbLac6S2LBxY2yZHfDcTEUo24ZBTUh4rLFhUMaf4G+T0E5glRflCciMBb5xLgdwO8TWE
l2Xl92Y5K+r9E8L/j5oCbqcgYwtT/KeYPEYika9tpFyXMsQ+MJDH6eLebTfdwnCcbsX70iso7cUD
ldhNt9r82KGYClsxXpJNNvI3vDcNqbgNFDFoy0rjJeV2E8y8E2T6v8YbfPiDxezxxvzlNJU8/UOA
aaubiCDU+inr03D0utabhzEzVeGBOyumpVDVlag5ppOqpceP6ZgO5clcI5ozlxsf/jOjHSdcHnry
gjgV4TGrZpSk6/whGwQVzWItHpkNBFX7269kyzs1QGVJyp3UhagfQYA6ZxNj3CHvhgIoT7HiqxzJ
OEMUAYWYGU0zgdZ4k7+NPrANGjdbGpmprCBArk0dfzvyZCyuWcOA7Z8Ii13qqo+yH2xtm3nwBMOJ
nAZmGGh55x+aOwcE8bH51zJ9/8q6AHbju+OzTgimp4cDYVOUpy5WtRpZUYDDfkeRmPfuB9rakMR/
D86l60ZOU3a3x6JZ7oIjT2lkTc2kbxAsiEeoi6eenyBQllSjUYO2we11jPytKfB0rCP818rzBt1S
9PPiOdt0/SADYCTYrA3FN7sv2Q1HoORWFur3UHfF1Upk2olQ4A/2EaJAHWBxbL1UUw2L/tFaLsl2
gtDwTLWV7L0EJ31WJT5eZ5xpgwzKTQqri4iuShb2kHXzFAD19D+GSC1LhUj47x/cNySbM7IEu5/Y
KtI6RRynUn9gu5h6kVCM1r3ukAGxn/QmGNYB6ZwHBl6wMDT8M5FSfluLwFMlW36iDXwPgCQ+xnCd
TqQ9u/iLiLUH2iezf8GxVlLuMK55rU/E7S3YFtihttBnaCd/e+8QoSXSzXX8pEI8YJ8uKs8cpvut
KKGbFiYPzDP1K8aVQqUxMnJ/PklmpOSN1Y1NbmbHTmHw/Q7W4ObZKTA3UgTElyJ7D5uZ8x2vQN4C
xp9cXIhAYeVmS5+LZ2R6p1S/RlbFnGoJ5TfflKlzNKoJYlp0RGyj9eUhTN7+jmlUDnjE9/5yY/Wz
0UVkLu+HtlDl953iXa9Op1Zjl7HqXgSmYAZxAUhetLMuo/wIZcE6MgYcVQXXftaJ9FByHSd+rUYK
+QKf6adh483LpsmrpQD7gzils/nSTAGpSAx/ocCQfCcoIQBObeUhzNkVe+GCI4KGZnTW5p6IAKMW
LYp8QmlIBVauiA7tJrCxofnqE3J3xStbmSRwWWYt5M8C7AK3V6g5MgmZayz7s7YMNVBF7hASg6ne
FGWfbt+9fP9BKcDeVSqpJ22Jpyc3liY6apdyn4vKMMocNDmiQR6pgqRYGlSvonVoWae1w17UZNJ0
WFnV7bsFgexbPJClDd3OP2/OA95hg92x/fehv51zCnIYEDBt6cy7fhZQp3Go26vuVLynnPj3BDwj
b8gShQLQhc2FYnQlHfKBdJeYK0ZoM5ZWC94c8gnowvBkZDleTJdaJ3tO9tf7QoigcS0waqNaYSDf
61oA3sAVTSZ/UsS3cxwkCUqEouZWVqpdM+gI3TZH6PPVwQ1eeLJBSND3djc9o+LG2YvuuMJPek7E
A1KPtJQqrvj+dkiby5CUaQFWHeIyNqlBxI6R5wNuoYDMMYXG73rnvgPIAjGEOT+QJdZEzGlJx2p1
zNSraNcYKzX8kOkebG/Z2jlqs/xbFJ/MO78q60HUlQWbiS/owPVzum81gFb8mG/ujhWw5a75OCFP
v2lZUDgg3/gj+Zu7POa/DUu7QW9bykFKiu3fVbr4Ko9PyUmXBcFNNNm9Pb5F/q5UhGhS37ZijTMq
ijfGCZoq8eCMCChAu5G6pjKYN9TenWD76RSm941di4j60c/gNxDHUdEZWMfJfIPiKiDn8rPVbRMe
mwux8MKv2E4mEcig6RmkscksufEBZJK4qyjzZ/U58Ev6ipPgUHnXZzJkJBb37fQbZtDqL5O8oM8I
aKOqZtyu/7zxfCAHrdb1uPD3nmmENSABQs1Nu8qrOVljqKDDsVzq0ZeKyv7NXEgPkIEe4XEa4hiD
qhzl4l1iDwg8AAeGMw+NZTZAgpe+pRPBECGDNE7rX7J2Y2MISBXEG0h3wYO8Y1sOs0s7qacMhQ0e
lRapUZ7gr2IPrI2JSLl7q4YFSX32N5sIqMQIcpt/Zc+zGc1QnN5RpeSsNxksVy8lqj0J4tniM1Pw
d8+9oAcAV785ZZI8GHNYaPt2w2/H+ul6vB9Q6JqyWD5fXyyjzvedD9T1cmXtX3XreofaakJVF6yD
VdAGiHrX37F81pgmGVsKL1vX+TFxVY9wfMy4/q3uSZ273180+y4UQzzbwopmONRKbDVZNObjNlPH
ncdFQ6XIWzTq+wzxy4jg7Vb8YWaS41cDc3CwrkvBPz5BcJelAMoDcPhAKKIajoJ1FZ4a0HoGlq7D
89Yvf+/tMrxI7p3HeJXvxigFQkf9nyVXmtj3YgQiXUs+AMYja5khKAC/nwpLea/LqVeci3H6t54e
rAHbvyUUzCQiBD/cS0cZGoohduV+3p8YUrMbn1mtOLkZHkA2fuQDlBTi++hSELYX7dGloL0hdUWl
1ECPJjej9eTgUuoEue4jPgrjzikFh2uxqbJA54ftuhjCFeY2RWabqCVWiytmh0F5l7iNt5X+KztT
pucGI2KYFJaAQhlwh/P+BidUXKMohG+FbjXS5iNQl9m2u7B4nCitSnFIFyjYE5NGm1tMk2n3z7sB
UZEMEnM0xq7v2AjIhjWo165ATEvvaXEWUVwBLoY2+KbB4nYExo8k/P5JTLpG2DquHYFVGK6r9yCm
bzXVF89rjOpoihy6QLWF+L6rZLLS29S8CpyD62byp+CZfPEcUr2xXyQ4hBYwAa/7OQ6pg0z3a4H7
fIXWaVwYOlceYYVT8y5KqURkWo71ruoryVSAnWyeEcyMDHXXTuvjoSemcuUG/LVXaV4F8nWulJPq
MW8YJDNO5R1erjTKxicA2PHQU8VROE4KLLV7Ami35+3Ttd+T7rw3dhq+0DkmTHcXCX5vbJvtHjpX
Rz917Rmqin6MDQP6SpxdnF2q58baFHWW0dbodmhjo930OQIS2EYac9zlAcZkRuToTD942ucmqOe8
Qx/zcZhIlk2w/zzYeIRofO6hiqXbrPAIveyHSO1NF2ura0wGUGhdduA/FkramwPwYrUmYrsUYuEI
xPZuhPWZbjsmt4VBmetUplogn9n+DkrNfKbEeVUvbOe8BZGayRK6ndTW1h2NpEhOJ236VlQ/Me8U
145y5MyTIgMhd/7MQz95kMfSiDHeCJyS3U2pcVglzFW4ISNQOf5x6J/FaC4BAIJOQBVBLPMX5HtI
IsOYuQOFoUNyHkkTaLRy+/haXLy+aWIjfkQvo9nIfpcnTI8UhrVbRx7cw/0ymzJrkvYVk+xvS/i0
lj+BUPmdWIN249N+lmrDt4Z4C7Naw/L3iNRh7KW853I1MMQD8wOKWnmZanXVKtiA7BiBtZupK5J1
/kVg7EAm9kwO01lvoP/2N3zD8ILvq3iuz9ALm/zlCGVGNYIayNdOpU+7dNneqDMDCQcpvwRuYtB5
dBPUkVCbczQbwIPFJ4q/oeOM2E5Fmygbu/dwug3EWoVHTW76yyhasXfWl+N8UP+Zz2l9Lhisv2qd
klEm8LrA+oPFkXyT4dzkc4odcH6Jhcg40+QBNS9nmrHx61fo12tWZsas6gTkcGMMmKDhoobM6f3Y
YXJ+4IcbipKIrwbpAUU6Y+LFpCw+amXER5UFtWUyTGSny/GYcjie/Vhqz9T+wbCd33RWbZzOpHC5
YOVTQIHNQBvli79IuEUjHK+d/d44bMqatRN6bPpilAr16ve6s0dv2iFZCm7GEmx7JilEL0v21fYa
/ZAux+Sx0QXpc5+8+ffZcNTOaDalhUTDRvCDPHmBh+ckpYvngOMjvHEBAyoIO6V+Ub6isT6X3H6Z
bK+GuvdzNWTdT9gqdhy/8mGtRyxMMXVUVN75vYYCaRdzBliiNHrP6mJ+w3jPOoqG582IiNCmdrjV
oLylaUprdcLqhBw3Keik0anvEE770P92tLVX5IatH2IBUsgmAYhgRvezGUsrycid0VaRMzNN7lJi
z6nJbiKRPD/NfwUTNiMvd7uKWLcfZjxOJ4REuUxiSxgL5okjC/MwgW8BeNm7xIPsdwxXiPp8N6+u
6ZPVx+RAMMpKKBMswgzysr7Q5CIGsaV7iiaMKxf5M2ZdteDFjnou5ihtFk1+vjbfbjv1AsNYtJko
KVWbix6oX1suDgJ/taEsiSS/E+IYhFpL+rpM7N/OYdcxssj8yopkvyQge5RWLWpJuRyDZ3MwB8lh
Q7/X6Dll6BVcmEYKl0NP0XTCb0hHHXyVWYbHYG1RtfZl8XyYiQoeHlt+2xdOKG4fkMzKGdnuWxlE
XN4V5NkQF6wM802KOiKP2EgaNWVKar1DKcyxHeIbxdtRtISK3zHevJ5sPg70VR8WbsVZUDWsw4zq
2V1cMYf8KJz1a2zDLl2tiOTf/S+rbiowDCJYvB/QAqCz1dA2ORckctMrTIyLMUS33gD/WORq9+z4
5RM8zkaYJJOO7TfI48naAo3UmXcse3PkWtDN3kwBQaB0qFhcEpzKSKXWbhhfXxUbk7lrwDlzqtN1
unB8a82/MK1GbRyNTKc2c4dt76hIxsjXm2unskB8GETFjYCPJU8+bP3hvpSkgBLlMmKRVCHlebIY
rrm5NmnWsnIyfANB9Q43NHhtoITKMm+2FbqFcdvYDFqx1g+EF+EcTx7AWp3mAx++lNQ9xQSQFe3h
Dk8orngTGO46mtp0yGZkd0M4+fkeBjXtXklzs46FwGY4ekRh3zC+xnTlS2pdCBiuqn/I62grPkdv
Qq5748ChA8t538Rja+c+pzIda75S6a0lfjAmh8SSvuqfY1REEFbj4cU90ADOJ/7Y2eEqmwXtCuhJ
b3bX4vAfta1tz47MD+SMQ6juo5BRq3yiFTl935be5UKtf4e3HouWn0gviQos6xTWAnEPeitL1vT2
ow4W3awUa7USg7b04DOB8e0FkYfsXrHJP6amOe3P0crdi13RbvttELskb2n2SKeU8umWqi41alGy
18/8dHK0ecQKM3YeD9Ht5wTt0AxXlzTtmar8+8NYK61G2f6j9060F+2ESdA1N6F4c/qJIPtLd1K3
RR1KhhWAMUttsp/dYcc0lblFvW/XpJHXVj/HJ/7hwKy8zVDvKCWFIohUISnZK0unfuu3DPiIX4sT
1ySMKH6bsszoOEYd8/6n5H3f24AKo5k6VFI2v9sA2+OwtT2rVNiGZ6lyApcpo3RH6ftGXKACMatH
dC/OPe/LdOCO1Lubsji3PHNKK0UHEJu7V6fqZOqqXckqV1HXB40/Vc2+Z5xK4YGpyfw0cEarI8qO
SRgukN4UTy9ZsuQAJ3YPxQoUhu6Cyq3NLfuKkGQmXi5771ZIE2+jVNWQlqisjxmsE2xYnc1+Gjmz
GnYxF0XqNEKGkHOCq/oN4Gwb5zQuFY6lihIdnnayKQdc4UqbNDsn4z8GSHkfgwXBOe52htzDdh3a
HiKKyZgNpGhhGlxeBhW/93ATnlMgzJJ3n6DV1Ze+IxyEEXhyvUIOXnEe20wU3cW3uJYdiPEMy7HD
mj00MTqPcRZm0hx4gYLewzksulqmLbWIvMTSVZMAYUnIltOeNLak9ScE6JWviIiljCJ51ya9A5Mj
KKI0Fh2JmDMH/7VWJu9nBfnIwVKVSe12+NyV80wdVo+XmgNZjvbEGOA/k2VOU4qNuzxRj0kfLQnu
ZRiPnVPsSYs8f0g93+VsuugzqDiK4M+QoFCto9eYKYnp+1T7pF81Plx52ilNTByrbKKubhKclyGf
3csNaD5sPTT/sd2c7w6CbUheEzlc/zvETUSejwnaGoG2jHPO8Q7RjagdLjVdgcbHSJuKyoUERV28
1zZG8ZlWdB7HQQ/h8AKO/0BJ4A4Sk7S+Os8Pz09yZGhUoTZCdb6bw3OUZ5qt+WQlyH5/9FXl1pVx
1wFo44hvDAwTcIYgVP8hghPysn89Cn75fblqsKT9sH44Hf4l9uQZNy5beTdHScpEd//hY+v5sCeJ
UF+JEwFQrGLyNbJWSHtrVzkXbzklPxMdnIJRSMe4hDADqrc7+B4V1ZSd8gKJkKC0aNrpCNvlSvqs
sBu6z9ehZs4dQYftr7koRAT5+QMw/YwI8rhsTxoX99kgAJ7ayifJR64pB6m2cHiuIrBIS/7tKh8v
w6zplXApimyS/taxRJv/sfLBufXE5Xjghzy3gZ7nk598jxVTwRb5R1aUaWfj/X8mfWx4RUz2TgQQ
CI4visv8D8g6kKKX9+hcRVqlAc2jkh+nO3VffC4E54wev287HBFW3S/LZqUznwPvOktvb4CAhRId
Kx9CKD/3+hi/fb02ZoRfNZ5GhNaeIKQgTNFPCq+Sxn7L0PbYQ54yJWAdO1PWdfRff7yxuGoOh4ry
BvUdLYa56Khm3NSKZERYdTx6oxv1796xObXLlVbxlvaJxWIihkivdplnr7b0ptcMsDozdUiTu6US
XbnsB/6Utx7mb3Is5lgozX/PXQ5TA6AFAkMDf9rQ9cNqefHyifYZ8F6VacYOwZz2mvcReEy/wnVq
7tiVGYb1u3ADSsOV3cLGGG1Ny4mW1yap6ppv4Trqm0E/05G9ukq4do7kh31rmhTzLnULouoVIO/M
MaOyTAr+ji/47WWqbF+B89QwLmM6dyugDS2GjZnPEnexKMd1BU5KJmAVxI0O/XZM1YvmqD8ypRHR
Jp8yrROD9aIQoe0fYoHK6RU3lq4rACwpVhTQdu7Ur52T/qhF20a/nkfO5Q0DDZKRwa/j5SrSFNJ1
fPT9WVigmAZ+G9zF7AFg1+Tw5RncSAUi+0H7r8hrCGUpi3CMaRK+ejg/SAllLvi9jhuFmltrqnS+
jkIwh5W1PFNUPfQf6gIJiu5HRBnRQJ4ZC1IoB6yjeC7/W9od6Ka5NTjhLyp9NTtCSh3+4C8nHIQL
rUmCXU/2Cz1iJidFlUNLwTHhqcfH3iwX2ouuvzTuSWbixJYH6pVAJ19Q6ECgb0mG88zjG8DYGJU5
i0A6NC7tpnZwBrWd/LPa7BaUufxAuGFRAL2pleCnbmN9Iy1OrEebgy4Q5O0tiBluAYKk0EB7yoUd
YxoDCvItszPT0IM2fhd1NSyc5/PVmoAg+irsfnqwkQoBgTy4fszTl+CQLcmRx/j6VFlAlgTvXo4B
5s9/j472Z+UhzvEhARrrvqpBXPZIEo6jct1T9r16KQbFeAEOcm3ZiMKO4YKK3S1+ykzPyA309hVM
MiTaYZGx+HjKRf8HisYDDvRlJV2WGXOz1n50V62R9EMBX5Xh7A2OzZ7ve5GfEsRNRmznZfZJt7Jf
WxOXEJjsf2gLCqRCblr7ea5E/PLdxmWtUN/QBF/u1UU4z2TA4s8syXmNLeV3U+0vfcKW16sbClD8
cu3pJVxZCoDaabc8wVyEiDh+RZ1lKfMBkRWU4NUgxlT1cRvTwaHeMIAUh1cRj43/OkV++Z4GwAkg
yiAORwPIt2JJCYjuo1cHPuy/QPidebFW7UPNK1AzQZKDCWlNqTdMCkFuaGSKKMlo+9L/DTQksvTR
Gqv0tR62zjNsSxDWnd28rgwAGoZ2JJcjnPN0OkfqHRvUGCkZhJvnvSWAJGkhZ9/XlC6tzLOFzJIn
0oscufi/H2PVPiSYUsENNCDMEjTlnTnKk77CEU8wU50U1ApfzXYd2PYb2QD+sXvfi4VA9ailcubh
wM4vRh6gVlMF218Yz3oW89f+pF9BxEkeQ5wszrZnAkSYVY7dKrJSI61QzAJDGAcjfCNHxrMf/Pur
Altc1+okhy1ar50miYmGY6NL9lse+rk/A7TppzmwQ0kyOlAHOdt+iEFkgklw8TYUv3AkCDs+f+O5
JMV6x8VsICS7u6DHil0nG5qYSeppwI0wjJD6OFxqJ+1pwfh27IH5qZOMmhroOnmvljuCtvrmTNLd
/PC5eilxTprVHyotzo8hq7ubBNvG5+4BXHTHGDNQvQxTJkkdtZO0W0m+dJRbYk8FlhNWzv3t7UJd
GRdSsPMqkKfV7zvCAugt9Q89es3dZ9Tt3ZhyGjUq6G1GMXBIY9s2cpD5rqDrnnh2Dz80+eumHd5M
DXNLYg/YMVuPCa1YRNCJjShVohC7xV5ro/xtjXPq4pvUMau8WZTux2R85e/eHuiEgUs+LNAdHSRB
1BM1LQgfnJg3KjEWOtf1BcW23GKJjfonffpIK4clYh85l8SYc4JuCUxr4B8m1l9TINwNlua51+gL
IQweU9C0GqT0FFb76gmk97qxoZaPBS0/GTAGMv9DVjYY/jU78oPFdjCxKGHV82PPUbyPfiwM17Fr
AY496UwqKKveJvxVJCD36m7ez/XgVRYOOXi13jxtddcP9wsohHOO/COlJVAD+ahqEWe9+9yiLu40
svDIo55Rz7bKAqZr/hTjNWx4wMh460PANYxpoxO02O1/uZQ18nbZxowWJh03A/I1y4Pbug09N8l1
TPjxiAgVJcqqVWV0LPOFhEwZSLTUOHcH2U6Uhkfie1aoszBWKpl8hcmxPiNKkSVWaBuElIVrMHaO
TEP3PysIBIe1SVKn16YxZ6bbSc9SuPh8d2ut6MHqtgft8tIOO//Li544hrkhvplLJAPlL6myib51
reiQA4e9wLBR+QJj4f49+4RecuHPhpOqMcGjQyjxEpUeckzoorZKS2xOBYZ/0HBY2F28K8QPEySz
0I16GxT1QM+C3xA+i/8MHnWRnsLXtjaokZSMZDhEWaqTr7ESSl8VLa5HOFV9oQKBxkLqHe7hlZyn
1O/y33PJAaHtGU9s5/T0OTSWwlv7AhVJoajrf0P/57B1w7mAQxs8xHLoDXl6JxRq/m6nyjSFmXs9
j4Blds7DN0J5bT7TuxbTUe1ptWp2on5wGwRLh7g+pmQrMKD3L8O0w/EXimJ0/b2CHYjFp9dFumpQ
z++oESXAJZFlmmoZfCrzQmFrqAMLhOvrUw09qFnWKfEedFRx+1aG34nE1qaa2jpGFjHNnGlR8Neh
wKNN6YUa4JYVcHrvloe3O/mp6D914L/nu9x0DyaovREYLv4feqWRdom+vi6ct28Eva1hzT36UawQ
tjJFp6mHndMILSoLoXpbVQuRMSMQBw9ss+5sQed7rvpifm+Qh4H3pUbCPI913Wqt49iqm0ZEuDSs
RaeHJoYj+L4o0JrTvF5xkOSwZ3mIbXvsHeuPTceDIaGbG4A8l+9WQzTgL7gxIrUrgBW/3BW+7HGL
RGXUXj469smjAWDbNVIfDXpIfIckib1ZTgude/iH7jzVTTw3br5ULmkAjR6cLHjSIMBjyUdrKIde
RhDH/KOvkrqsPTEEPw+44sOGl3/UPbQ7EY3zt6MCL0n+J7dNHMZw1GR+68nVHo8+2EebeGLJITDh
7+e04cZMcPlJChXCddKOy4vBeURUOSIfTyWdz4ee7IE5lXRVshY7+/Bf4KPOUiCNQmBsNgVlqm9w
LaSzRvtt7Kv31Rdv+HF45sLxzynnwJKKYDHgJWFUwIc5Tud70/rNx1nwE8BKNOjcVkNrNsEQoke/
KEm9QT8ICM1wPP3kpkBe5Z2rz7nHb+qqVbN1pP/jwBcH2XXQmQximnuP9rMBsmx8O6qfd9owKwkG
XhEY7VOIE0HaV2YQXHnjsMcZF08W2fTSVz7AUao5sSOKUDqCu+SEUKbjGkHNDzOtqxcIHUv+Qobf
DvqXVBgVnARCY0qBiNCae04TuzE5LtUe//6PYDzqqEXpEuxYC4TfbIOBVIrYRAjvYy63xzUALMtm
H2/bNxXNVdHRpsC17JWfU7FOC5fbNRqj9uEOIVxPfYVTUi9jgcxpSNE2hmYuOcuXEYm2vkgPli5X
Oa+hflMQM9jEUe+2o+C3iGlJKeH+TSb3TurhvvfdtgSRm/iHLjS1fe4UDq9Guo/6pofNUk0t+iT4
+yb3pvHEiMEjjX6doNsV49GUvbfy1vuTADM4Rx3XvKcY3PEpbrOxgu0jPiR2UhWb54v8t0ytUyil
KiNHCJkNYWhYnprhNy0n8EVQ/s1hcACkAnj6EVDoFAJ/NIegiMfblTAp8qawaNMXhYNayE/GYeTp
olKhaTaiDZkOMJqHf4QRvJARPWIfX01Dh1qJhmWI4mdcH6UHVMWcw3CeaBhO/ukwftjKbUIpi9K0
35EDx+SoN/YXKmMllv+aA0ZB3+IXhs61Oq8XPot9pA2L8PqdyzM07SVy6uyYe36JzRkqUi8bqsML
FmF+p5kwgKzgbIMZw4VP2pAU8gi4SZn5z7scNmZLCCf1Hu4rjCc+tm2/eOXFUDUpSNzrCmRVnKvk
58huvyMOiwD7Sff5ev9McEr7xOFNJbbaqfTuhmsUdkYkWawaOVqE/eDp8wq86jtukyULwwTZc2Qz
Ctvt389alxEMZ924mwJa6bxi/iUu8tJxWalobPnXDpfgHILNcoDxiUJWpAQT9c7E3Cy8CCFTVkoS
YzZPBCpRmUjtgPSHYjlj+4QlGm8e++278LpY48V6U6e6lXZAY5cL4y0vzOduAEUgGp6UawWYKWDc
irDFd5RcEr/TyVHggfn61E8BD6UvDtCw7cWfjItG0nXiNoMgj/BO693lxdAr3vxrTvhigbhb5bhI
96aB/E19EC2R8DUheNGb84jvIre3WnzoKnCjTS9Bz3ZYP4SCoxv+rri0/fW0e6c/FFfhWXk9Gs4I
5cuttQaFebdiqQIMA+tzn1r43s2LHZJ+tyPVHYo0TkP4lPv2m+OASPX4WpznDBBUdBeqG3KHaaM3
wILL4qnqP8Ak3KADDO0kC2n57CcWBPD7sPPfAg6xXLUEASeX6K9Gl+VEXcqUYp9L+6F4p6tZD16i
Y4Nd2WPGH/4iYNos3C0eGT6QTzUACQDtGTH+axzxjyPcfpPD1KngDG6VSc3f39ZUNLawov5jatrq
h/ujcmsHD/CexqNTlGsq+YAG9RKd6HKBtNuVebq/hKc5l0GgeVG/0rays6N74K549LRTHomkpb87
Zfv25tw6cE2buXa3tP7tlN4QFKv24zZ6x0YjdmRJY1HyFLy8kxWdQkRkVK42ZFR2qmcWs8QX9uxq
UazbmCMPefzRffzScZOEVcFv/M4GwxPbt3Yq97cfYa/dNj5g7qDQzC2tHLZHVQI1/da63Qc0mK0k
teGrZ45OYRMLJmejkMxta9En+VI+BsTpzUYmxD13pDUQsqFJd6HKDQRxV1iQrb2L6UME4Vss8kXu
+QHmHqHVmL/jRTjDEBiivQMS+t4q+gIk7xDk1CYiCHZMYyHa5HedwOshxezNAftPiZONXGPSoRg1
T7/uh76cTxc8+FzPUPrXdFPKV2Ra/Xk9I1d+Xo4KuzvD2zIIOd48WTDECOQyQU3p+nhRJmBgFU6c
8oRojG2pSnLKAv+4XD7kny0MZDQq/0cyV1eyYK22e3026fhHKB56Un0+3r7h7zeLTK46kZDX8j+y
5AUB5MNw0ezEaZgCOhFlaBRqCZxwgrpC7z2kZZowCC25OOvtD5LAVDdKLLh0m8ZjbdRfpJ9DfzVe
uFyyjN8gdT8Ls8CK0dIpfV984Ay7bKUh0BX/9aHMlPYeGzapGrBIKUGkjFVnM45xrtfRtKPmneyc
OVUlV/MmN/giBZgr/PZUiX5LA14Wc5N9Qjx6ORDpPhi2153HFcF1irEJusUkeDe7eNLOELPP25ue
KmV5k5URp5DPvLHgHr9HyTOmjwA6JYK/p//EHAMdB6KL0jCcFDhUNdkE695sahFF+ron0BQ9d+Y6
7sxZngXqrt0bOkTLbf7To0L38uGlbv9+gPgT5BW3ktaspZzVuC+9AHNp/nMCmgRmKTZ2cphn2a8O
bl03SbSt5zyZVfV1RhNi+ihNuZQPTtd2QbMnHS62bvLhbYyL1Q2CnzroEfWndmRztQKx1IqI6FfL
rxcbYxvsDl2lNZpE0aIAd5zPgyv07C60Z9kxYc99ALpjU4j29DMibMVm5/+svEdlm6+K3XzRyMGY
WnCAi+kjHiBe6vsma0ff+SlSZRwiEZM+4JZfvuzDRmudJW9m4R8Wuj5OJbEox+S3HgXekXiEKS91
EvRcdgYAGsBfUPg00vMFeMOvDtZQjuDmlWyMJ4l8WSUo8IjWRAvD5v8xH93iIPwK4JYTvjRkMk03
8mbdlquTLMqSRso8y2cfwTqZMrq+8ccqC072bYCDh3/dtmT/nt2J1/9XgN2bSDgD5OUpDBxICt49
RDZ/qpCDh8bYNAJm2KxYJuZy806KiRfJikiDzMqaiu8sMEkhke34xl29kV42GYBIT3msJD3xwxsT
0MftRDu9e3Wq1TXRe2pLv34jGTvmuIpUhjkJOwSg05NZ6V0K+D2RHUV7/mhUG2T19GpPgojJtlMV
xjmV7hcoBdPDFaqYcniCIfLUNH8ePaZgGMevjN0o6t3+UgCnniJpCm/TkZYs4rHKgNBztPPWBJ85
7uiNCAZ/LqeT9lE1Dc1kJtQvuSNsXXJWU+RU4a8DZR/9XnAhacKQbE9tfj/Pt7Dk46OB4vQodvWw
veqXzoO2uSA/g+KZfAhVs76gjl3IvywMUWVTPFxs3wT4iNREwH8ni7QBHJ0ae3OQAkjdDNGUPYTK
MOI+EFCTBLUn9ulneS652zlPtvlYNZtNj9CYhizgOnnyzRyJzpf1+CDej+wFs3wG1p9GvZv88qPD
YroHnTAzQktHoi2WFmMj+u53iEap4P9N/wr75lLWWjJ9zlv1U43oyfBL5Ph90GhU6TBsXaHRIbQY
ZzDByOZHw21I9gmHS2XNMxh1nd2t8QJM0msbE6g8Ban2kUb/PKXIV1uBvWt8GKoNsgZm2N45jCZG
uYTRc62vZ3+yxh9K8VKFmLALR8OB/zCO4ow2XEjOrT2u5rvuIj1yDpNyDMjHxkxyaxjLtjdGM+Sn
qrPc8IVM+TBarOaUudYUFiIZ8+w6J5lVEK5c46ZZS09VFmDeRpfDoBaLXo2ckWsPUWP2OclinFF1
Gdc60Nb2jAVLXu8TDKu42lDy2YCgkPaPzmeurZhpLr1x55o3urOK+x1TeM7aOddYIt3SWfJyJ0VN
YkytyL07MkvtexqaMu32QbDY1d5H878K1ZJcWOQz31tR37uhKZPkZMBmPEIX7A/kcmdQklekINLM
xU7J21o7SfubnqgibYJiqD6S7JAML8WTBng7k42FKCO7NY0Dr2/Wf4b1niWYkCI1GNys1+yxEcbq
rd2Im7SqiUgLbEL1lOSJBoSuc9TuWXDuJ1g4J1uqiEVj+/RgNe3mRePcpqrJS42VDI3h/ocjnugQ
R9zGiZRJSFoCMeJPNyEY6s8S72oNqCOfOHX5oGaugFXpwURISE/5o9LkADQdRbTA/CCbMHOxe1rT
LXY7DX4RXKMojcGO3B6df/pVQBV5ykhnOVYKqjsle/mPuiNhB1OaA81YNozXTbTbWz0Jqf5bSeBR
vgpW7RR36LytyMUf1r4i4nf51LBIyf5DnP5eTHZ7IuwkeJyRuXKzrRQ/j4CxmA4eDlJ0ogzsctdH
qdT60aRjA3ZmDoXvzl9dFd89VP3seZ86sp5iyGrMVM+09NpeZSR0TIIolwN/3A9Uk+gwGNJul+Yu
yrdgLTzFpqD2jPFKznc8PS/YP51kQvSAs+rsStbiHLLi9dStaxPprNF60avvHAQqrXPYwgrMlyG8
TgmxWzIuKkH1jHhXyB5AKHsZ5eN9deU+2E5VcEv2K9pWiWgrtM0cUNRUQd12s7A6It+v7DpR0ETY
I3VFSlAFTs9ICp4lNyTaEI1h0isfsLi9VGzy2uuuSvEsduln1uqY3Bpjp9suKdKkvHN8YZpHS85J
ImpL4McvFMm+x2szPSHNkOMOCVgpFc+UtZtTJGDm8AoaDrM648m8nzOeBhRHpF59/bAXadYkGGG6
FVUnbKKReqdZllmzZmZRORnNVGndAGjrmPHceaAzLmQKn8HTl6xF8nIlhph/NOYWUjAxBVzXmYU5
zcF4TCGysnTgiaP2X9Pwb3OGZBuCuURUrtwLwEQDn/8fQrrotz3sZmzPydltk+hK/W9Oix6IX0t5
pszEKSkir2tMTWNvbb9ifNnyDYyBxuTxMOsF12M+2NZlwNSh/LDkSjRoLdU6GYbuDaWWBYqJ121n
zu1Mxfx7NjJmhBAPJWFMCcbcBC1enSTINzs3n73FKvuR3m5aU0tdTWzz2x6RhAg8WcjC7zjqqart
mAYEpH+4cIDksuCOt5r7iYaiiyXjkkBh8CL9MDrg3bOP2XAn+3jU1SbfuAOebRGkvOOTCTUu0TIR
Gox/imHzo+ZIQyPzvgIWzDRa75Z9Y8KZEToS5UsNqCXKzFAVKwfsXNETG5VSMbcoxrSvpd2Oa/qE
5SkAnW/7KAXDa26elC7t1uUj0calh1JbIUVt3YnXF8FlvWJEChcUjHuMBvYIo9xs0/OqQ4TM3InG
+AhaX+lHayjkLljED1/cARIO/QL0063I0XLfM+1gqlUu+LB9zB0Fb6VkpNX+xeq8edu2AOStdlLN
tz1cLkAstIkmSIouHpytRjsQ8sGgoABTKHJTiwtwYdhMy6MlxUgPalSuU8CaQ2BWBvcXIhPsBVt8
gjcG/owPB5abH9iy++1UNRqd7xvORGYPU7a40JviDVk/zzo4YGp9yP/N5Q4lMgLkxezgLOWzZIKP
ku85UZ1L5vpKtbDhd+NS1+fqXSZ2QTllbQquNuwCpIGSDznddw7oHnk3+M1r5ys+2LJ26br2SSDz
LvHraUZ0NBVYweiWcQgpLlQluxrChCs2F4HHhbzm7ZbjKckXYx6bp+CAhzrpRe0vm23xiTvkqpjV
DQaIDwDBCnP32FumVPddfiHsjQCuLIf/g1TExECkvT6gCtQKNcVlz/cwWKU8/sZgLYE0heKCpGvU
CMbLuICmDgnJ3y6LKtEjndxS/QYWwj+S4yRf2O78NZtxuBJIvJ0cGYRXvyUERaC9g1R1g2xhNhCC
DeZKf5T3zxA335+FchXl4WnpMXtlEaAVDfSpYGGCG2W+Wub+C7n/PPebqq/d17d3dzWeJcwH4c6H
veMA5XaiHYtCcUW9jByM9khvz32wQWEhSpl7vzfilxn+QWPLSqepPqjrTBRO6LvrRbK8pXUzMLsj
i9X00JHRQ8RSrs7ePM6814LX18qNDIyv0aK2LlRfM1ecWNl4WRyj559aNMrhb63sb0NsjcVaT0tD
K6+M8A0WpWVIpm/hc1Dx0xm2cjVzGoz7b59W8U3yooffWI5hoWSoRI9TPr/PAc3e9XBZNZyRxsXy
Vkw+iVAuul/4HJcKAizG3cSfFC0O+kCGCpOtu+xQhh5gzKVPPRUJ3aprqA8bFwTXQwLhtw3dE9ma
8dc/WKvrs7R7vPd2GTtsCVmFKw7G3Cv4U2DOGdahUIB3XUz5K+eqI/nct3BluJxz1fPAkiRX/Slp
h43AQEDekbuRFFqrhpSVk6sLjGtuvIDzmEANt9zORhwHotliTlLk2OcpT8XTaKsxR186LqGjvqH6
9yBuGYP8cFjaEF6woTyVL9TXYKWSRLC9Erep3p2V2XUNDWxp32DkIHBf1vlO+niPV4lE1hWn5GUM
z7b3TBz9mzBpA/sPy51y2bs/0JHIjVm9r50zbM2oEc9d+hD/lnQIZQ5fvTc28ZVEVU9mJmyvs7e7
g21ymLyv1HRjLB90m2Nu384EYuZHdDIWyYZjXLsOWUFUuVgaM/EpdgZiM+pW2Ia+bblB2Ydl7cG9
bqWen6ZFk7rD/EARn2XzHOyGRX3yXDWgemaAEhg3WpjgRMS1GNRIVhxwq/1OhKRS6DIU8zjCWUNE
UuukNQlqnHqnEMJSH04wOVuF8l522gddcs2gwyOjJtXw7wqT6eO9H0CfffjIylvl5GRydRn3MyQn
7/XdEwoPy4PrQUR2FXoc88MOky3oMFIkuSDQnbkztKIt54yNHDqbGUNztvNtfE0QPJftV3n2Gok+
BlvN+8xb12TZCWhp7HLQvhtjK7t1OxUhmJ/bD/PTE+tloHc2/Ug+e+66qfsIv1NE7L0Ri32AVzqi
bROYjZP5CjuBwlAdwHFTJOWacUlx7BP/551qiqwdvP3PwMR8x8xr+mwvjJ45sFr65pSaXqp+jJRw
K70n/G5gBvmhjmX8oCSy69AyBS0A8fsJeX9/7kVQ5pBsJZpAC/NeFfMGxGdmyso+wHX5LL5kGwOk
xSBEPYNoB/w0qqMJo0TiEmONDhkWQF45Qgzi1PthsHluAcy4Nv6yJJh7UD8EevfXSL7hOOEsQD8Q
ugeWJsxPUxjomq1BdJ9xmR5YMUyCmuzqMtcbBqzlpXwhB5dHDWgfFueNGQOwefRMe5lxERQccNBE
NU+j5PO/aetnnuW92Z6L9095CIEgz5ns45JBKIOuWftsxgFKih8WFIFry53PAUw3TlksaKEu+/tK
mq5hzmbv3wvVxb7aO+hpWRz9edJay0l7nxlBZThnOwhDXFWhtrIoz5dKyS5jeqb7y5yaYwBWwSWr
oCUxrTwmbwlDddESYUn6X6H11m5UwSB2ckBo5idegvyreWBoGPi55Fjsl7QnDjyzk5UN/H1lGe1J
z34jZSwGqK/mPmKlJBcMLD+dLgz4mj4rJRAwfuzBJA1Sv+9EkOrX4+n4cWnnINmeiRv/VgGwankX
Uk9rMy16jKGSvW/bn5vVzxCYDIBAUjTVdqg2eHsuhFSo2hjJdjnUtzAm+IM5gio8dCyBhax9P3ot
bhrhqgF19KY5P+DM+aOZf/voFOrcI5uDj/D0Ij75k0Ix4vae8QG5RTlTIwyc2Tq4ktE/lRPS7Stn
2Z7833lMwkbVzZ0InkpVt9osCTNTw+CMWlXkJCL4trd7lql9LY/nyoyrqSrGsxJA/XkF6IpGv2EI
8n9sGz/NyFdQY5H866DpUPeR+unOOf6AL73bpWKGMrW0onU7qf2KiDxpVcPW70GBwkLAF3DpCqDz
FNoGUsaPq3Ocfcz0ULIJ7d+Da16SGAnLuEjd8FLvcEXlqKd6WskszO6UihqSc4t3iJzNCzDA+5cR
qZGh81RoDP5pe5TJh35cYKH3a2HfjctusuonnLHA8Ega1jjG4vCXyLbeL1Zx3bWyBxkf59+XLt9c
jKv94eU8rlzkudovn3NsRgF82Y901zKCHteLJWcObMdzs0rHUPD/+ALEOVsKlIMku09hV1pLrf/5
TJHKVFz8s7lGANQq/j9AaSLxIg22P2Xu5bxG4ErdQt7rsXjcpnZ4HyrlEmItB0xcHpGCD0yet47S
mOpYXd1/0yX7tlfXdXc9YydHbcoffQD9bWM2aKOar2skJTbqqrrVVdmKDokn0OwxevpZRe3b5wYv
UCqQs1JvKohKKp2w7p6XeeU7SFq80RDO1IuDtt4YlUogel3uxQlya4SG2Cc8hpEeDaT1JIZJP80c
P5e6BFsjDr6mNTY8LLaGY5srUKV3VbcuBl+Xtv+5zfHZ2++XOJ2bgDhVppFMSwVuE7hZRcy9W++E
B9oAzP/RNpgg3j/24ju4ajmPyLpLtYzz8vmGWTybdFyzHMXlOIOnxc5An5kBgqrPf5fa5d/M728+
62J9FgscNLWG54WddyWpPfE/U9zpgfkDk2v2s6Of8/dszX6QtS+yC8ZbjoJvLNgqRHxcBrnEXllD
VdHWSsat9LoNweUNrmrZAE7BueeGhB4rtM4VLwasPEArSAOfoTN+7K6gzX+c3VFyNcnByo8W+aag
pJvKRfKMAaVpDO8rl8mNOC1elmEDw/Gm8PdgsNBjumQN+vk2iFK/BSfth8cKfa/bM/SRYG95BpSu
5eUQ+9UA5y0DATcqyt+250mFYhRK1Yt3DpSHhLhBTNmUb0XAoUiWl7aTQ959EYvANZB+sb/8VOxe
dxDm+4jCVOqa7eOjODenJXQ15pZ3Ak++ucOkaQiBouvo6E1E+oCeRWjKQMdH0PY6SUx6fOtnKcEu
CNLImGT3Vc6VGAKysXac65W+HWNS0q1n90xjj1MD16SEJnCgdsN6ZbDqNZqEBchEkqFl/nZUxkfR
yIeMXjObKoneFNYr7kNJ/hl86aXkpJz6Q7ytsRgEG+0XmUXdgK6TxD5rwJgvAS8xrDa2+DZTHDES
ejdTSYCoKwK/AD/sqk1m47HJwcu/Brel+/sksKWuZmzqK316uSVyRMVVOTPK8UTooF9gBILZ/aq+
l6Mjmhcd3kKxCN52Ggg1vfJkuAwbpfymDhV2ueyOZ1y1vKlzbTXJQzeppSPqEiRCN4sc8DYQSmqM
H0AddRjY0ZshI74CgWpEd5Eych/X3A+eulq8jWDRf+R31GUV5uK/fY5ClFGTWEBbq+Gr7aL1Dl0U
lkfWkHUB3u2D2nkf+mI/pL1500oC8EXLYUJ7Ql8RsXezioVwwK0977rDnTddYLp4y8la6Roa0zv8
moxz0hhJQjyp2sDDGC85iImJFiMJHeMsHAZ33/aKKLVSOol5X2K06d9lfaudtTEtxGMNKmqNUsUG
sHPhYhawig4EYx+n+mk0ZFK9d9Dk7vB9DFnspKrnmpGQPey+/Xw6MUJJ8z1jys8aHNg+Hq7SLsnS
RlXqrtzmNwJbFb+EPiSgMfeyiHUtjw+jAHBMrR9MoyrdQc1DTRK0HnRyqLTTsC2TqTqVMM8OST+X
4082rbkReIYDNcGKsf09KBlvq3U6r1YF3ds7RMjcY+iGI9551rrtQ0ddJ5eXDRTSXEr37V0b4CAH
K3aE/5RMwOwEOGZhzOqkBhSQb9oTUxBvWUldqurIQ6fKnoCEPOhBumhCk0xG9tQ0yUPburQeQmvZ
Dwguddvp9H5OakOYBa+Cs0Eb6lBACtIIFpFoRZrh/yW7Je0kSkGUHyW3wzSMxaAIbM8ToD2C4iGf
HjMrRE2SHBYVOkwbhvq/U5Gd1x50Kf8PbgOXByLIyE2y18l+llprLBrcBcn3J6Ube4NLkKPmxcc1
4HTqoTOxDRwfGAexFZZx54R0fVP8OtEufyT38sCdkUtycCehajO8XIcvpJGlPw6CG9X2ktu71qy3
H21oibbKHUjv0IVkixYGUlM/KBdbyc+ZeMwPafBnx1egnBxayN1ZMmi7uOiEAtLI5FM9aXgGgR4s
5h56HzD7g1BCZZEK6McnO3CMaOX7Z/ENsD3JTCXQ2xuLvYakkroOkLSr9wtBkLxPUyobtHGSu4H2
7Bk+w7QL5KCtJ26Kz4Rz9BlRHT3LHVfPS6JyPxtuwGsXOS8gB+C3j8SFQ4ses+y5h4CXkc5KbTJS
XhLOesTDuCKxpoSIt5ZSrxJpXMOdpsjXoFnbkU4Ja7o8N1Oqs0c6yAe1jzNunHJ7vpCv/e5hnZXu
RhuSDXx5TWf3nnwaB/CaS3xaMuQ37v2QXPjh4xOQDdv0VD1zYXZb9BKgeIM/4qIVt1yB1aHQmXKs
GO1dlhZIMxCk1JRkD6BrpVxtegk5q+VGX2cAQqkb2LvPPpHPTj1mxqDrwesNm1UOGHAgP0fxdlVG
Vf4lNJZSFYZ9QGKtqIquJFb/M4R/ohVxOH0rUt4JAKH9RnHqADS9qKp6hrE8KZboqchdHecqMp1P
2EJBDzlLhfNQqO3IiYMBhe9zlOFyHtC/4SvKiGZJ9YLF3cYd49Lum8h1z7sqfx0lQN8eLSN4Z5Q6
V5EwXmAs5xISdclJghxKKMEmyvMQQRQEUv00NfJDLNYn/iduZLNlKbPU9llbRomMRmqcFOBJmI49
oR+FvvARmo3dpSkM00qvEYCs89xRozCuxMeNgqAMsxSh02YQlVU8LP8URpxpzPw2JLMtZDl0fE9h
PBGNsq4MMJMR9lY+8X8nxKyWJMH86lDpXVq7+euhSnTR/oRnoynxudNY1pByO4400U7VLMuw7OCf
3SqJDSW7B9qtRlmdVWUAEe+orsLUSW1vlqibCaSyQ48mMTtHTiNzNI8hcYbiVKQOqRiNHiQuDv2x
QCK7T9RCZkvKAzQxWagjhQFwzUJkgzi0EiY1kshU6m3zJI8mqgbqWnj03ZypRmdt7J3mODQkVI1t
Q9ie+lz0jbvYHmTAFyINEyuDYDbNWlGYkCmlSacrtl+//VcoTQb0BozVue9eQMta3vbw8RmbkiKN
Lamzg/9lNNtGZDhVPV97ywLYW1hZoAes+kPP8AtLM4QEfAEsw8qygoW8sLeFIDYSyj9ihL8AUI90
VAtujSY4pjZaRLgQSxYm6tkn9JMIHkCi5YX73UiaSWAmC7QMaOwl5ljZR3dA3rdDUuLpTeXY1X+9
qlnOsm5vsxARucrhZvDggGi5SkUerx4up7a3Vm/t8t2llUuDOct+VXTTQNJHvqIbIZShG6tpO+Oe
w1k7D/HL/TQ1HazDwTAwhCE/NLw8C7KUjwLKBzNLhXC4q2Urny+UEy2b26Ny/UpCpEUWFbvN0OVG
/LoyX0+1njTCsvxjS5U7t7cbyRPwxlNxe3OCGsQ5dQ3MQskp9OPsUrR09IkGgQkUi4mZCyoWY5op
uI/xdYdOvyiO4Nx+OmoOj5FaydBdLKBGxR+mPxwC2IwRxY4lDLX4ux0Nx26AWOvr5HPoby42S3CU
A+QguM2SD+6bIyGAXBajZJzf1wLzbTSlPV40Bq39uGSjtYcecNOFH25qdnQkC1UZTtplKIkuNBoR
J+ALIWenkOlo8qZTngwkFrKS14srsKNwHWHqurIblG4FfcizeKb2zNyqYsWcg4NaqtxtJXflLryq
lUXD0PWKt9cE5R3SqSHCj8G23XwDbOhyD9ePqC0oCUE4ZHHjlHioYWixUsLPFHYC/pN90N93qDD3
dm486xdWFGHzlNwzCx3sorvDSWb6qYI3V2UaK7UJ7Ugz7r06/ktT4BkWWbt+//9SN/C3p+AIDaXo
r4Bk5FLe0+d0+Lj1tg7aWosRPLsZrYCZdDEjgEXScgbWZyttnAVLRejunW2x6lUH4OlQDEG5esZv
+p6py+tSSy5XhiWpas98b1uBweI/83+C0JoNZxRJuAIUV8B7bPzxBXHURQZrrKjzeGNGTicV1//M
qLVJ6+X4AH8FlkqEgJ7GPVsNlYJrEPNQULtU2KbHe9y0jgKL13ZtpSikqNpxG88E1BU8acCQSx0l
6JROyRB8SrPNkSyRS38s5iQmqgcThua6G+TRkI4ueQP8QldRcDVnFhv7ox6eE3bgzX1bjv3ggGc8
eaRghzHu9LD76UeEwdmfUs59UqJD2lZwTMB/ODrbSJcWJdixpPs8tkJXd+1LAttRIa11nI046Fd5
1tGJqUFdXdqLny8nyGVeJSJKQ0AZEkMhEKcgMuUwnScupZ0M7MCg4wEAQBGwO3GEce+MGS+Zh6bf
i4jLCnaQTvhQChg3N1cVprmFy0UOf6LoitKFOEVO6P3idoPm3uE5fdK3Oc9Jn17TyPPbIsA8kbEu
lZjfV25JMXOlS4wRACmd4rr2lxuQJY7FxghX2bHpf6ZKPKVdr6ysDl2Z9IDsM28yo0HMfS+RFNvr
jW2WmwX0eBLz01S71UYp1NA1709GJHInEes0cEb26p+KXZ5BkIjuDPUI6sW5Sw7wZ/KiGPmcijVr
iGwUsHUX9Zswo9+oqMD5B05xLiurv+NXmmvy9ACcxMzHzYpoBfVUW6BUB1nL2Mgm96Vsq3bh0vIS
rOy8ZPiuQHZ/ChtkdEzzeJ3BpzfuCRuqrlHko2BRd+21BAr8DG74e7aIzpRFUy/XcrL7l2krb8RF
IyNWf/JiCaGW/rqxLLKcqJylW8Qubnzoxcm87dRaJQasfwrqcYG+wgQIZbgf5fwjj8p9uwBktPlj
qdMVtxSlMCfeJ/OQFSw7tkcITT565EfWGqo9yzuRwVVONtf6mirxE3ijbyCRcUE1M+86L20PymFa
DGMz13iwmFnpfprBnorrkj0XkENeBfibV4WaeNE9EqJZK6ETwb+DAvi692P3NLYK+0LK9KmFSD93
WyVGI5b0db06F3MNXeJJN2bYZPQR7RoZBUyf30UsjFZ/6YdOhd4dRJTBtiNqqkjoxINhn0OgMrU1
AhZsYY9jvS3ELGZDpJcW18thFtbxUgstCP+bx+0z1AOojyXlIYSTl5QXcB0oWxdtglYx2KCnruG3
FxdUgH7hj9hWRPYtB+seAXJpsMFljJxICZR+iN9hyG2X9Qw5fWJh1Lfp7XimByRBSJHOZBXcOOxK
ZbMQUMmkN0LKYxy6nRppzoFgKWeKzpxYEg7e20XTYSPDByko8W7bGqBFCEg4uMXoqk1I6opD4CC8
FlhJHUbqSeWIukRitc4eeT5AHkI5wIUn/P6fMO+7Qnp6eFcEqQsH2kcYuZzXNNOp4K9+JR/HkhxC
7tW+fXFVcR+a04zGIXLGF5ZXWtlThcAhEjPRZKB6Aq64kaXahLXVTG2tCPPDmpNos/23/Cnc4n5p
FupKbwqGtQFH5lPuCEHuNBxM49t5iantYW3yxnEXh4b+z+9UtWHeA/nSGpXs72uambGYP5UazNLu
3tbCgyERo24J1fLVl3pwGUojg8NuMrY1wFTjpyp1H1Xsml9ZPGonZQ3e1fc+sNhhnc3NGoD0p2Bq
9cQVLFDbT65y8Nv2LoeAST82G3dwgTSKmgF5neU9rmXpPoa9hA3PzTKmxLAa1ErVTeBugbWiDmVY
KfnPnn1PMpUu39Yv3k0NQmpM89PmTLlkGznESLWr+aM9CsJ4UObZCgz6oI0FgY+iRyqXbV3a9kdy
naG4qcf+AlsAbq0y6Kd+UiCb4qAc4/pCFGz9vejAhfVz31HOg9AOLG3/a7VnTsnFQLUpmfWblyz8
oShxgAoNWfRgyA/XajeYYpCRf3OxggSx3nBKedPmN1jjdcpqsN/znvU+MLCaYEMmjp2k61L8cthi
1zoaRLGvs6lbJXKL6WRB7eAKFXwi1ZIFWU3LbvEyRIbT9T9zUWR4dyK82FVN+GzFA5qgdYJBZiby
4MQT5fV0KQ7A6X18/7CaiZriODyK8fZLr7g7yK8eX8M/jOx6eDbEbDZr2tYiKKrbORBYk3ylcCz6
vFTECh3+HOl8IzKi+kAo4QS3NuLb9fZGcXJqAbKXGVpNa/5+7kPZcR7KDM5MPy5tCzADntSpUPIU
EItIfCCD20cv/W4U9cbmTe6ZQ56NeDlYBYBtBPPyTCQMZFxTgiBJmkVZulVtxWjTC6z9nGCnXdWd
tDQYvBWPvg2QbzIyzvW3DbfIAfrfpU3imM9RGZHLhw4FpK+Cy7k/NW2GoV7Q2durMYXDKN24MFEZ
7ec/it5HrMHg216PAIYhOU5o0VNe9BV3GtB2Vb/Fy/prHIOYR6NywyOoypb/137uDXDiAnxKTWWJ
na1UDlAfVRXw2bsLazl1mG+7AwjcnsT99xYC0pId5DC0dI/KdUEwJ+kuLOu293FZRZRXoiafbLw/
a3ZT6byzycCjZMUBJxAjGqcuUCm4KS4XSphiCAdmNBXdp3t4LId2bhAlii9gph9OzUPd9S4dpoXn
Ipg9OX/P/izcQNQRB+hviKzXx2qPyTj7yEHjT8tzWxYnVPT0ImNp9K++F3wFkxhZRITZe+r4hn5W
kKvCfceiu4ia780MhMEbEyMdROCL8aWlsO6RbCtSaiVTJZpzhWym75VO03uAYbbnLQwfat9BuaOl
rCEVyrvyEz3Rm3DWeiSmp7K3q94i1aZy0xWEhwRSJDGhws9LjubVEN+N5W1WLkdSoIrqDg180zpD
FiQoBt/sZc7+GLKoXsYFwDUOx+54jvTJI4+BA/YhPsUtsqQ1+o+wZ2MTv4zshJoGfdffuyfXodtX
4X50sI+Vd3RAJyky4yVtEdUvgSwcsHr2ylXy1tSIfsrJrjG19YWXWpBzdcedQSDKZU4dxy7JobUU
AfRkjK7P4QkEGNHOEdu4roM0lcvKrB5LnHZGOpVc++FmPGrYnSsEW+GPRitbGC/xarYS3WUbgZ/s
+DY3OZIPu04Z38pnAJ1ZEn2u6RibDkJLjTKHQ412mfDj0g6rHxEZNwdWSYaz9TuaiFwKk9YvV4GZ
2DHQ+P/kufzL5j1cihmY85iGIthugIxbfnEeeesUnuOewYvtVrK49918tZOKbear3M9KjmTgYxQN
6G3lJKols9m2P4sXehHI3LaFAH0oaZ79fhW9jpIz+pTfVFAbOmUPJpNRuNAs21WaDfMZZtP+SSzM
gqDQBL7SJtJVBuwVF2IwG2JPTCEMlNj81hUVRhquEY0VdRrITXTRpRqdYTgdyEqW0yeB7F6TJSN7
LJ1DDw3oadoE8BrdsmOClgU2KylW88A9TnWSAnJ57oxD/xy8yL49guVhNvAXIBknc+Ey/PzvK8p1
LDljoAeK9NuQZ/Ea4C4InUVABvsokUn8fV5D/tecc9N3XBedOasEbMtsV+h7QmJhxSqTi1aga7/J
U7AacEiGja07z28bR4+HtxDSWGZvTb63uEwSaqbKFO0JHA0RC0caePhkE9h71uYD9BntXakha7nl
E/TxdoEKsaNSgwht+nL9Abb4dfXmoZjrZ7g++3jyQ6f0JhMQhR6/s6z2Jlptw1DMQ2NiGZgOQU04
jgkItbfu9jRJz9V73vfswa8ehgAag5BIGSmzFT50/xeNE4kbNG2iLSx682ikt/at0hBAAU60bfgg
3q/Mp56SRufsTOxUKxWXRucos7xv+rPWrRAGyqcqkHUp/m0M/m+z947fGDynuDcdYbTdRHZ5Jovp
IkSHws5pR2WgjtCmfqZmckp/qYMGm0AISiidTj0WkGP8hHndzPaW8oXMCSY1wLrJjrmls7tag7xj
Z2NVbTVK0uHzleZBEJi13A9Z4WSabys2xL+LR1F8YN2DEYchTbU2u4ZcsQWzj2pO8wwdIB+zI3BB
q7wPKOwJGRWNTxwBB6GYQppMGgerBNM4saS88JxH1W2GJagDZHJ8ugn+g8BE4hmr3hdyzzczT2NE
rhehNt//VRrej1GGl5rMCPK7hJ4fk9Dp47nM4dd2Zd8yhQyT4sYJuGdyftojwBbET93Qr2w8qnKN
9U8ZtOu/WUtpkfNKxcrS32rCm39hnWZMhm4Ip/Ros6UmD2XkcAfqcNowpliauv17OpWl36cNQz/c
vFMtKQ1URuWcFbfnbCvmhUJGvcuVLFph2H29tW6yKjBXvqOtb7Zay8Jv3DXKJa4lAknI9rRDErrw
tGI/WuMMHgjLzV+WL0LFH9rH9HVxPrIp2VqEge6R3NbUUuyxxLFcK/u2nDwkqgsV9POkY3U3tIea
Fr73cnm/oUPgWMvBK82KtgxlBsKzfzU/hIndj6rWEimuWfYOQ5rQVNKlK+n4OgmL9meFErMqZ79I
uIF+C9vGVyuys+BIRkVlifTRltHBW9wL8+qPIA5Las16uq8zobswEwUfwXDTojChk3053Fjr369u
PbXEmSiTPpwJkDMhfdtlFXIZtRybTvvHPs2477rTJQv83M68e70srDT12nFpeBU5Kfw4UlvooCY2
zMWAE8w86+fHC4EmXz8xIXl1hr0JotXVvs2QFdeNvqfiv6XwRYHypdy4czywdM/1VIAq89HxqXd0
bK0IStEgOtqWRyD/ilTMvHaAcdDqDsEIJKLVO9UOSpWXfO08quroXik38QNlTU38Jx42rC6s4dDQ
MK18Mx4mnxgfPxHVCfhc5LjVn8lQFPqTx9Kb3TOdQ50PbL9Ri098v53mU541cZL0tVpYd1WOJCMx
aRXFPJJE9EaMkx3pQvGN58chJI539saPH3HyFpVVcwE6muTuqud3pXTNfjmqcxVk9Y9Br0dEgVO4
H5OOVQXNMfK+nj/kEQYg8GbvXCxjoiAAnpMQ5w9nZu0zVB687JBbKYSUuQj4jSwteWKEQPbiw2wF
GnpKp1hDDAgOl5bKLOEK3cfMqjUscxly7pR+7h6Oe3H+fv51KvoAINIeNCjHLxWwrNJgd1ve1ax+
3zTzqPa1Rk8E0jFo3jXcxIk5rEY9j60RYcFfjWylRqs83ENY5kHKABzpP7gkq/ozgPcPfz1M+Juu
ZW1vmsW+W0jGsR9CedPuH9ZJMe2XK/I0iYF2eoGrmtm+CLLZnXyhOsd1pI+3FmO8n1JMH+L2dMn/
F/fS6GgawAa9QOi/59DWNfa3Ar9hWj5lZYnn2r62OZEOADWXJ5e0311jGIteqTePOzRZMow+SI0C
KaO4LD46PT4IdJda91N4HzQNBADsI2ffxLxpObnXYTlovB0oK5t1NIzY7PlAsjBF2gmadf/oKV0O
k8CDiaIknm9XjDMJSm7xE7VbXtbOX0qsnw7cju7nVzOUfXaFrCjDw9TGkslzCJqgrHdSPBCVlZJS
GzhfJbZj/ndODEU8uSSpHrvOTCTnknEXwVKwJ5cHn5D/9kiLLxZg28buq9Wl+MjAVew3BCMRK7p4
f19iqnvabBPLmUMnYAE1KpqKcoW6lTkP2D/7SZXQ38znS5EfehVe8XJeepmJc0hPibOK/KH0aLfx
hz9zWCQ/pS6JiwYpOHSxt5ZRt+ntqNgqLb+qp4PUD2rfUP6xs36KNqyMcKxWJAonwlyH5eZadg9H
pS7jiFOeuReUSyfiZGV7OJbWy4H0+pr5rCpWBItzxtxz/c9wo9BzbB4inMrDhRANq3HKMmVWDoaX
Z5xhlsBT8o0hvW4WCGqZzXnwjHCuHM4QqozafCTLHCsZVKOglQfORT9Xv88WRH7UJxOvaPGfZoTf
W+g2BPHEc2tdz0NF/EvNnsmhf8Tf8UeNm6VwveYq+/z4PnLxbOKPeX3OfJKGoVEKDrAp6NP2TOPh
XDGurVvO/yl0gy2rcaZcj5i3UFb7Y8YBW2TSWk1funykzUnSGFFUuekAQ4NveNAgRRccPdJpV44v
Uo/xpK0wp1Ysr32/VYvZR/fSjiOLT4wxtRv4xjB1FqXzu/4a8j+779Je2tRpqsJzMs37ESc3g6jh
VLTnglzellpZelQh86EN4hRBe2CySKJG0NXf4oppzXdcK0PBtiMSeHFhr6Ury73UQzopZ9eyOrFc
vd6hD39YrRcMgv3kDjhU5gFMXbeA/Bu4TkMeESzwcd7iNfbvt/zVJE84zhGdZxHEudWARi9nHdwV
zvkKtTvYbhScN43M14bbZndMeJhx54UK0zAM0cs1LWXhNteoazR3zWKjvpmBDeoQ1cVUqEKeiIqH
OsIzcA6Tq2701l6EVWrB/g9rABm9f1nbgvG0ufB2b5L8up++6dmvrMm9GPc0UAXXCwiyjZdPzhwJ
kD7y8rR6A8YuUki55BkkTdvqSNd2DRIgkmfyL008+/lMTacxbssGQJgf7HDfpaFGVjjBflRzviDX
BpQ5KL46fJ/3138/GRV9Ob8HZgWH0Kn/TJM/B5L46eOX5Rq0jWhLe58Z3blcyniVOz8oiyMReeTi
ucxZTROEIQLcPjSrrcVGe/9ZTE83Fx1SV3rLtdPCqEo8veMSsaVgI1G5+YEH13+E1zvdRgs8BTyO
IQb/D62s8DZCng6h/3o8qGIbtfVJ0z7KZq/RRmQo2M8sWbRGREZGCMPxEJiU3+nZQqR9Z/oPT/hs
fAwazX9JnbZBwlF4ZJWwyDZR2rGiN84Hv1Ljbgycojs50+fDHC1qPcNLQ4R5VglUzcOPdv2GjPhD
IItAd/hPmu0iLnVzeZ0mDCDOLPdLMwPZioq30sm75jObVFVDTM1VMZE401el4b78sDf120bM2bfN
4sC8QIDvYgfjDfWo3ifd/WRz6aJWJZg69YRoio2UdFRdaZhsw7GOCha4cWFazVL0RJhDXtqya0xw
oCUdBk1V8KW1vGbzp3/cy1KyXmbG2+eV+3EWtJh3LQBYksCNmk66/KPpxq35JlexhpyXUYJfpQNf
E5SI9j8Vn2wAwDQmffq1k8C/iNZQsGVFCAIHQQAJC2/sXxIwapvy+ZBjcAQMskTZyNTl9JCFpRfH
tz5oiXkpEL9KVLUPqosnrDZPs3gWzdNlBBxHfbqyofmysbwbgb3+/mLTxyYvud31CXr30x6nt8CJ
JWqbzQ5BEQJuujKEvtwSp4jX5rVWuuKq4oc6u9fUMKshj04CuAczZQKcxpxGOi/RP29MFll/1VCx
5p3XQehNkmSHPd/ixCgWTnaFkBvYOEpTfhNU3bNjMBwS/65DNqrFcmfTo0J/T+4SNpkazH05c4f6
Nse5Adm/KAvpa/Ypx2fFgw4jP0+uDBiVT8Q11hLMCd2606U6/XomPNKdE/lNeC0W9Nxb06CH90EQ
opTOnnQ62VbeGtyHtzCFzh+bGDCYlAB0peirX6Nwne0Yi8jguM5mj8ceLVgiQfl47Z0PRPerZqoD
HTnr2OWiUF8ook2lRIniwMXq/cIvrO23UDP4WWnrVuW+8Adrnt18zvoLy3LihUS7HSaZyPzpvWxn
G/F/QlpcrfEwvEH7OsyZpsYrwjYEKVqTED0MtvCBemj1YCk/lGBcYxAZuZjn/fdMXgAmcdVeLDCN
y/RzJQufCj4OjsU0RLLRA5FDDSIWOfNIVDIPJRYoA9VfNBDox40/pwCJS79J+uWn5Cs9yCflaxB5
HAAhQLBcTpjJcUPmRhXvliPL5GwUJOANej5TYedBCUg9oDyXWBZHS6GZST50C96M8WLCWjJ0HNg5
kLtkAfbmd14eu1Q8l0pzLU6R916RRaukClvif1qPTBJpSoz8ukNynapCIgp1pW6i2Hv6+jBMb+q6
xeiJ9AeKwhklHTuTKkBn31aVzNYR81SGIVWYKVFn7YZYJ3WKYX3pD6TgzsluAAj4POqTcckLNvo6
xpX2EmsQkUiuHx6sDrlt48cvEci94ELKLXJxHMrgp7CRB/rZlGm9HLJ9kFodI4Ewq7XPm0O2Xxau
YiQ/2Q1ZkZc8Ev4XqU8neXGCUuGSJahe+ChPj4C3FQLDTRVDgVMHOoTRB1pAY/fq543zDLnvRytO
RmQnQBnnkvA8i0BAMJvyvf9RR+zDSiKOmARRTlq5ZU3Ps1oWVdK0D77cHqKVdxJUZEremYAW5Rld
qHP1qB+u0OgugcmPwr9XlfLrouuSkjsG+XGEKYLJB2t9SpsPgm3AiMT4stjCYng6WXL/dKbsu5aF
ShjgUI9rRNVfq1tzT+uaB4IALhVRHgqxWUKx9Hyw71X1cTzumiO5zHRgZPDjX2r4rq/DR58tXItt
E9u1R50oHrqGpipTFefcCv+wVV8BX0eJIqdIOwytb6UEgdT/SVh3c8Tih1qd46EWqc5ExDYGzqYd
5FXtdN/QNOcnOh8mK2YrhqzXUf6ElvoZ7V7XPjFASHhGY9Y6JU2CSZuFs+Vd7m7CRrhXUJ9p7ZkR
7qCtStYAkMvGoDOv7P68RR2pwX3LFDOMXv15YBwnbqCV0TSObOhE8SnO52KvOAalyCeoWEBHWPdJ
avUtbmokzDTtNEgrQaOSQDltIstL5KzMXSD3uJBweDv4SKuwD/3Fge5Az+w0ML1TPA+DrDfoZhBy
s4WuGaZOwxq+i7JbyBwEdy4RYoLQUe5eO5cWuiEKbai2LmDEmgm98ZRUhT/n2jJhDTtCvwja4lY7
OPYhXNYzvstWDPNwQGmBxgTC+DQ6cfPDe6yyMcztepSpBmllrDX/atE5ZuO8u2Wvk6KqfQVzb+xe
0fNRpTwdYWUdByjy6ml3p4mOAX5Jp9QuWEKR9qC4s6I10eHkNiBfgr2OqWzGT89XLr5vhp/JQX+4
Kpx3ZM+dAn4GBUUHPp+7vMSa50zoW3zcvg8vRoWU6AggSSio5su2rXOw/EHflwJR06H3eyQYnHoL
HL+juT9wuQ7oJUyy/dWdhpBYWjDe1akD51AqOyTA2HEFmvVmeapbKpWfsDDZ7/I3fNqTEMVlKRXI
Vw73aJJPnSkAYLnwS56Fw8UjSNzms4XB6r2MVCTiCy+H4e0h/f13EWFD0afDbU7SxOdhMFNSzvVC
2EyeoCXhbOnSumA0e64kzlD1tQOOZmOEIwKe93H2rSPMWb9vUnZ/uGT2zcAfBjLyYeCE5+fq5kPw
6+lDlnmmh3DaXEwgahNusW26PuNtqoN/fh7x2nz3sPNWfuF/lPSc5Qlpj4vLNBJ3HcaPjMgNC6kQ
on7mMKkOWUhVxFXUjHxGGlR/YyZxdODLSYVHMd6SiMv2rg6CWLsXfVZgInUzPJU5WnDAWJd96Cit
tQev+OFQITWrdJTF1C0kuPjgFDxXR8xwzUTm9OPZr8w/iiI3nl6ALnYCdaOD8enPvGSD7oeOzMKl
CcQkzhFGP8ejnlhSdj+odY+DmGeLw/P+rYsNtk8PSELf9p2FOnmpVJoIQqFS3jO6u6l/n01ENBlP
BLqM+poX4K47gaKVJK3SWezLRE4ufDM+2JNgIkfU1iLW0ypxi6nymU+ndiTDM1ljM/VUQOwSj3D0
DkvLDizC0uSgUOJt7Txt7vNVLFcftlEHVrnkO0DpiPnmmjLHnujbJc8BusS24s0JLtx1OTh73jM5
FoRoWOOT07YiV045S28KJ3XyDRQKLC66PbELrfnVT/WijHvu+b6lFQBibEDQnX908V7Js59Qd9WZ
Fo5x6trZ6zPiKQvMdg8TxSHMTc7QCoKFUS4tGqAx54d16ThPDRgq/JZhb3lNCDniGxAUs+IpWwNM
uST/Wfs9ZMq5lCSpSIU4QVqrn990Y+57z0eVJ6jvYytUWiLHV0Kh8Wf4rl7yKpnPkm1dX+/1cXXr
gNF0O8LP0syr/q6veRLK+CimAkbAdhqns+2R5Rj/id8ia9ViiG8efzPaOax0oSMpVw1Ktnaa97tC
fi2LQOtS+7+epxbGz0Ch0xymyUpiPB6NEBgVbDiUWfeAPZip1+vZF0Nc5Siqd3H+8iLqDcanT9kn
Z8eBZAH5BVI0T/63nzkDyJtEcCXXc01baNTAZM+wodZBrbjPujD5P0kDuX38bbvZ9xw7qkbSEi4H
vncYPAkQxLwvX2EdgxCwf84FVfmyZomvaIWM09LpAZJWAERrnx0jbfWTkf6Y3GEkvmcdq2dLUKTG
P2fYQ/AbWLQ6e4izKUah0tzI/QTnRp/FWpLVYIB5E3cnhE7bnk5lDo6QAM1PGuIy0P0QF9g5XRxs
M63aAl1BWlj8aRGfmDm6XZbuI2F3kRG25kxyUPjGATz3hXH2ODNP6TQpPmRxvbHxiZVkg0ZothHU
ZyaECYzzSfM7/2baXDIGPD0+KaKz3P1lX88/tumeIyYmzvffQYeycWSm5qUzx3Ra1LLSkOzyewhM
KqdgPygypcAa41VwXnN3QyKwtIBvuRVGiLbGjXN+B113K6O5p1uDMf5+oA1jHRRKoOKP4N/lySaa
znVEXEKpcbVcIum0pXnF3IADHJfWaBXIhy6MAR/8EBDQ7Z8b+Mn/LSgi8Q21uYSaLtKGEGtywYYx
wpWpghzv6DJfFJ7Rjsx5INToR6xKmmGVLyPE7BbRvCfScaew3acRnXXC/41z2Wh4RD/gPl141NwR
8CTVKVVJWtPnsqQDKZlAsAInx2zyqFbwCdHiNbavV+tA+/wAfV14ZZaDetis4Igo0oc7YS7gPyCe
5kDBBYIhwBDGVY+qg5IN4JTbiEkDcorT8sVco3YibWwFCKndDaCY9wgCSDTO5l9tkbT/Eb3QOS2b
8bWHyIjb2c4XYSFIrS4EOokSw3yOJhLy/aibxuZ0PWm+xHS8S7YK3mYlULlo+IvI2q71/QMcsgwh
5FR3KnAuhyv4YD11Zm8atH6FgbajeqUy0ovKQLXw8wb7rs3bRmMT5+rHjWedkf2FV9XMz8iqzalM
+q6pHoc2N+/H8ZlCWcINdRBF+25r6dmMwQJzrN5xYNUdVcqbjr8dnTo2gJcmZXdihe+88QxcdJoY
lVZKQSW3YzVEYeY2V3i6phMMYkPOZBSXEHcx/k6aW40LCfytpWQcC5jcqozO6G+8wJI6ALLnlAA7
ov4GwPyqV9Y+J7W0qOf3nu3vuwJgprNoEOHspXv5GK55Igy4K7DB4FB7R8wa7dj5AOsfqvmPCror
4/b1ugT+3ml0Em9osi6pjW6GSrBSh9IgbqTiz9NTRZH6H4FpyUSeRnqXbREhR+NQLzAaY2vWL75R
MiyIZq5ltGqf0bxD+5jPY0vTkzRcN0DjoGvS9MTGwUzcjSxTLHfZzidXu2rtphPDLENZCPtDxx31
XF5nVoMXRxI8Q+WSEy/cszVykUOarlIuAzb4fXwoYZm2yq0wuA8cnnJ+V1UAKwluEtc6KNDC1pnX
wMb/8S4OM0x/ibX9/2RApOOE2pBjJ5Sko1w+M8oSnDbx9hcfA7z2Nk4sscye92HFV1Ohup+t0DWy
XUHohLV86YiMfPfaTJ3j+EmcdoCOKFAbq0Gr/QKPi8twuZyUEWAbizvItjV57uNxgEFJ+Pc0oO7s
BgHrZfy6tRsB56l3ve0CXj0PNWola35foIdaYLJVcnhzm0WB7C5HfZSSei5Av7LqBVcYYJPdbMeE
Kg1KnNDWrmPMComB2cSNPy51ZmA1NVApkLu5+hvcLBl+g7qoDekVYIOpK4nN7G7wTu+W/rUWROrq
no8n6nKBD/SKjFymfxLMPTVpFJI1mYmdOqc7kGDGBpMYSTXNxHKoAuqDebPt1RGKRQZSJpr7+xTH
wqCC+cYs3DwBcmSKA0kvDoCp2H6ysKHe/6wtrK4ZyQEDJucx91NFmDLJDASNLwWGV7xF1i7VqBgF
eVU0SE1LvmWn4V1ONIrr3qkP2r0Rje8u2cjMqnvrnrimTmgFMmdWTvxsNprgfNWw0w0smahjoEzf
QK70efPClxtQ4NPkJEkImi40eJTDZGgzgyKWEfie6on/1rdSc9RoIxS9RSp5s7znaKyueuHOlMrw
8blLXaIVJ/gMbXVB6hCqMYR5hlBCtHhNyx9tzAjUpbx1E+MhksXkiBnncsMCJ4g/nQILIOSsp4YP
hWsULkmUTEKhx9diSw1NoGTwDrKQJsiwde0pUVwCB+d8zbb8p2CUtVjXCLKSKVnDghE7Eme1T9vF
7naMkagmssQGpkkf3ytorBS2bBrCYSYk3C3WYEHUJyJ7613Z/dtJ2gh5/S9h/sUD4OeldoZiNhTr
R3jVy+OXZtIzHcg9MXJWFL8VBc1X1I1xpCC7+uzr7n7j8AhKS1X1LWtN2fb7CA0IKSP9I4Qx/8K9
5gCro0fAml7FEQPxy4fY/e47Z5OFUE6AXsgtYGsIpjN+CTndESILb3Nkc0vck2RkjE3wYzfLmFpP
uAJsIX8ssN50PM8d605YIINkYWIbTbZhUf1hJd5p6Rbs2yyAgyQ42fChT3j1dxTlKE5uEGXLq0wq
aKTU3Mo9hLOuTrmMQa+vCAT2EnZ+ngQ9LB/1HR8Y0Ta/jtUKr4xSBNq0h5zxia0rwc2/4BHuW3x6
V1L0fyr/QubqhhmrUoMAt+NkpjzESX+L/qgNlFHCInL6o+mFXB/OzScSA86c6ZLXiAAi6OxiNYFA
D2XKXRgEiDf87keKU6PuucGys0BNfQD5cHo0EGdKtvnR62kPUcBez+QLYxyBzIIUnbKiFtWHzFEp
INTPP6hCRRd3PcY3P/O7dWGsDQLKrVMwtKL7ikX4qZXNAlDAWL1O9cgLQbfCwr1063nFb9VT/Uq6
0MnuXwv0nr5/nToBm1J2GqpDgDYaL57YhBvqENbkEbhAu7tmneAkTpvsVanF2kzGcGPFhu+vmaQp
YWEv4AZzFreOrdk7/oJIVTlpb3aGOyHeMFgQnKVgWJ7E8T3tXgkBO1oShYCvmZheG82vL6pdyDme
SFrRuy6yQIhnzCYTH73yZGk1H7Y9Z5TQ8gwIWZTKzRvhFoUbc6fIqaD+Ugm3fGG6o097UCqyNEgi
W+OpUFSC9dr3wGsiTDCQGEO2rIRZ+06mPvq5wgjQ8a9tC/2m8R9OfVx7phNUWWVjkg+Oh9Y7FAx4
3YVROrCrn9JAaRpGb6vIwt2WeO/81TAHT9TkohJc3vFCQ1Oouhn/mfIaePzVdbAn4UUni6bUln0i
h7oCM7UHPtWQGZ2vFsTrdj9B+fP08nBupadg14unsbcArT0fREA1ZGvQhMZTKENp1/ukq0vaaKRn
Yq6xLy9C/It8lL9FJKIad8+VKe2M34KmsudLWz3WE66Ey8Rt02/lDXagnjhnNLGDdbV3WXRl/EZe
bJwCkUXmk6VHV2XZoZYW4cGoQuLcvCUXy/HT8MN62mUujNHNtHASd2SQ9Vrnuto11pSwGmpmBZ5a
5VzbVQ2VFBSCmi5C0BkHtsXpRWILK6Y0zEGj2xWpYpQJdnivq/iM3L4tGOikgRVF8t5B/K5SthWh
WvGlG/Tkb3FXf1SUHS2iSpFWdCOQOwJbsFyz7z1BF/FgRnPTct6a+Ru33t5BUIjcucEuiwSi5of4
dE9ZtBjQCLbgaNXi3kFHvIVkl5OmQWUZmjIX3WNC48+oUUXEoMya12P9yJVb7k9Jf0QcGnmZHdFS
6hbnJuNrhnpdLc1gVHDTTXEY7XLG0dbqPobY9ww+8EfqdCPJZhnfFAlZlZk9Ma8aBwmG0KHPU4dJ
f4/oEyu8NLBLhanZV12MQwmYHSr/iwylu3IwFl761rtxAyXyU7vKS62yHfwjAjckTRMcyXQoHDGb
NWmmvsXjTDPqaiGJoJ5RG8XCMx/WVdMulE0EPkKRgEg0uRGtc8Qj53YUzDH34qVqt5/l51/Ukb8g
1KUePFZ56du8UT6VQoVF1athcf99onwdjKB5lfbvJzEpGXzSiItG+tZ78x5/RH3/VJk1nL79amtu
rY/7A1tmvpvNhgLI6vzkhfQ/1YFTY9taZbbNX+EvqM37wsJZVv/Sb3FgHV3MVDyqk6WV9AVphVRi
5q7vqhKBggss3K5m31XbILWKfirsmMCtC6fTnm1ODletMyaQ2KWXpNaqXpIo+q2bsxisfGMRr9vD
3hfnFQSfOgVvYcga4u3mZZ29YU+P6piW0ikNmCkn8Uq0K1Qga3tI2DUe4wYRSF9Mon/VWP6ecauJ
JRQUIUtyW8W8Pqsa/xVBkdnGyNYo75V3/ca75RdWIEpPEmqKA55NkXU+sNMTpYaksR+3doZDsuiD
hZragnFGsbobf1sQmrvTesHBwjSQn6L1qZTpafNX6ofeYBeBcPRc9e5mG/Bzb7yiD95aMgfJDcmi
Doz7bX2lJi0GSumMV3vpVtIkRmAG88VuJKBOZcaDp/74fVjwjzagg5745/UTeF6Nan1qoZR5gprk
HGXYQo0GVoKqYkCxvcCuhFnZitRqjM4YZbVIECnxKBxKqzYKFZL5ILOSQ4qOhXYchfe4mWMaz3na
qK/R7aazOz8FE3SBPJZSYHmp2+A7/df+hDcpIG03A0EpKA8j4XPwzb0kvf3yRFWt6B6b//2DmDz2
CHq8wif5evqsBLMyBr3+ii8yK0JYH9UdIUL235yGcC/UmRzFMWp6JxTG08Q84+B5rh2U5EZtosUe
AKqWrrcQ95lQ8vzSFtyzCJ1bR2pQeHmYJ87irnjjaU4adbBL/d3TEhlB/HV5ls96Y77RM1I+aIFC
2yJl29JQIuwm929S562QMOeO7cPfpVwVrPldhTbqMwUFrnTult64VBF4LAeRXKR2RqcJGRjaMMWl
jswQiT268TmWGOrzJ0BlYDk/41si/vI+qPsHPQwcs8asPfgm/AWoodwjtQQAkFDIzl7ggR1HGfby
9TQfHRUVnkvk+DrOxTNdPcRucgBAaSYrdnZ1PFD/qegbss6P3N541jPps1SHVfCFQNRCyRKcBkJj
M925cwfWRgoSDTZMBh/PoX+tFryjs+Txzwp6bDtF1o8Lfn2wpOf9BX0UTRXr/ZtnvTU6b6uBX8Bl
vFgy6pl+wO2mHX+eQlgpw5UvNNJdREIK7bPoSseSu5zPFXnG1H+H4RwIr7tWJKoXVoJLMnsm+yEw
ZkzVIhkLCmDVOKL246KUfrj3zmv+s+IzEvAXo093ZqHKvUYYFc/9kh7WdaIRPRDFcQKNdQ/G92r+
S7EAf+2mLP+u3Wyj5KaUz+PPt+aDpSriu67+LW5dkl/wOOrG3wt4RQlhg4wxd84kGdeI4n4IV6G5
ztS6gT0VyiQGrPYZt0m2LZTBJnxH5cHxLXVmuQzoKAgO6whyY+ipbEdo3e5gBOWZhim9Qa5aBkv0
nCXr7ks2B70kLY6ADtZHvjRD85lcUocEl2PKr+BrkX8LB8bWupWvS9ycj0AcjfqGHy6IWTzf0TD3
25n+X4+rcV9Un4J7MMY4eoOpS4RHwnWtePAvdHBBZUFX3Ul29Cu4m6wxD9qMjJ0qZ2OFLeiX5Tk7
bQAPJZfMIg8+3Y6IZUC2D5dT4CD0C2CTrq1cinQGR54zmfps3WvqUefQYxAj+B6woJ2p5/8+c0zw
CFJ2fcSuqZ5wPNgncAtvkdi25GgMtOs9dnCswV6/pypBnG+2KJ7LzYTG5Sk2JGGAQU1L5V6s3ObP
2ocFUOBFDh+p1K6dWxg2t2eFXzjsIDha/9oNPF0JcT0pjkUM6yQ3teZlhtNIUb7Mj8zNntZ1ieYv
yFVBcPtm3aTbMhS1vWZLdZO5d7iW2NJJCbC9lZ/aQ3s4aMBtzvih7qPyKiRBDYmPwUmF58vYbcSY
BwM0dPnZGXmKe9+ImF0IOx6aXiQxMFOzzX/yUQeSnv6ZVojxM4H2by/YO5/4UNAJvbyWasbpGHhS
E082Hj/oowcxrloXkS2k6sjmZGcSYSc9XORrQWgVQR9DgXF0JBGYQ1u89QoJfaYyCkxaXgH1JFSw
jH+CnhNMhAKWFgdQDIIuMr2zzstw/HSzKiLLSDgiBAJOfDU3NWwguVCi61p0UevMMNRrRXNUwhjb
f+R2OnRZzrf9aV1ZU+7TELMpKzhaJOBE/vX/Sj3msn+FehTe6dObiRS8P/62g+r4J4hNyKVvUAlZ
NG7Zq7R5frYBStZQ8anNhJ57ToXV7uKSYCUKjwy5zcsB08uXVrlMtYuSn3cOlqknh18ICb4/4RbV
XNTkB8tXM4fpFtmHC72p7sD1Jix4RZ3T4R3JSDcHWbOPDbvILFkb6ZUNL4LpLGV5D3Ho+fMWzIGA
uTxcIDxut5jsEgqmVyKINvfGuVp19FARe0uE1QHIJa2eDPNOM1OU0pes1uFM5DphLNcLkuiWTKST
thTBnqcSTkdjGOQVOqvMtYCliAtkUp9De26qIK1nwK2i+esObnZrWQV93kF55JPt9lIzQa3RnM9M
D8gZcR+iCfXs8bgMui4WivVMsdiFzf3kX8iTp6CY1lle2IV+fFWLC3Y+TxHCnW3y9s4A7PxGtdnc
7bwsGEoz3n2wQLZX1d/rLfnJZ/gm/IsUV9b95hjeQu6tLUX50CMqLQrNlX1Znt8IUdC4yrff7sLJ
fYWtkDFTMKMnoB48mXR3qwwk2FuoScYrSCWo9EFb3x+htjX9WFqSefegLJXpauSXOigB+aO6Eeqn
Zz9gq21yDzREDmeDDFZGAwgNj2a5nmHjBCszrmGKMvfwqW/in1tmMH2aU1mzn8kJpt6hz3H7KGYK
SHsK0NmhaO/9m1uudoHMEfSTmseB87y0O7mtt6sO7rjK8bFgF6OtA2XfGOA1t+UUAFdKrR3RAkPS
IuwqhFWJF2xKrCyk4qGBMt1KotZb+OmkowxDswvYLb4EXD8UoOpdYxjDcf/YjRd6+uzBPEUBc2ll
w2SaDMHX4di+XZrtL9unwdPsTxL2wHO/Mi3IgPyUGtwryZFXqWxtaw2vdb0MUe8lIaBxlmM500VJ
u9jXzncsA0K7wxKgdrrXfZbFt1I3IJ5i8zOv27kHXFJjDj2WdwMGxdihxtZS9mbxag6T5v5lxkYT
ZWeQG6liKaSZwO/UFY1NwLrjRUTDnk14pso77Pk8rHBLO/o86vudT7rF/TD1+dRacXUA8NH7TcLw
mdQN4Qqx6847tYRC9leDcZZm+j3nZK8WjHX+Ys+ubKem7CwBZrGKT+oEplNmaQW/kACo4ZX5YLR0
sur+B4+0p/ipgTcilRsyPp7YFaMreFFvPfo3LnggC58G9QHub+omkk1NZeTm/+dzyhezX4ua/8A3
/tcbUgk/ml71hdMlBbMKNxnLqZ09yhbHyqrjF8LYkEenAg6YxlfL5NyoO3JIHhTMR3hVa8OwOv+G
MGr676XmCrxqINECor6FqAMOlHG4EX0+SgV91g6o6KSBtzsBtii7E6Sjv4XSMd4BdCXw0V9LqRj7
ACnti5mYoY/iA/CzRycB1kSIMJOM3ZK/ySorcozshavC6yDzVnK/xn5ZAOhTLJzRAuvQ3jGSro46
FJ3Ge3ffUYmFpNLyzIWXC9mVLXj2K7Wi+/SiBS8o7lboWyK0ULmCrHSxvhpWshsi7HmcXAJlRf9p
gRV5edmKNjRWxp63bZs5lT+rRypTir3HCijNXENVdDIlfrWsXk9SMd4crMsGurd6nawwNCETLZuz
LgFZyYFdwQrPxT95cuQwpPrxWj0z4sBe4qCGEAkXPJeKkJzQ0r1p5pZGLEbrtQe3BhBzV0HuZDmZ
Q7KaL/VCFXixeY5htHlLZm5K8y8gfdCZsud24+Y+PUwcqhhXxYmieXC4KCsYyZ2NW6GoQn7R+Oab
xhkYXJ0jb81LUITehsektvGN4TSeZYchOZZc0/gpJWEVLbaAXKZry2nzcDwH7Uo/6N3OEGA7P3Eh
BI3jHjX+ouw3II2SQXFH9JCBni8YoMR8hxfrtkHndNQzpocDmvAaJtooNrMM1BSH5eDiEftjUe1u
YJNuX4Tn8JK3R8t5q+Z7TCmER6O4m4OcRKBcI+aLEKYpCTskuJpFBsm2pKj07blClJeyTpqw68Zv
zaiJYKRtYDou48etKORFlwkZtOIl0l4jmMCFbU1zkSZHL00EgG5HTP121gQ8Q69ZsRFqqfWJiBRz
dI2P2n6dxxcBOA99MJyRBlNJTcfAHOY9pJUAPJVdkqFQDA2p1ACM/hAApLFse9B6knXKcsowTpJf
u8/yNhBc9/9wHJdC99g6tXGk9d+9h2A7HKqlHF0nruWrCY//66Iwim+/A0IpP2a+Ad9sjrqJfbLV
EJszX2aLAq3iU8DB0R+j+shKR+37lqUTZ8NLojh1/ZD3YettuX/zKMNNy1HPoaiLGjF/Foo47Ejl
Ar2/9GNi7dmMGB7eWDp6p24mwskT/LA9eEagMwCZ07ZerT26CMoXaI8cv0uHblK57ZohxJW7Wl3D
mbL8N4JqKIjbxTIpLuVcBXOzDQot/pZIx10DqqAmDICzPqkdP9JKSrbHegEMly//sT7SxGd6a+8v
hNY8GGyCdLG+SmoA/mXajmO46Gx2XO+bmKcAdLkv8YBWdMq3aBg3/fkZedyGYHEL74SVX1Ile9IG
mQqyt6hc7XjhwRtwkef2PacUo3itqlMa5ciNrDO+2h3Dquc18G41EWcXDrq9L7RgH1F6jCxJF9w/
Q9Cige0fNEEWCBFOPOJvTPFYeaE5VCXgxCh0yDsa+J6YqUh7cPRx0GIGVkCaZBvDY/oKD4bFHVYR
NJQZmzMI7UsOM8jgr+q2wxUI5sHsyXMGwCIaCoKhMLobXjWWn7ZLMuDyN6Y7TL7TYskgVnIbrpmF
zdxOqpS9vCCKkk60xn5Tkibxk1Srz3Mg3s8YZplZJjPNZWzOSOVN9LV8zy8t4r5mqqa4gPoegZnJ
EsathzNL+uDHhpaW67UE1y2dvN4QuDjpl0bXcUac6e8NhH1h9o3btKpyn76rXGWF6j0tgoyZ69Fh
ps94wC4DBYh8BnHAO68bS6l1yUAXDXYCepeeF1vDcidh1K4KYLEpRcYvggD339Vi1/ynNNLyU/5e
Yj3xxb0LMIUr6OCA8VHxaUIDC8vGw/r1WKHhav8qwbsdyiqXBSHI4d5rxF7O16OsuJQISYF0ZNT+
J+YGsGTgCX91tbRDns1/ei54M6by5p2j0QfxPti+KHQO5b++fhhjK68P2aiWhjImVwhoe0bEQWoy
EUePCYA63TNqBG+zagbX5dtV2TX7v2bQIJQwv9d0tG4mo7aLFS75aYysFn2RXpIVcKhrz6AEnSH5
5JTf5Y4qPjkGXTQf2oPpDizIqzi6sLxYncxSyjv2yhIOuVmVIeGdpXAfcMaMpqM8dg1boRHIIYL9
mxkkwLh2+ZGRuim2WZG6qccYRwYOjKj1MSeyOLKShmnPiHeN7AMBrJXHX1/f6hqHzSc1o+Ie8b+i
evWV1WtDSPKskp4BcsDLDdE2sv6h0A54mqIaH41wAozDOmeFQXHpl7+pKfX5bU3kZVHechOvs53I
AvupPfpHg8aI233Yo4KK384HxrnWPGKDSsFTdyevKLiUNyVDSIGS50dCMYHYfWyVi5cwYWAsSdGV
2CPMSab/zraMrCCA34pbGrDi6hkKKesqm5miTFa7rLLbQMJP1bvbVYKpdN63hi/18U5ubvYittkq
b5xufP+KUwmVLcRIZhf9/V1ogDrC8Xvp+kMUyiLVIO3jow7QcNSfjVsbjUbaaam2L9nlQQiYoaGJ
6dCZ0qbVGfDiWk/z32vHIth8Ejy60m7ItVGCx+i0byZ/FBFRVxIownTkeSdXPBwfzzTzxgBrRP/5
2KgbQk61pv6FGIAbxmE0yqYwKmK0NdtD1W8nQroL1H6FSK/4j0hAA8xx6gCAbJex4be7wYl05ePW
fwriY4MMRB6QSA1eusKco8+GUaNXIzjtUEgxDS1sc4ecvHF0il1JMAM62JGzJg17KIA9JW9SmTgv
KlX9rA0r1StWfRJV68iKQkX5WEt+V6uhy+2rcPyBJ15Okv0LUZh9/PO6FZw+a9sexIWFlXiqMWOm
8kYUUumbJqFV8arXJsRLKxInIurmMBgQLct4PYAymtUyIWWl0TAVpX7Ee/ZKE8AFvZPzWbX6pBPV
/yNMj2or0W9dERmve3AFWI3cDLukEOxmwntG8QJcJWpHteTRVAu+5CvXvvFKrd8x7SVrdAKXF/w+
6KoWdGXrES7Orb7PH8FE3YhE2kY+uSGY3rob7sn8XRbAOsRYs9t0Du89rNwT0EvLZD+8BPXc2031
qsp7DAyrXYXC9DSrUrL3xq2y/Z31OSQljY4JsGVVhMnZ8odRwMxToZ15GwxgkxYmNgQV6bzQ4ovz
Kp9RaIA1hhgHNb8rrNwGOGsFcJyROQthQUgEcJs65CgpQaF2nXuQIC3GzmQMj4YXU2kr/uFOEaeh
Yp8GfuhHc4QQhVjHRWmp3W7fRjlvtFt57pjdigF5oxVYovV7SO1GOJ+fZI2vCMyg57tV4xDpar2p
y3hGMf6U2lnAcbpGm13eRhccN/6u8HI6pjSZ/vOPN+34a2YL6zzC9hUMVKuC64ouEHH23rcjBlRq
lwuMIgk0QMQFtyWHnQbt+roTPf8BfXjipo4o7BFScthsrPQC8BJt/4NZg3XXt1ka330gZRsdKWAo
XmsBBkwKmWornxqqRF0kK0gRXUOUeOaWa7P+J0T+P1nyMQtMALUXOsCPs0FrO6peIzkZ+81rrTCf
wkELe9TnKpgBq1SiWVPEUkmmw4IBCPm0sQ0ZxKviyRZ54Zr3qSXs3bfJxRNKoKnJcGJ+zEr71WOX
i1nO46XK36/luv348Nz5BOZ2PfsTIrmG0ogQnJE2b2PIIUxC+R5wi/3gxrOt5LHVCSmzF4jg+NzQ
X/vxsIWIW6+4KC4g/rtlNrPn+G2sA3WLMOyVitABAQtIaW3yQ5tCABY5Y6t4+JdRPPA87hgXqON8
w3qy2igkytvBcNDYP2WL1M3gJd6Ao0oO4ftH8TguEZokbc3vi8xoAutPhLs9fBBUn4evqt1vcOGH
ni/UC85Q0Ulo41lH3EudkIeDhC3AlGRmBsJJZLWm7VtenCDcUzOoyXH2N8n+MWhRtqffYg0wnzXh
6nNYH3mBZASf2L+kzlKJlUnErU2B+vSo98uM+lYLWht3DfyHflMYrAxt2FFeaXMixqWeONSitIct
U3ftSKnB/gmrASgn42nN3dkMQR39Hv/heBNX+p107KG3m+X9FquL/2Y/ZUUdhpYtLMJMY5AQCVHc
UWau+EztpjEqyQQCFWJUkveVIdFWXGr7+0qvcrOPjqxC9JfZi1QFt3tUD+Ji7JE7wLMbgKbWfQij
6kuYot+YsI+epNj4WCZmct24r9bGBvy759IF5KtiJ9WGiZaycQyO5dKH5lOirv9ylU4ro9ybVhRi
D+j56ffaTy3yfXaT2regfc5J4UWiUrH/ftPgsGoD+P5/8Pu/tWNgdPDxWKxvbRY74Fp0O704JHP4
RC18nDbrUrgWCZOeLjWY0GNnhm/0QjSulFrVRty5q2sxDPtQgsxs631aqndcQcI7Hxu7GrcPb6P7
KSsf21mU+ZYp/86WotfuNT0M/jgPNxeAubU7r1PDSRBoUkTwObZ8PtsLnmwhIKOk6V0OaCcZ6srh
BG5SgPkpWn813XnoGYwp4J7UdnQ7ZPyyMsQbwioyDubgFlcfe5/JpbuJSK614WUvi1xEO4QUPSJq
ojGgnsi+++nPC0ayEu/E9q3wbfmGqI8lPefQAWlVzF5AwZBYr5DgXyWbPLS6cSAwNZMg7TRM7zVi
VTOCJFF6eZzrFo8nuTMPItCtHI1ZXZC8Csr0xF7tkxUuSBhkuSvqYZsacRx5WrB5MLPDIuEKb+dO
1PUky/Z0MIZ1oGz0HaBs/uMgZAvH0ZgzZ1K9JPMM/cnY4zdq36n9bYal906lFvQggRH7H/5JqLbN
wmuZfPzN2ay1F/K1MF39QyuqL2xX6gd1YmFwYb8GzWTp7YlZSY7zVGa9EQuzkVOsK8KsisACObrs
qiKne8M9V1wNrOTfAV2u/J13Px00ehoFCJwP1e5W6mfv+WVMWNgAIJaHOVbBdp5mBJYwAC1XJbWu
3b+Bn1ElfxfvfQOraKK+slmvFiWkaTcDIu8xNwX7/+1rrVdrfwqvxuaZ3qLQhjsBehWmZpEJgJoJ
wtJFUrOcnb/inADDMl+5Bams2xaVgDtdUjrJMTk7DZpyFmkAWX4bdinLLUlyX1kF/jRX6iOYdbqd
Es7jPnmVmqgVUVCeW9jN8c/eyaiRqQIZiM3TMeXoyNMxxUuDdM8Cx8cy8rBoANw7yPhZrNZdjnw0
/2U8ER74MT/Fearu0+Y9jR+7Ipedu1Rk/nHBizyApoHCHCifcPWvEWuGSMSszjgtBJRu4Qx6GTni
zLZcWdgV6zBARkdIzEP8aOiktZVZbFflkAJAfMB5NvFm9CBSx9+rETGG1r24fvMd15hfdsfVP1rm
RgRTOsdAoJa9BGOpET+/Jbapvz5uF4Ql7f0HvyZ2PxRONpCJKQqppJvK2qNhJOfGUM9WZJUfz9r5
X1q3fiv9mSUjG4YN4cYg05UdhD11DMHVd6sTODU6+mXCf3tgixiiW7b+0r20cXHzuAGg/zQz3d3J
mrnqiuiMAtaZMp4YKhXZX0+ujSkm48fF3cFVgx1KsMeaFV/URYs1QxQoSbJTIGxNOoi+SNe5GEXY
W6PBqfgzf7ylj58lZtpUjnic5XOBSO32xUUUbfZSGUPk8Wxy1Qyd0zGpfRxINl6tSATUe1wOeZQ0
SrJmpgWXBrKOi+9a35D2BcYLuTjuZYD4A6OhGmPT/wRbJPk9Kk1+2ydG3IQuFPs7pQfo9bdHrsts
Ikk9UtmvtYAlMbQdC8YNckaTPuCczfDmW4gpG5vjrcd6hPdI07HrbilKDxkCPVBvlm/scMAkzX+f
AplwGIbup0lsocZwZlnBwp39uHnehxL4bz5hZ4kc70Xuh9tQ11PY2q8eJfSQ53QnK0Y/IYu/bHiT
DKphselwS0oFx07gFiXxYRSI9S6DIwnsiUQGxW05LuYSyw8iRHRGdnMtuBkpLDIhJRPGw0ZvGo3u
FPuP/ovzgW/cGlufPr1JRcfElW4JD3dFW96NHmZCMpgT0VRMzmm9gNipcByK5xrhd90t1Br8lpNc
cNK6nwtSCDVeAPfVa0Iy339bw9p2mvdegLWhhCWs+MpX+uBcyMJxQD9vvbAxIfFbOEEisBIK6vqk
51drY+3R+D7hAcJi44V6KZSpt9MvsQ5oMWflboYGLnXoTqme+DXKz2FmKqMXM8HFcY3lOO5HyqRl
Ex4yxtzrFE9gtBUysY56sMqBdWhRMw2qGAT8PXsvOWB30YCIOXPk8yTGqwwevAZjD+hv53y62JjF
MssZ6b/d+g0+T+obNs4Wjvm/YMB5haZ2p7XxxcvW7/3DKi2eNDAo7cmbab6MSQWGEHwnb6d1ghVa
YKylq/41guxOvw/G4X1sq5uM8UmOJCHU0FG7TGBCi4KNx9Rpe0uIm9erhgrhsGKYg2FFoGTeUsLd
bWTDqeZ6EXdcdfiOdxaSUE2SGMmbBhbAgxK7NnunmaobJzI9sdBMqqRkkkHnbYzyggqt7kuR+7sW
27LlNHW8lW7T+iWG+MRMt0o5PKNPY+Sawz8a8oz/1DJIipk+pBJHjHFPCMWpElJQ0LV/pEQ3YH/j
HCexuLSpEPPwEsCY7eyVA39FLhEZrZxPRABQQQm2RpTfJLyfS515ThpwtoTMjCXBvX57O88XDc8L
prG2dHCXt5CVWGSpNVPYiMLc45kRy4JS9IEHv6eN1UKXhgcVC6B4NRJjrZbT0uwQesiiLLT0bLVf
PJXgfs8cxpsr9ALTtRmdSwf+LX7RZIlw8NhE3Gaj7/SkubXiuVc26XTaPlZUqlkdGJaBW1X7pjIG
bEWY9ybinCebKJc4UClWvvXywl1TCWCTXNWw/TqkHIvWWajeP2Hqn/cpJCKk4iCBQ0kpEDcmi4PS
iUFT+Llf7U08W7Fe8nqRk0gHNGyrPX1FiHUbzd7Z8O8YSZM66zzA0vDTEZ74xSf3aNihUU1atS3K
ZWBe6GkETpDGnqs+J5/6DBXFih9lniWWzlCvL0D52XYCJty/Xp3kGMeiX5HUlzIUhOBUAHjx6lj2
+OBsWeXgFb9eFo1+47bEI2HJxvHz983tyIlD81wekTwlDjw4dF9NpACXNX6S5PlitILYgrC1Pa2t
S0GU340ohjA4/67m9I16wUgDsHXgc/anyyJUAKL407v1BSVutJ93cCHA6W8fAeEFF7K+vPJX6+Pw
bqv2wCEnqPbIqYu/jfKHf11kU34edwCnZmeXoiqvUiQnBrV9Xpp9Q6iV9RzDYVzed+8aS95YrWC9
L7kPW+pg5Wp3YEWnXaF8q1SoC8hBCyzj9bgjKYayAynNzuX/H7BBjSnPQyddpJbS2N8SgvhIbkDe
TBfhMbxZscgR95ahP2Ei/gWDmnwDt0ZkpJKhOlfLJ6YbpLzrZDpsj6YJVUznO+ZdvFtreYsATCAu
0317lq90Y1UfA0kn9IDEo0GZGD3Pyx3ZwGstxvZTtW+xOJ8kP2Q0ewibn7KkLtMZYiZip4+0JyCQ
64UeDyzQNW4vHVvPQrRrO63B5yv/yUeILCqUSwFjr5x6vL66DNThxr9EQ7O7UXMc3g+Kny4VD5T2
7QABnKTv8B+b/Ptoc0phOQsPa/Vbtp3J/PTsWGVYnYP5jU2OED6sVywNj/FuInHi2KA0KFLBrq61
ygtG7ObxL+4c03GRJiCidXLOJYOxmk27GiCgRN+ILxFtYKqGiQU94kFHppbMV/BQTpm9KzEVLbMj
tbvZRmZ5IGMUz/m12Rc4NbUz7e2wg6Fbnp71Qbf3CUckmDVDRmZAK7SM9F/PTGqy9j6sPBfMD0mY
Wi/9/ZiKoMRlvQtP9rvs36BcFC1u+jpHj4GXSISADjpNekKL2jvGQiTyaXDgagg/S2kIfwpFYJzt
GSJPqLNrNr5K0g3oET7cwnB3lp7s/WB5e0nDJdPBi9kv3S0UluVt3/1ULtrqQSxmRPzFWMoj5hLh
rhGpXUerH1zAREyi6cHsGbDPdFj1XI5P4T+U/KGCQffXuFbert47fUnBuDMSbVV6ccrjb276kzI3
TQEFJCBZzZDWJSOMM1gROfBiwccbzVXgY4mSvXibfV3n4SsLHa0zCTTxn1aP3MPtkCqGsIgncacF
R2vDTXMTQzb06CIgW47XuhDAqmigGk2Ura+AYkCjfGT+VNhen2h8R0IBIpfOpzJgCqIhCQF/dUrD
AQNtPHCah8FXFeea9JPMnvkvig38eFAAVYSUi/hP11HaC160nBjvsIwGDHW3mOfyoUi4b7YwslZN
bQJWj+SeI2XEifMNexZlY+xYJjMmU1V4tB+m9DTCPxae9Bw5tCfakqDWo1kaboY1Pzs6t6kthJtv
FnNgce/jphl0oiY8Pbxf84v8EYx83J5Md91jhU1BuCt2uq7qqPSzwFttQt6opHeNTLBKHwo1Ibh/
kJ2q19cjTAp0kJq+zQbp5v1hl7ZZ3vW0OADgTSbUUP2jkvUw8UYm35tHT9kPecL7JvR9v5+3sOZ7
35iWY8qoh1hPmDqoz3Pe+eWr1j1fFP/io0HIIs+mX9+IXAnz8pK42C37UeNjLjqsGzFeOXD8xAaP
fNDozNLgn/6KS+3w9eoF5Joco90fE0cXbL100ooxMLS9a0Cof9GMqKUWZT+ovDYbk1z1WixwuCP1
jooWYwr+46Bbdvw+gnk8OtEqU/scbf10Fwc+IHCtychRpEJC4DdS4d7Wo3HGccuYvLoLzfAskvWb
5bNfnK+ushO4RnGpVkx7YpHkw80yF8Sw3YKMFROssnst/7PNfVrKHrIJUdaVV/8BZU0hnvtmzpFJ
539OmFsPNRKm6d/JP0Ixh7z9iFjyJ7pqQQOzmGdle+lmz/x1xZIVNZZ0zN5XT7wM7m6t+KvY8ge1
yBPnp9bxcsdI1NrZBDnf3r2F0NnMB3ezWJB61G66SWtpUg22Qcq3oDhNT8gMmyJlk7p6rSPDgkkz
0xszsdiWIckEPvrzsxUUf43WvoyXdUAG+Rpg0D/FV9fqK/JpCEVdRsz1cHhAJL12OEDYlRZX3ifT
3DzPNR7GDmV15ON7OzqE3WKFN5RCZfh6q4tXrO3XSnc4d/nOPYy0Kl+K5FmtIpobYrMCiRBz1wmZ
9+gzJVB+6tz6efLtPYolTYP8e/bqs6/aqjwN9SRph+tLylnvrw4C7IfACYtooKCN6+Pi+f+uGB8G
BiZDAXhclB8QTtr7Xz/te85JAwxKXeckU4dNDEQMwoVAH1rHV+x/C6FyjTEVtqXU9iPbFYFm3pNa
vYf0mDWhjRSxe4njdpBO/M6DPZPC+nA7o5g5ihupit4205SSQRr1MvWkLJhlvbIzDMDnZe8D+eou
SvupoZKxp5j4GbwBYlDrAJqsRiIDqhdrBV4hVmZSnDcDzY8Q04HB6PPQZJ+mEDqd+zj6EF4mErvZ
liYuhv6B+haYc2zRWIzXtf0vKKzGih8E1Vf40zz9swvQXYN3xY5viY51Vc79nw8dY3xkgkHUe4d2
rGYOCPZAUxbly455RgEp3utty5PgpRs7rdhfgj5PbTHYKIrgBLwV5Dx5Bl17eUiR3pyoJlS2OYKH
3H2uNuZZyuzsrGlFRf/fSI9H7x+RlBaiGE56+LVr4HUHZNIBKUsiVobTxtahLr3gIsVgWf1QKmu4
c7PvqqmbMaoaGX9HW5Ohh3zsuc854D6oQKZ8MaHeCgmxDiD5CjHXecH0OI6TIrzLONHpoCQcNNQe
E1xUBFJ7kCWCkXacpvPNzWHjXHYDAMonD+NITP1FCkkt4LRqcnkguCtjOfh0mui1kK6gknlzm4sS
Y/I9hJyW/eQHzMQAwpLbwNnusCO3ljrF+BT+bbFtXZmPASx3bPqzZGbN08iKntMlZyyyZIiWW+7F
NmdRmP3JvLekiIR5gZu1gF9EIIgDJGLiwm6uEtqo4Ju4AzqI4X8g8rmk9ya+RrPlbcwaleDgL2ng
nK683qBnz4riYTT/HbNPC8sMMp6iRNngA4K0Zs5ecWN1npTYDVuaGVDzb+rYwAdDMwCqPgiB2qQ+
ayaI6hwmKVgy3+Ub2sq5NbpidI0EhvgYrmaWGyPXfKUN4rmincy6ki7ff5jX0equcI+2K192F9iR
ow+Lx9WptAvhoD7yjNbxi6Pv2pTMh1Fcrde9bNg9u6yeqkDJdeiF0MsVEn5h8g9/oOx6wRNLP2SU
eFc/wEMdm/8OstlUYpS+VJS0fiV618ieIMT41OQ+ioz3JSRvij7xxaQE9c7IzC3LMcO6ZGMOIwtv
qpRAxTpDiIUzS600o9SGluwVSg5mU0BnxGajI4D2VaMdJYgtoL8Byv1gtq6837QMKvN//A9+p7g9
ba9tF1wmpqmBXimuAv7qqKMSMb2/eoLIZAHNp0RyJ0IzsvFtWHQKYbreLJ8QD3OhA2eXVXxsQAOI
auPNjm9YPlbDi9mnuBtEBnRF37ghwPxN5pdp1aaq2CTkwE05JcwdUaKNAamd9mjknt9K2N8qw7Ki
V2nqHE4Ze9O68QBNFwCuQIbpth6qLiw0f5l5f0XhUFL+Vq1eV8HsyWoujmQIUqM5O33KXpn/kvjD
RbqahdGmL40/kl1VX1ehYmHkuyTQuriXEgFpy06XWBPOyzHyIyMsT8miT3lTswZU6LWujq5bDQ5/
OA8nj+MWvDUeswqGXVFxpgQY9XL0FuhqMmpRiBhXEpJNxIMVK9Ts3bGOLIgjVM4RVCkomMU+af0j
GIT3Kgh0z7PsFp7vkVdbBZXjifxyvkd81B3p6C13oBwIfv35CL/2nBwVdhiqTcn4OQYfrBBWFAqs
1LT/UXybNnJ08T9Tf6Zc/EDxWosCJYZn8nOqf33oLCkPpXUQtVgkYFA8h1+N9e9yS6IrWd/OMyGx
/tdITLTylzZDE4+yQ4sR3JsYsuf3GscxwZ7hkT9afeGaMqvl/UTA1dor94qLKxVQAoG7XHN2HGY+
U+2+199uacqT6STneVsacp4/CCQlI4/zxdzszIoFhirRnGCa+N671AXKfjymfGxBglTqxPLt9qjI
z8Q9ndkZJKUNtmizW4tqtCPxaRAq/CtvnVhbRVPtQ2IXIMm1TVndOy2lMaDmUasL5UhJMcZ8qh2G
omj1KQAIs2jvhl5bUDZLWmDfFABIdPn9gZxTKPwrBIeocD9Ynq9YWQnRlv5UXBp/Y2Owi1pDNZX3
kNdM5yHLmmHCrvJ3dU3KE8KU7wbTqFUx6CzPnZrS/9gHQsQbTBd/U/iT3vnSpCRL0rIdT2dL4JYo
J9Qpgk9z1ZBztxb5v3DgH0MFFXiHglOGvu1KlRgPSQOVyyXNNLsJk8HsjTfLsupMjsUSnb1P/D9A
Cr0dIx4Ikrs5hSU5fORIU0/nFw018lkLukffMm5zEYQ/xTuc8CIvgZi6dyIGmVge3pMoBCzLJbO2
18nLhjpKwq5ot6hefTsdQOeAmEWyDERmOYNLNPJqYMEy/xaecL0tbu1CXXISBXSN1KuuMPgfboro
CcXfHby8Ytsw11eK73I8HSFpZ6qj7QVv5YyOViPAsXd4xkf1ontaz3+TvTHMGUSS7n7qvg33e378
fzvQhQoTsqm99UTzXwUREiF1GVynryGWjMTDvpL+QLAa+OCb8ooHcO19dwfHRdxp44lFrqvfBu7M
0oaSOpvWCDmU14qRUDfRvImtEmtpiFVaQc55VTwjmePI2fcGP1TcFa7gcNvgDxPIuTfxs1YEC+zT
re6ebnEHri4W6+goMEzcVPAMfvlTThFjb7ogah0Ri4OMad3nfWH4l4Vwnmko4yH3RudaBAenRqhW
j6mmFlN3YIoIfFJnmUtuPe+4PyNCCUzNGGpWyB6zDPgTe4Ig9422P4Ln52O5kzE44ID1Phi71Muk
3e7wrOz6TDLOQH6SrEZGwH1c2SUHZoA2pfP1kHffSM+5i0FxDmNX+2iSnTbkMdyJky6rrfYTVE0D
Sa1fhybh4/xabGknTkB1N75UFYc8gcXT64hEsZRVRXpuvb8Kq6Fhc2Dy7eAWV1KGQuylYa3pu1gm
tfhYJkCcYKYZNxBo3mTJ7DUZkGU2Vgk5hTejz3Jhy6ZOsMvwbsFMbB9lfXZRNkwVURwk3r3J+Vgn
1jRoqBWahdqDLTSxUU/VZkfXckSw6pW48rwTt6khdUuWWN6SD3I1oysoMgQbImWAhyImKsbScwE8
2MLrq5zTpunICsSAB0YTeVLOXehN8OvZAhzdNoYaO+IEhtZT2Nh7GeSGdDpCMbY5o3DRk8szAbaG
ac+apq/SwUau5OjdTcZ+A1EKvRI7hOc0kfXcVpmeX5fpLHHms7+/pfH4rucfZDN7dYYx8nPfIAOQ
5aPnEb9KOYxgHthAlZTntMRlfE7GgZkUh53eJk9yeZfqSIql5blYvT53RsR/MckTdsFkJDUJXHoT
GKA23pWdsRe6Cc2C06SK62gmoW90CMcJN+qwitgk++TZbI7mK1MrxpBtYd+XZLiuYd3iJ2bZ1oBE
5lH1A6ievVLpdv+DzGXLCwfxObQ5iJo/1T4dhFzPttZfxFJV1AZMz1I+DjYAHHNpy9Fx2sCi42oo
lf7Y98r4gTzwzUfqwQ6gjRv20whl+UOZaTI4nB08vGqT2diHRyiSOsIyLAX/18GIKM42VKYp8Ip2
Y6A13qYpBUHVUUlN51zrljMBXtXxwu0txvwgcs4pE5Ff1AJqNvrhCx+Bke379oRWYqJHFjX4MiO4
BQVNr0WbjodBOPanyEgmS+QtB2+vjyWeH02i6zPO3hxoj1malsvzIoQNljVN42YjkrYY3oiphzjo
C4Kui9Z6Zv9PuidmAges7BB31Xhi27mUOQWpLf+7qEhXhRT3d/GhhRxN3k+S8NzaOrmEywblXLTz
6FT0KvoRWCz8f0fEefxe0PF2YoT0RY1Y2Uu3EYs4hGbKQaHFWHQ8SJF1dDs9LJkN+XUOkzOPJyjn
2D1AC/HyLwRX2R3jdo62x/QPRzbYXWUM1Zm+m8b9NRsGOmg4s/AlGStmpGm3mjUI+kiU8FVU4m9C
3GR7Qh4hvzeNTn0t+1oMCNa1zonedXmUza+FD8O1vqmHjX08oTsUQdSWSMPe4+BOOlZRPl1hZDT9
0ImzBcmp7VPb25vBWAFoFqbW1UljR4tG3qLt2It873kh9xz/e0U6pQKCEKOxa/KWl3l9nKoojg3w
fmygmi8qdVC9izI63vMhQRdR4XG5GhZudC/4Qm8a05eNqI6RtL0Frs2XHAPTUJngx1zwF0X8jfE4
hbOsXU1T/RrHN4k4FFoMLRBAakscweCAPKUDs0/6hWwxsEWh/XnlUnGpg8DpT5mQ6j55/3RtXfOp
Z6Sa5c1W8nZV8IqEgJCNr5JjPQ7LewaE+ljS8HGPZk0t0YySBMVvUi4z5+9sMmFuTIbjdbZxN6u6
FoZWD0gHmXY313GCW9nujwfb1yNc17AsYUd5GWAFVrIzBEEjO1iwhJ6C6GMYLSgLVWcj6ZsiAiwz
uJB6eZzKDFizodWjuQ6149rvGEQCZgqwW0I/QZRtBrkFY2Htc3kS0/uxmDCfFsSMBvMN2o/5Q3hT
my8oUzVDa8PcN2tBNL3NSg8gLBzKr/ovRYANuUcRA6pDNXhyPahOqPd3wca3jaIP5y4IC/KURucN
taZB5LfIGuKFqjyQNQn4ChSSpvKQ24jsSVdb7zyR8l5Plsa6FmMFZX6gE51esv4ag6m/SQqcrvFn
Y7ttIDFe6mEnytbvqkYifEiVUh+fvorY6dUtIiIa2TtCthU2HAVeqytPtUQyBTTMRndK8205AvoD
aBazfbxE4NLWCiTMLw+vHbtmo0aTwEtTpymrwlt0CWWACqO+wWmd3mR1mXkZE0CLkY5cFyV+PcUA
eOeNkF0cH7G1xMje1IxnFiHq/9jzeRKuU60xRiCrNaS0oys0ApVPCnOhsBeuuy9sslsXkKCZcRQ+
IGbSLg55RMTtIEqIHSf8MlLFxZqbxdGax1kieI8jY2PMpbi2nmWypCLus0joK3FQVJObzFDsk21e
GVpC7RQb4u1oWpP56/25UIlgLtAbE3rVH3cVDwG4f3ET/w7s7UYUU8Lj2BCh5eDMTlHKyhI3R+Zw
hUPT9s1oFZSY7ZTA/JF/lcImmev7FpLu1uH7Tk7iBXOPV9NliOMhwvuoDwFAjQai6bwdzdksSikd
5zApQ1Lderju8QgamiHrG3b8ZjDJZEkuk/EbmpQdfyXEYSlxB5ehJxaDIx2481nM6wvjscWobATo
sR0tID5UG4GPGs2Q/SsOzgPQ+C4qVs4tYcDq3GnkKdiHUo46bjE7Jix2NrBH89lQtVHEwn5EfnDX
KNWt+XSiPwItZxKB/5fgPhh8ysowob3xJfnowxwzkCBBgf4z1PvKGj8aGfLXrYIZO7+jcyG0y4Ky
BroTTM8kh2lQTcyDK6JIhYNYffRQdILmSYOAY/q4ItxT/hqjJ9+WzXMKa38kZujs16UUj4Q1Rf1N
Eche7eDwVE7WFNTWtAo6ksmAdTyXwMy2u8Movk6hQGtR7Y9HRou6BazEHVWIE8nkOMiuPf8rbs/6
gwg1y0nYaXWAfkUpSloYvA4MPsmH3Sa3icTPKuX6yDbfzGu3OMDMCdo4cIrhGo+1pn6ex4i35w6M
8YQxZmkJdAy8vjLW4cLWCR8rTYNZk4I38Oz36SKSw3SZPj2T0agZy1uoXKPLKnjWfi63e7gN0+62
XqbCQMKiFZ2MCaUEyNPiI8dQcDJ2yl2wpWY1cnnCVM4oYLVDvud14NFOcG+0wUtaCVB7UAxF7OrM
+JSyYS/8KU+dU1L34MUmh9bl/qaFBrOwk/rYtPI+yBQwl3PnMvmg3Z15wA7ROSP79HfXkTt0MIkd
XIlzmlqpR/nV0Enha+r1ZXW3ImOOXYT50Sljrqfzye0R8EZtGVFdek+BThXYgw5nWCmh5sa5zXWr
vmkw/zLy6E2vOHuMKeocfw7DGL2ITyKRQyk9UK+dqYuZJSdaFmamt56IzsL42OYaJGvHRvDfRaOS
dRZf4u3MVvpmcG5j1ATMt4cUbILMV5/B611an+RfpgRm6hAUyLRDj0u/EX23+RXQaeI6SbqZpl+y
kvdeqBhaNn40M9bYjKC07lRoGkPmdBo5gEDgzynZ9oRHVyuiKf8maKZRz7axPT1mbO0Kb1phWWzj
FMzYb/jM6k7jVFLXSXk7VY5QHEUc8c6OY8uQKR7dm39dz7Jk9LhV17M7F1Y65plgnOClxNQrFLIF
noQ3CNOogk96HVC0FiKWgEFNaDOjuMduHHacWBTDuart/amM18oFfVPIMrQ1ylspMPco4deKO7bY
ApXX0A+z6qq5BFl/QYOA9J6TWuPKSeWTQ9BJ66LLW+APYr+gbZ6R41KXedOLo27vu72uIAe13C68
FXdkRSj6w0hf1aL4f/yV1Ldf6rPslG22PWdjNuLRl0jiieZLT8BG4wYFVMc23GzdM+JvLai3jAnz
mWEQnBLIMOfgqOgQW2/JBkBX0VNLYElgGBZBsk9RdUDC7hamssICi/t0YxYOOHoUlp61cr4kqiRE
adNyimtnPq4GPK+jkxa3CwwyVeP+je17wV4w1k2E+9e4FcozoYMU3HS68SO6TdVncwJAsUoJ3Xid
KZy1i8eZbv8QPc9b0vQ2LdIpGYswK8LEJUFnbDnPa04sVTPy51CaM+wQVcTwNAFmWQBJ/UFGpT2P
P0annorRs0Qpp5h0A+zWs1ouHLly/X1tgduqEeNOPqPWhnPB4Pmpmo3Bb1dNTCWKtW6IgOgKaJ6p
wM9/VXfsycpY7HOIhTfwmVbbuIX37vzEQ9Q376lm50VylSBGoibdYcY6Bj4eDdKvMKeygAcezNfb
W36zGpcTOkyGfWu6eEuQbT9Mb7DD3LXqMkTm8BTwgLi4VW7wsjzZH7UVItVgQ1EBAMs8qI+7D3QF
PbFBqGpLHpk3lBiFaHzrd6MiYpaNFPJNQ0rj+ZKcltg3a8Q9Xol85A5MwKHwostBJ4QRKz1GQPeW
dV4rMdMhdpMCKvQmsSO2gq5TnCpohTwj4SptH4znospo4YnEVmUSCsoOuqnr3PbHuynqJO0DileK
SWb0snhMjGwtZUtYBXXbUN0P5Itw0wFhZ3DKvWmMrrHdMCIT1y11ngFaJn8UQiRvsC9XrdmkB3JB
1oQN7AHv0JL/3YiWWfnRI63emFXVZZ7Xl2HO86A6mZXVxXUUaI29QeAYR5PyKU3FoLYYA6KJcKJ1
XjTEpIi4YHnM+Fvv/P1JiBcpTyHdpb7JKifI4sNOnQB7tNj+7hyFUkP64Xz3KNJ8gcpSdnvoh4tt
bnWX1VBGKRUE91D3m9KwrJROmWIySO2vstInuyZ+/jG31bG5G86IBqhQThm5oXEMoD5+HfowODVA
ArrNrwgSJvayk5UPLfXamV0yTZup+aCuNwwc9wthlpZ6OuTrLe0p5Sdiff4jto/WI7H98a96ueL4
BvDbpdrsQM08tEMFd4BATHxHzAH7etj8hf5yECExCbhdFqjJN5meYyhof9N2CPSb0pve/2lmHmJ5
NKAum1qLW/vbQrmCTkSRx6L+q6VIZ5O0LAm/hqNRtBsompvbjxGDX1dBg7Ec8hOEfGUZenGmx1qL
kBVX/F4WgSiYgWQYVPw+MtE52CS4hw6PSNEZvpAp30mQ/NSK+bVNxW+VRUM4rBWJR8kwnzsBp/cl
1PpmU1VPRLqMBetZtxJmS/qfg1vHmRdMCDJmxMGCX6aIezdq+fR4NsXb6i3W20iYa+iABa8jm2MI
Fm+5xyTY4A4Y823+riwhr/++q87SNebz8tOF7p66Mlb8ZliYxjaXDJDUpHnU61l8FvOR8a1UkwjS
iOhcYSIuUfyHC5YPOWa7Spgqjq/CtEaDBCwZYdurESOtJgrxFQxdQoJjnqUc3esbjrHztcMvZ8JT
ltSng2dUNZke8CGFC09qlJkoGyOpH90Fz1ha3fa4mE1qD4jb4oeCHuGrAgJFIADjK0V/I8A+TNhK
hbXgLnzkn4TuKmdf/WMSNrlOUcJhw7bEi3tzec2J/DyoFAq+rTia/xaKCPI15SAlUKcly1yTXVSY
PX+8EFOGVAcNdOU5hdgS+xtstUUhta4o0AzYb/FhB3EnTOpIGBKVuU7go9C/9IIU7DrN6wl5Tmzx
ThOnv/B7KUSxzg+fowmUOnudSotvYSNVznKmCVrwyRiObz4d49uiM2SBWUTi7Duspm1rnazir5sz
Z7R+FL6lUWTv3ogmpDgYxQKuflQDG7jNBCjyCVJNrzkfSfRkSnnr6Go0W27hITMGnlnzyK3K1l8K
Ug5mBXSZ+ByHhGcmYdRIqamoeKuVAZT8V5XT1nJiQDJkItOHY11GLkvKuXwuTEL7F4qWl57QDNsU
iBOaP4j08j11rska4stBYlg8ThWmZ9Gx0rSXiapBzjzcGFYNnIgJjFxexy//1Z7hDXOBnsCoF486
PEs6T7Yg7DfldfrJF75Dsl8MoHB/0gugjDXQYZlbNBnVETCKREnnNVlBPm+h5Y/CMeX2jSYfTDlk
+AtseUYX3sfAozbZQdgk3cfUww9udF1L5XUbnP0djn1BN4qMzoKXFnw+KVL0u8zOcpNDD+odThTi
FiGyZSjheehey7uHX3NESmJONYRwONyE2SsKLHt2rOnX6CDsO4x3c3qENqajXEuh2WO95SorP5qO
IefuwpOl1HHsUserZXVW1d/+EpobJ0k6djHbwOU9yTXz2d6eg1AW9cmzXMpY1asFOMlZaJtTzspI
MGBCPDiHSE6bmn/2GFyQ+sq3dew1gF0mq8JhQCpfQJgOszFcYgol8S6OTM3jtL48GvK6PSxiyy86
LOGFtLqkBxmA3uGRhfxpqbxrc+MHZcUv4ku2wHpiLYdBawyCLqSEKzpPJwFGMVV8BoCmfCNzKOCa
uwMbrSP9poPsH2Km3aRBWWRyjS0NViqhRjEzW3nTqZr/M93EigmgijBnkJ5puOupl7DiC+j+HeKU
vWNkU0fTQLBU1gQo10OWme4h9fiDz1nafMhcLYootN+64hkrJqRKIIeNgKyLkCQMITSvIZDYjmNZ
W8WnfiE/3QopsE2gOlZHsp7uGucd5Ww3q65so1ry8uxmwbOaACxUu2dIkd14a2fQf2KSMzd/12ZZ
7dUVy5rt1/uRYzGqommkcUC+yTOAvQq8DnqAqDgqpyhtJxR6zMwGahcuNIvqsyDs1dJh8nhzaEKu
y4quWmCj2mFRhMg15MKDaLqcbBRwZq3mMk9a5QY/Pzh4H+74uFMNIZ7FYNhj4mpegCPlBUIhChi1
44F28SQqqBA3RQWS5frZQBDv1+rJ4+XVxUxVYbbcblLJyiiFT7Ymv5Hheg429Y9n1OyL4IxzOT11
CY58RYnnA24UWwvnBX2+OXxlVdRJ1fgTsy3qKnSnlJ0uPBjn1U1nY66TDudwXA21Z2ky0i4RgG6H
/FGOXLQ8HEwjIeIY/kJiFwUds8sjxc6XSXU89ALUX7qY5CGRTSChJUMsiPobAe8UlCjKirq4xWGa
EwK7sd8craSFF7ZkWYHll15u8eSRYj1M0NPqcOiT6+sl/zpDcR0kDG/5qn9uwmDnUdU7cltIY4hk
SIIVuqBbbTQBwtKangCW1YXx4yzTdfnaA8IXRJIroysj710rOiPVEBpfbsqhKq5LjTrO6YrMBKzZ
pGXf0EKyBzyWvWeMZiKhRPZeqk+4rf95lx/ByP2jkftLsSqMV9zpOztuaOf3+lXbQLwaOnzNZl4m
syE2LWpAiMVcuV3+drY9Wq25A0BEKPsiVrTl+JByC2w7Ouzyuw4SyQEjJ9asoCTsDmtfhO+aIQZ5
9kJ5BHSYYuXRgWMzsYOQv9zsQENkCDPAeyBioCPSKr4fcbVLF7jEluq1WheK7B3DFOYbWrngdi4t
EEfOODaIyEmZSyQI+oWG2vB8nsD//tbUtSah7hBSZMlRl7mdlJQrgBptoEuqG7iYCUI3sGKP/JdD
aljMhY8HjB/yAsv751FnkRoePdkEMC4aV0Pl/MZLbZWq47ZrF78CwfsYLlNFXuumg3z/Z/r2C7LI
XpZsA/Ws8iqHTiCtsjgP5zXSCdv42epAh77o4BRCjCIWePJFfcPWJYn8YupKbRAOGOBDP70eMus5
f9kSF07C+fYoSZS+g6e+wfZvXuMcD8Hsbt5KXtIIB27MNQ4dYPqSHga1CCSte6VHd/LN2hvw7PC7
jt1CTTxDiVEls00RmFyH9i33p5eB5N7EaXznkhypyBEaVuyCiBe63rRWuHtDRse5CnQd9hG8qo2A
ontPZmarDC+mYZoWH9c9oWYHkVP/D3bKnSnuK1KZsCr4uGCygHitN6IRi0j5+mqr8YTLurqbTjD+
DPxQKMYgWaWhtecnYBhgzjigHwLFSjKj4ppAlkk9x305ltt7JPXRTMwlaVswDs9NyD3RtYL0XtX0
FP6uJi8Z9lzwhFD+ocVf+kvx32xTvarK1MIblc4Ovh6l//aD1hDops6d3uLpgdSVEgP6ck6F44ko
dr4ReMNpIISoiVYNPPRmhk3Uzl0O6Icfx4dGqZDqvbJi45dAvi1xDaspc0g+9fR9yS/k2d5ETfOR
eL28pe7tH9Krqd1dU0z9SYKQNu3gs1NIA8+PY8hyQP3hsnuxeHLqoWhjRKNQztFBiUChbT4DT3tH
fe5y7uNBR4W3pxThY2bOOTmVHkbTXqhhTausk1f1wQARlMhvtSmMkJj1Ot0qZUTiDqWuiJYUVT5f
fZTlbkBKP2o/TJj8SVZ8BXJCWHQ2JMURmsbXMwOPH9osWpzUJpOC+jj0j5yPC60rRWzNasg+l/nC
oOwbkSSGkM9ye5Img4TFo99YYWrKHRmkJX1AzpJIhIMbfEnbxiTsgH9JA7u5+w7JCcaQG2YU7ag2
1Ihyz9gjd7Y7yVSycfe8x0hpYEc1K0sPFXMgSzox++Y32uC+OsQF82EPxrC/j2NRawIlL4dcc34K
20cz5LonPPpJjZDKcjev0hPBAI20PRgJv0/0RKgwHf7hFkxOVjmJda9ri7cB9rxD5e+eSATFbuHa
N6WmA+Bpz1l9GxOUAUsOyl2vW/om7H/LZMpAZxN4FqgZ3QgZrQ95P3shtDUoKZPJoZlQUftLNP+4
Kl4cODqILiLPlkyWh522LlaCsZ9Bck/X8RAGasIbPXTW3d3O2HISTve7Qp9kSsxts52gMWU4ZRuZ
c60q+xL71N1UMuHkj33gGizIDBO83+BsEQNrfm0V5cQ6ONgwXecPeapreMouYgKA8IF4UibG0HYT
+p4fcthIZYFxaXgt3Z1YHPDyvIwH1TX5LdD0jpB7ZSE1SdXJEN8XDQZ59ahdoAGTSmJTh6cJ7qGK
eAiPAGuMe2KjVGhFn8tFoiT5p5vROXUYc67h8iqeKxn7rLELddAOxjyYrsACW5+IqJY0xprNj28S
JA51prVSjb4DtS5CZycc2uj/XFHP4ne9QKgmTAseU4y/6Lpw/11EXFlCV2uoOfDrNfnNME7ZKXvG
D0qCL52PaKB6/RuVOrYf7NTQW6ReUORIOHDdv3bbFMdA/XKbqWMdlUn2o1VMZbpEgF3Vuhth2uhk
rHeuS1zOfr1/oS4kevNStyn/vrsqhMsVK7o+iFvV5MGrqBZboPafCLAnu9rgKQYuK3RaAlVjiybp
pvSjoNXcXLGE3RWcGF6KghJnrmk16km6sFJonOb/1lOWL1D7xUPrSl2Mj+auHutOZ5+eHigaOPID
I3QPe9OOSYBoRXb1jW3dX9oRxcdF8ZvDWZdk156cWP0QW/NQnNeJMNDcS2fGUZdEfRogGGOjBS61
fWzarehZma4SeWgNWhbdlsMA2FDBDEpYm0UGhDavMBRjgwTtm7bLLwrBPoP5AQ6IJ/GrUnjdKzwW
upPmTFKL+XSMcWXIVDAwV4urZmcp/hN4WznkdOC9cFNTv0XYm0Os3xTWESkW3yEjbnviHJfeId/Y
gEn7BSKqjiap7NYGEVStdY+iTfm/ho/WFD10o5fJYHTu4R4RtR8mZwxHOSMZkt6v2KdUQ3cMUVwl
IETPDlgv+eiUg4pj3nIFbgX+IqMLe06DNlDpar+Zxp7NMoL/dC+KMMjPGYazJhaO4DNjfWs32o/5
KXNRoYio5DbxXpPyDhEsq9/P+XfynkksG1zTWco1FAe/IO1JXK/FBAXaaAT/0NnEUqOr/NMeDkUv
SG/hjh2jWaywHlW7/v+3m4fd5H94h9uxH+ODUg+IgkbDJ9fzy8aj37vjz93ZUCKGPRnCU6C2KMDc
9cMP7ty0qA6tC5decvunBWlFQYdnkjSnVeBaU+jiMpGEtwflFDnSYyEXdPJB16H00uG6KdJmZUky
SVztLqym1ikEdXFYmvNw2sV7d0Hh+zivkKla2fyU1puMplB2qQQCbVYo23DOwMccn6wZHf0hAwqK
4VJZJStJmEbnkXruWu19iVfNsnztzFWzlQuE48pjTKLslqGRHtfXoqfr/4jh7fm+uUkHjhWcvHsc
NSQDlMqGMxupWdjWRgsRXHrvbqZlB2wBlMM6ps3AasLvZtbZBF5+RVUECHp5tzDpTE2QtA6/qFw3
ckoYcEDVvJk8x8ksPuzVzugRg1b/JPSJ0xQYdK3FmtV1RbTrvPBAiyf1gkL0JeuBcQdss7Ry2zo7
zeAS46adtf8VpUdgglMmgc4R231RCkL070JiEY1cwxoaq8bub7VT7+XlRFWaeVoFvB9rlvpeug78
wjVrfq3Dgn+guzvfpBBPFNYQCgfelz0+F5fjZoDukGjwTFQv0zPTUdBFWQG1zATJMcPQSWZ+gPH/
U9XG/8Ma4RZpvLOZGufYtswgq3RXPbuwgU3Wgsx7PYNPYAyusSZ2qdRLrbwP6SUjWoXbZ1qrvoyB
M0PV2uKhReRfmJXBJKXLhL+XyijMurabAITZFF9d/FaHtIb47chUHtmvkYqztpSnqnkG4XnMVdw+
f7bUJsh3QNxnCPlS8N4ptA4e8i/5BQr7O8QISX5d9sPbIWQLap95HHgT2+KyeanvZGeN2cO9zjqm
gfsUYo/mYtkmMWtYIpd/uVfWOMveYS/8r8kk36BiK2CMYKm86DDGo7ieE9VIB2cy2qH1qxOxiuM8
IosWxnjN1vRKcmPtQ9Kw/Saxw9c74TVvPR1X4nFC2bb6VOaBQ+1q24gLrUebnYRMGNQnzKXlNpxP
UPc980nD7nTf56KDI3DJCKQ7ZoNYfssby0qMRWSdI9cLd58Ib2KndLwZ/p3Dd9KzamWDT7El/iKW
hxL2J0OTVeZq5hGW/NiRK5dccvvpVdDGk+11+jdQ9Yz/1g8hxRLbwLotYJ/x5FJW2uiYGHmnykFF
xMhhfu265L6yxVTpr7I3aIL3DaWnorz/enVMJv69jthv9lD0qRtohO2dBrITGJyqkamOiT5AiTdz
NemTE43cy9h6QltWkPUBCEFVHTudX8g3h/SU9BWrLZm6Yvpng2gg6xnENFZ/oWXxS37PMrUN/eRn
S/XXR6XrxizX8ZZjB9bBfOQMXoRlkvmevqQq9KcXBSUfffd0O3QoYQhEeR2h74qoKG80jQRV8i2T
MZCU3Z2Dnt5Gcqsj7lvBoWHtpFrZf0viyINgjXXwfX9Ri9noq3DvwnyhQdGOcR8OL+k0gb0/ZCZ1
pbRJbUQuzA+KCtQc6/2Hwc2rKN3t+1pvU9B8iObaU1iFwt3iJCHt7hS3VgsSA6SopxanFy7/Ski6
sqsIyIFRFpiOJsWdRbTsL3Ll5DErJnDbMAEKho0oGtvyknBUVRelK/wiPSLoWz3y5jpDXW4j1y0F
sbvgVBLjpJuXpODQj40Lq9tAU7aU19OgGFVh8UTpdRe60pFT2pegwbGIDbc6/ya0zwsWmOiilA75
GxdrDtg9arzuEjxY7cuegh45SHdDF1v0R2pGYyGMEbGkyjnh5tK9tHrNAECJanvASebeJYlnZ2kW
QTBfAeSp6JJF7HUup59IOLQnbUJDFG4RcJghIkuT/kdYbrPgnREqz2Awy/hvDvjbMrR/NwAJJoL4
c+p9OON5nn7um6yJS77WwWHivXqVO4gxUcsOY4uReb1angl5UDMe6qg/2xYTGgTrXAqiGJkThWaY
NeIHkac/Wj/UbHJB5ycxLTbCBapUvo1YLYpK9m412K5ISekiZHydFFF6um+qKUdR3My0ik+SklYO
/sOr2KNDWi5BwsMikCNjsaMKpqn56ajvh/JO5gEZ58v6gwcOtgz+TodpkEGnVoNw8X0yfPJ8XqLO
fK4mOtzK3r99XgKj6P92PRZixVYu8O2VGqH+ui4l6DhbZ2O1XjsmQk3Z80d6+rOBU/Khu7azPifq
6jUwfXmqCoH2IbYpExG+fQtEph5JmSx2ntq919vYLY13gwuHDOEzAyp8bc1W6DVAXAWgFujw5R0U
WNKYdpWT78j3hbqqahhl5sN1o9rwC6KvmnyefO/r5Mw9UbssKm9wNr6Xkd1Fuwch3tPEh6ZzD0WP
w6+u/DuqBW8xyYtXyJ1cfNvmHtNAaVVtzcLgRcrYRnhnde0qPya0Fj4GvzwaYWklmS56EvmEOaky
HiaVrLRL/n5uRKlR8qYu567luUkG6kIfiXRJ+y+hh2+ak9CSmGUzWy7Q1+nikQEDfcDSzCb0PuOH
CEv9lFD9HE5GWXXhLAiyvdjuWWxDIIBhDzr277OXk6bdwlQ7nAITQM+srzvWHvOeockazCC2fm59
RVhi6rS0VKgdKs/F5D2zNHI6mPDQU91cU2aT4RBoGVfSQ1OB6yTG0Nt7VjyP68II/VLkVjpmyq5D
8Adh/BVZBBk7gVNAqUn/P91yUR8DcWIv3fsKIRyg1/TOKsuYXy5jFxKXKChuy4FMoGhVfZBJHxgC
l1Ql6VaB7M/jZPkrOUXslRyUs0mCnKh3CZTEkNdDRZtbtbglwLubOf9oGCiQpBy6kV9xVuHlCWkw
gYMSwxI/ldaZP0cbomPzW2mwrM9o27TIThVF60B3ulEsRZS+TVp09e9AnLjBM/Yhpf1jxtnBAfYJ
DbzME6JY2Yr/yM23iAk93RvbjT/p1mhbyl3Pz2LF6Lv281gwgZ6eGeI47RzJiRDOb9R2bKTXg1pV
SKThrNz3iILnu39cmmZu1OMcWrLWjsEbJWHosc6mJx7MFCZe1NkxA42iAER2iMu1JBed0CzimTlC
cDiPZJqlqzksaLVL95h2jLU5/fxD/8NgTOiKo3h2dAse5uWSqJgKwZbC0B699FX2Z6/MdQqKNa51
7yySJY2v2hBM86CnMIOTjT4YRLDGFOI+PRJw8Tu11WfzwhmOFx54O8KzV9WKjryzzJwr32ss6cPm
ZdkCCuDMLyHXRqswg0+qdFMe8FF7V9HYHBG+St5u+J8SlsVGGYLVA02bjaVYYhzCVJdi9JipwxCB
0TiH4mqw3zEwbfIc1d5d9gAfrJCOmloyuCr5YjQuYYjVI6F3aZo1uv3hR/GVqfsz6l2tz3hCR62K
F7Ts5icR2IQ2IuOq+N7K1DQJsVr+46euxOf5SU9CIIgTarGcA4IOsebK2ULb6/75UdchZrG54+Y7
AAuGCkMdg5UjTaPEmSvdSLi+mdAUvnGQCx40UetivnsLPcEeH4q+9KEUsQ40Fc1mIZrUBkLfGtr9
FTC9DRYdfQYIPmGZ2PdCuSGXlIbL6np0R9k/xMWe+6oU10jOYWGAiP7g9hdqxZ/gMRDXsTfw+qlZ
2vK3G+aHW62FUDCLSrVRZlrccj4YUbsItFLiQh/Aa1b+l6QPeVLTF0pAiWI/+1iqpLc4z+VsUaXK
uqdsQveZYleEvKGVJAgCTyOOhojAFA+m5Kru9vLjae6dJlU6EtZbakjxY3gP16/pd0MC6S4GB7Nx
FRRUlDe3YrsagKJMgZ2C8wIygOvSMuHGw/wjbAioF9CYbERCaQojuwSubqeHdV+sLNIgkdug1xV8
wU49I1rpVoIZy6U6zchVAnzsI18eOISV+B7i0iBw9PB36M+2yWNBXfjhiNMj+X1Bwcw2NbpaI4PJ
gLo0n7iKGFtASDQ3Yg384p9pxxFCSFYox9UebKo368jDQUADGrJyYr9aW+F2WtGsASPGl1T5rVZR
HRrrKm/mn3MJbYeJK0SXnBv1L66KBbxFeKPEUmBt1PRKeYoDte6S3juZAF/V7v6FVt2+CGlck4y1
ac0bWjSG1ibHCA0aq7J8wRmkgvGBf8yXaFqr7dgy3ckIaL0qzF79Oz5a2EXU6zMR5bMQgPvOXGuk
D5uKxiu6bRM5/tg3B1Vp57hjxtg8Gsza9G2J3yseRtxx79kQgSeSxpXgRSJguD405GjLH135bwvb
GRJED2uBHmUzM2XydYziPPtRgFCu4dErb5n3u5YTWUvmWvItk/ZzN7tccwEbP05Znzo73YErSt47
zhDjbcOBl+77pQ1IPB/3qxrThAIDa5ODmdT4rDW67UkOMnNrjnBCughEcZE2HeOLiBWQiXgsoKYx
zmb7mZjVyhOJlMt9ke4mW2HC/830R+XnjUGe/1H6fOOgvRXNtaRHYoPDOtCxB/Fb6pY0Bu74GQZM
BRMxHQ8OmFPNg64+QOTjgodWLQGy9O6sJAPrjM6kpvsNeAz6nnzzBEu1fIZvPTCirVi5Cy3q2WpA
Q5vfy2FSGcTTINIHND+HOf3KOtHcJir3fmVpx/VJhCBfzNLcy7CJmpBcy0oOUzD0VI/1PeTlbgPS
lS9kuKf0++YIRYSsZEyU465hJlcuOMX5WQc1MjxyxQuFTorqMWAPF4xJOFYNEgju0nHaxE+/7OlB
JSGtg0Za9Wi1A1dFJ0lDD4RETiA8F7hf9NxIIYoDLWEa4QNtYzo7b0Up06cSxuXTYlLvlJL1SmJk
jLwbxEKjB2aWa19mABJ4HozPgbR4ePYg8WU/VXzzbZGC5Zh78AHMG2vFPShk9U6LlsgJA4O5mOMV
xfHE51Psjqz4LRgKOJ5U9Wm+sK2SUzRFS/hNu23Bh5tVSeh6FdjSrY82itIBhGXdOw6KDTz2718f
vwf7XnfybVw1V7gVJKCqQjnZTg5GW9RICR0QCmefY6iDkDL1AuGRBPXULLXmCm3QG2U75hMYbXZG
RB8z5Kxo/hmOyRtPyCNRBAKBOCWwc+rQKGC4XwMp4v6IBeLLQmFf0zEiwQUZaMNpbLNZP+mbToMU
4yun9RGr3piwhY6Wk2e+vKxOOM6GVnNcLr5INpZSYitLmXaOD4uldwV6AmfAu8Xcy3Jdc64DP/0Q
Am612uDXtjmwxfpfah+JScCu1GOmzKaoFNAva08uR3q/jwRUcixLcoE57EKNzxf+FNlnmkSBXfmG
EwL6CuBq2wF+euBOitZ6rrgLr67cmLsaaVT/f1L3j9yGHO0m9Hht8maiM28g0mPjOUbk7MemAW0r
IBNdqbUw31FBF+WHX/th5uW5D8/PjMFso64PT+2ZasjbsFJ/A6IUC9uWcyPsSs60vkb8qq8CH8Mw
MsNc7HnzT43rrQSisyesObVQZvWbfvFQzP+JWCWzaLOGn/JZWR7bVFp7FHF/R3tFzBqmUIbj0eZ9
Ze0JgIbuUJPc1n3u3IKN0i+tKf3LGxhBMPFwcShtrOkpl6Uef5NeSqaeoimAAf/+pF9fR3EjSUk9
2EFj/3670had2NUbMv+BZ5eVApUqYmMEnteCshn/E4eP7SqwtkRVjVqj6ZsChPwiF9Oq+TN+KkGR
oL3yGgtqBjKLvkxpptsLmy3v6rYfNd3KLnH3J7P5Yl9eBYuHSRVw8bhCCzLdKOvhLMNg16d8HSC1
8pJSUlw2DR5L2Qivg1zMcIEgzI5AvGxPmFmsOUB6rhic+RBXUJf32l2o2gEFOXWaf3ITq2J4kO5L
kWeD3kUc4gaF3LitsvVWK4URiBYj45Aqiq5oTLvsa7cWsavH2g85qwO17e5S2lXZpUZkfz+MBEpS
RbCbGtDu0T6zBtTv3yKPAiyd6YFprn8RmLGEO1iVJFfchoshrmoQkT7cl6wjPyCmUjzjvBP3scpE
XYkZ/M1Ns6Yj6WbhSTm/O7nJklzZO4Dct15f9wey7XJ2QbG3BarGgrVHCvoxvlBMLGfg0YHfUR6t
UrzFvr6nJ5xmAghrsPkEXePAPVDkd/IE3VweGaj7OIK2abU0meAl+fhpvhbJci+NshFIc5dV1cvL
J3BxDYsIgx6DIO3qocWrOKCjZB3jKpYt5II1HFqNf8GYWK9Rrgqjr3I+CkWe13RgGIj/ebg2ZHTk
ZVhkApg4Zj0swGIUuYyVpbUG0Sywe0iqwsy4pD+oZifPlQ4coUZKGzsnNjEcEP1kOhUWXFB+VhR9
9oxoTZNYcNSlLwOpRzeF/3W9gHxIXksnODDetXUWIknqKI5afI1rhWaQoIfl56cmCXHwIMiXysMr
K9ghQ2w28VN4QOph7sL6JHiu3otRChOygslLAU5BlgicTSiQisVqtpPfovPfE/GBujkvegjYtD1k
dQV8nN8snijher37//pPF9yTu2QEu/HxG4g1+mNy4jqUFAVUR6V97xTB+mlmf+Nyfiu5wZOEAoj+
IcvuG/nTKH1f5AtFYFTX4OB7httAYyuJ6i7uslzwx6dhmrtHkS7/UHJi2p8LgRtowsFRBFYGL6hw
4CoeKIO/R0ato9qcfcbND3dpYo/3/vgE2Trhv1l7T5LkfjrsbgFWtAYMbOV3ZYdmYDa1AkSdCRrU
2Ct1f2ptd6fykt0JirastMb9XV0Z4G5GBfsDs9LzK6s15tWNFep5CkothPZgN92sxBNV6hmoXdnm
T9bv9AfBGEsffD2O1BD4griqk8Sjr6Iv8WTJnoE+ZkVUPSQjTGUqPV9NltOp6dgbguFT8kyeegeA
AEZJLA57xhuqqgipREXwrI5aMpeW76/HQHS5we8xkfLMS/6W9ngeC7QecwxUd7JeUUPD7ZZNUGYx
3ANWvUArag/NBCJpMoPExHvSE0sHsSsgDFPYLna0QNZY6sRLv47Q8upFmDc2NyC+Qp9kU7HGRGcs
oHrF7kDaESvFCL2+zFnqmLdAMwvcmHhQWobyrqSXZxm5eXi7qwTMeEb++cdtVUPMNGNitW5NQL/q
xBRYqYZ9QJu6CwLt3Y7oI7p5j5jjyTuauPllh/rTcgzmUqrJD9FIRed1OJBfbYD6kb3To/E6AgZk
O0vY7th2zs1O5pVzAks0xTIcQDoCBZL+a1x1IrfysZbLZsXaL/Ekpv49wo3PQiafqepSSLzQneld
Z32NdK/tEAzeM4lMipcSWRy56BsbfajSG4a+bbCqOoCJPCCryTbSWsvV1Zt+tbpF9z6miqFAhHZX
/2QQrI9myrSycearifGtHgE6fFZCoQZADsedFBvm6U9fcrGnJIkK2JXnABCz8f7ezArDE45zsD5U
o4Fso+gYgpqBkDFyuTGrPU4r7R303Xr3L336VXeljjbklG8Opm2hNJyDvVT6mcSbg/I29iEBvSlO
L0M887u3UEGbBsvkk7QsgAt1/fBNDw9ewJhErEOH+MR2lPsjozcnQFuwk8qpDD8Pg+eUYczEq+0d
bVCrxnSoDURtWxn4aiDyImnlndo7vzaFD2UxyYHj2UYrrHGy+rcrH2RDkS1ygww2CkSQ6BkiPdLW
9A7sNwd0zYlda0O9bT5omBAfdvcJuKi/gNz4uh3ibjppQ+4PBIqGJhkwJR25GDGJmhrtARmQ5fTo
Tf76w6iS7Q8NvoOlvOnj2rmSowYjOaxa8Ed5aswZIYHdbKXgAE83V2nKcgu+kr9Sg19gZ3hrYk+C
uADDzaGodOs1NzLBvMi3ld4KxF2x6YsbTPmQj9rAeJUapVJilbDwMMVkTH74/ebp6anZMiAcLIaz
Gmm/Ai+iN6naNC0GFFL/NxIOEQrP2yGbhojJxN3rYlrUaiqKA+Brvds3mZPeDaj4+7nKlHHA5B0z
qjOhhmSjrSAqoLFWn4BQmlpDbD6wSNkE7m70y/E2Dg65YdHj6ck5s6Sj/yPZ3MANUqlVIQQ2Am2W
eQZY32eJonS7BdEVaGxJZxtfEYTTF+b+hDMF8lhpOOU2O5kTb7dqwzSBfkT2TJIoh9N1DVFvivPV
qiARswsyM7Gq1zBru6qC9LvSJzOqq45bSMurKtvDAuudx5XfVHa7weLTWxWj/e6YJJdDeHN7jSVw
2glipa77PvYZDCGrilzqzUNo3mt72dFTfN2PGGQhZ+6bblOTs8cShFQ0gWeL+Y4tWKgz3HCG9fsm
8gUzc9K37ThQl2jMJoc9d3BOIjfWwqUOyyrtPkSml1EsSIFMHlJ+WgY4PkDmgHOknA37mgNlexWs
/C83KFm/dKBzVsfxT9yaOnOGRWMvyVP0JmYiFEW912iUGnlQyBm+rSTF9yxz5DH0Xekyeg1exLHr
heoulTHemlatLDwWtqiU9ghuwSo7seB2fpCyHIRYSWkutlqBfYrAS1i+8Ym8p2HGVxFPcrP0+s93
hpqwXeoG0CDIepozoitQIlji0SQM72jPPcf5IIhg2oR96C1/g+LJo9z74mQrKuYRmIdILL4tkXrA
ruMvj8UFV3Qj1WTeK1XovveOmvd98DTdxKTxoAFtgbypgf2O/Pjd5ggC1XqI4wZO7YQd2WmqYR3B
GXmQ+XYhKfxTXhhYmzVDGoFo9WuAdgPyxTCnRRyN8RmVOEacjekPwlObjCjgWuqSPfWZVvzZT9Ji
ETTv9iOxomQZha7vM1d86NOEBRI7ygqxjkz+I/B1J/tDxwWdfr0LVS5fjOBFFLlIBsTM6aevOGxp
B4qr1zLoqVV3kvrHdCGZP7x/h8xEXhwg7F2Kqs/HajGM9ebh7y9z6Hl25+OondiX/e87ADBLAP5d
/n05m15qvXEmY7ZqzaUUvSc08i0M9sVObc2ccTj/4uVaJ9hphR8fTG6Ler9IMI58HY30+e1MYuEf
XCyCRUc7vGrv0YlrtXxQ64ijDCmbsJm7/13pUVoGdak70l+r7UDfcIDr91ZwpMA7VsJugIG9p2Re
PReEK/8hjo10S2O/ACEcp//4dVKyNapJq1OuCAZsobI4XY3T63JmxuMm+bSJj8F7OBC+mqhY/qYe
RX+ushdWFMLz2Sdr+8vJvM4GsGwrj3V9xO9pidUGC9pSDMSVQHPYsinfWDl8xqzDbZtEkxlHOyYg
MUA0JuGeVU1lIEkiFY7EOFgGL8vUjt8PTUmyRlmnR4kInxqWxZzl57Ikvia4Q+ws+epAl7t2cc+d
f+Te3S7UClgB26XTFKeTTaDXWfd0mtk7vB0IBmlK47EsLxRDixBU/p374UUjDyJjFaYAXMsywwGV
8OecqJbSIH2V5XSIbeNXDi4F/edZEXCrBybB35+7mirx8JiNXe5wp6nI1Z/rI9PfYoFfMn6g21QK
TubfB+YO9lIsry1mZQ7zZFoOSanoUT2kHI+l5BXkZXvbglHA/3IjOIv2VOs0Ohk7EcWW7wf7AMWl
T2SZL5Z0r3A3GThsfVROcGg8462mm0XjPbPhvJjdAuB9rB3EQsD3knOixjE4T2ITdVSnR2LqsKEP
dzMWGcKcpev3adINeL3+1qGO6BTepqO0rKoJmggeOVstZJnRXZ9DGYx+C1c1RTpL0FO+voMu1en/
qVa21twJFdEAyWtluj09TW7wRsTk3RjLnNIXXEbHJHm7n2HbgreqgdZBi+Wv9j+3q/VvhwZdQQe2
uA6tx4czppMmaTPxHY8xRcDlzXkmwvUcASjHeLraiZW3viLq3lLXq27qGABzzwSDnoNre4ULSlFk
1OAyV6o2BECI9Tk65VuGGsOKfmzhBivB/d4bkTLB1eEyNE8O0iLszQtVn0IIDulBjwmQujt7yEAY
ZdYD3iD8fK6wZ0jyiMpGuntNPAYjMGu9uID46hrVBT2XRKqeQOEM1zEwte584eq7fGaNPFyWcanS
odCVxsBIx0AiyT7IfZ6cZ8V8s9/aGg4c1UzkUV6+h4VN6VHNXJq5V2n7LFEJfb8mbfSmA7wj7IzR
ZKTwy72emYlk4DxbwEdwwkeV5CZ9SyZ7UctVkfQqB8F3UGzkdrxvPRKpWqgW9ZgJuAwJQKWhXIUN
q8fGr3UEesC7iDpKrvaMX8lGOiY1EJM/qdF49begnZAAflHicqgeJTKlMvWwfgVGdFIGxS1OK6HJ
WxVQlcFNIDI9QycjeJpYF3WsN5+IYvxOBe71b/y/llLy2K6JzWynS/pGTfFkuXMoYFgaS2wozx9E
hDoet5e5WvwF0Xzm6bWDNeroJdz+0xBEgYhiq7bMS0HqZPFKzVt4075VYyMZY7kmDYdbr4O99OXQ
Qs6LVIQSgi55HWiE4oDxZHqvt0lnWrS0tT8Mi4iZQViHY99jEpUBBK6zmumNnAQukYx2XyvZch6Z
oS82u3Bvbp+MHvUvbE5a34mYyzJ7xj1Gk3m7L1bGbyslcpf0b9QOf6qlyvCw5D9I1VIcZoJYLxyy
//kDPVam3Om/GBJYbx2+TrLdo9yRsVbPT+hxZmjx9wvuTKfDfjxoTI4Y/T8yFuMaKmVv5R0OWXw4
UTQUbVVvrW8yY76i7MIPw42ZMlmlM1F7ps/YKxX5Lw4eMseRDGqBRl6ftmkY4KYCuM4Q/6jjtua5
l0Iyg5NnbDfqyi6uvXVqrTfp2i8K093MxdNt43LmrZpQ8fQquo1Io91N5qkVeRJ09t29y1EGPQdd
Z7LXyKETnTTuY/PdN01FVBppCIg18UX65kuM6rhMW82u4abCJhj83ScFOLeqgLEr0jG4g4V2tDBw
OlDC4Eb6DpXsq2qW/L913Mq3CO4HIQHmbfF93tYSSU8qdVoA5L5llJlT8xQZ92b7Z3tFzWzdRO5d
GIiTBxf8WqD4hAWMJasBrVzuG0si/A/cO2f0Ft71tk7n/VaOlaIm2k9KEpuKs2vo1NyXR0tTgeWX
YjM6MQEqP70v8iQDyvaRkStDzod3KzLQdH5Ou+Pzqvwc0q3tqpwIOJFF5lsRBYbOrXFaaaB4qggc
b56Y1GfdALNvKfnS1sqYBmzvURuoCgrDol89aVr2SLVVnG4h9YPJhpU4Ni4vlN2jBaQDaVka2zAF
TQlgUx/I1yqGqmlKBs91kvqN6/BemHpqw7Zxw/SOPZlCVZS252BnpZ6Lhql2gZef45JAFO9su0Hp
tKiXSwwNUUZkpbzJiQso7HWwleZbnlwj5YMXwR7YYY6MfXR9AuP4mQnbxiOOyqz5ZpBt+vLeLxM5
HlGQNJjCFcLy6XY94iqVstblrerawyB0YmJXIZUqs0ChmgkFK1+C1gTCKuppkUEDXhsevj5DsrXg
7jUL5YvRnU/6YC9bVoQht6VixL+U1IPhX3swo+cyqcXA6MCp4FUq/pHT4jHvp/betoDNRHJAc2dJ
W3Nozpn8VrHXYrRwNMaxyOL6L/0U1fT9RKDSXCDxDkO3jlb3dDnMoTU9jQ6bGqkfGnHb7dj1nU9t
qw8kOYN3St7mdxh0oJW5sQLUqT2ud6dcXPTvFpwzQTl84bE7pix6yRhr73HFzegtq9f1yx98cWd1
ug5Wrypsd0fiTgj1wb7hWMuUnvfgphhSbncc2KMtsOjflFdKlXmjtoslHd4fpxRMb/atabW6j0/1
bi9iVP/xA5eikuupKbzzX0GeG4zGRYhRAIEGXVQLTtDbqf9YASdmN5nDC69RfpAfhi9/b+/QLVqY
vG4DqPc2y3v2smUQJJZT0XVAan5qIqm+uHQ53HIiLvjyaek44mQPvF+46L15MpDqUHTwQE+d2RS0
jAS36CMhBSH+A4PX2PXjkJ6IFRVlEKqV9XExltF+/V14JCsNLrruq2v8JoewFwUil35vyCYH4unM
POzKwrdmOx6BkwHeFW22RI5ugqzU4hjAcqoRgKDFh68ZX+zh7M/0rJYtGMwPFPWzFkG0d3Q6Ohug
IM/fy/JeA1YXVumTA9JKxme95nUPGXDbzZHl1zhBZ6jTNxbCq75Gzkb3rIER9jQfl7zu20JFCv3l
klfunSWs+oPw/npLH2UfHRZXXnF9InL1vRVbet/fpGISXag8BC89RaoqZspsu8PI++SEEQoli3og
lzFi7RFvAG6nMr+nR9sEC6NZYh/v0mgjr0QVEhIJ6aCn41zgeCFTuitMCJuaak/rJnXEhNkkZoW3
ef81XcJEtHuCck4uhM0zqdfw+0RMh8dFweXjges6CE79Ysem6bZZoGGcnCsfGHaKDQDxnsXQlVT6
VAG41Fs5i0cnsSgvpi3xuGqEcGogqKreits3lj5SRenDD6GrQIWwXreccKtiFRVNls74KF65yxho
+U9Cx4ZgCAG81tr+gk4eQzpcFu9FhR4ga91qHG9hwqu6T+zJPD3QzoWQDlBgNb0XsjLY2IkmGBmn
dWp91SLX6Z3X6oDY3GRFEdXRM0IuIFNXvRw98s1M/sHV3gkLWWKPdSblk8rJJrQzYqHDovSX2615
2qRl5ZWhVc63g9XuemDk1xTf09+2sjYdBjFdSED6n9PY0lFSoHN+iWMz+b19Y/ca77mM0qxiBPq6
fmm/Q0bHJ9Oix+Kzex+NS2n5XIZMFHaaagY9+nPThO+gjtOdWsCjohEQq/bPwyrRj0z2cEqzYxS0
d7dKS4A+Q1BzRbpk9yhNKjEruRFo2d4y/m4CtIDKhXxFeFNpdJ4W60xF/tTi8F1dUdItFu0GHSPn
dN10sz4NVa8bEkd1CgdUowvHvTMlYbTzA714JQRVYyg9PNzIAOsK/4pIK5/OD4OSQNfaq3iHqSjK
SWGPDniUiK/PIS0KqzFSJE1nqDNBESYKm2ALZ50ppPeKPitnERfZ5zBYJlHEE8oEx2537N04FT/1
hu6uXcTEjh/40sRhpf37DXLcGT/9clP/tLnlvOmE/n10/7MHBhDzWFlK5YoPIJFU862QIgmzoI84
s7QPtrdSTDAxSkSjusVRCYfa97nWciu8/Ge437k3/d0wYPKWyJtTlu15N8CqAARfx/uk1TmB5ETq
w+nZq6XVSozvRMRg0o38NRzNY6gkvjI1qUAEBY8upJoXTD+RTecAlv8f9Lq1H82PSJm5nEvQmCpb
Vfva/fid5JuIlFHco6nimMY9uwCjlwD5iVmNp/82e8NbTmw9g70U6HEjgj6MDFh9hcIJtqG96IuI
9Zt0PwXHL7vCAlQpi9uMMHQjTseQFaGI4+LJu9jLrHhAm7R5HObUR6UaS0TaKbb6XiEullaZ0E+V
bEPT0Rqv/tUdtq8jH+JdiBNA+jJWwwp20VH9O43r62b8wMhzB/hW6HuhQMvMGzqBghXV77ztt3o3
ntuA+06ogaVEGD4qKxmOGNVICAXmrTFkKccYkWUEMrbPBoeGv/gLQ8jcgSGpdq0vxh4OBQ1lioeL
1M9oN2+COFVjkPCSrI8bk3ximDaxKW/9e+QS/xPoOn7ljAUtYzs6kZzQL2gDMxIrETcOvHYVciCh
jBveQonHk3JW2mNr0W/F0xPVYh7NhSv+JYAdkLzse6rZbNw1yTM5WyWH38nMW0AxCXmlZivrQNor
712U3nVRFQJO4um0/RPwFsyVM1nike1dKBsCW7XLoWmwKCJHLckLNBybnuc1VeW2qz0MzoVKkf/4
k1w3mryrZCGuJX1weA62CG3EpO0V3c08q59UcIdbgvHrdxIh1e+JGPH+gvwGxDmcyb+wOaUxIam0
tiLivYoqu+8mgiTMVv9smB3DjX9sa9hL9l+5wthQi+nX7jemZAnuM8LHPoQ280Mc45pYhqw3r5si
qT/zw5LFJNXj+UbUpQr6NmsAea/2znDulnwDDCYXnQXOfRXDQoahVS/RONRwOyMrzF6n7qkAmCbc
k1TcK2UzsTYAZ8ktz5tDnI24hgzAaDXeLehgWiWgLFADQQ5BoioPcxUQCU5PZ1JsNiDGXEosP+J9
rIQ6IGSOjncYCdyUNPnZYm6w4Kf5cpL88mTiRhUjTOxEMB+DsXy5bGS6q22ihhChTAgEA6EhOmvn
eNpKdHhgc6M1klvpa2lxTlwjLsozIC+wLLLOcNQBV+VwWD2CXm13gfbizBdkNtsLqA+yCoKJhyO5
7mbL1nyj9eLc684+P57J0si5bWo1OewPZlODavVr1GP3KqNIlEWXdBlYl1lBOF+zNQeXE7bRGjeh
BmyGIQ3RNXsnqlujywM17I5sbAv27+EBxy7L3ClFvZwhJdiRrHFRX2vVXzvbQAe2JR+P3wtobtyT
sdFJvRmgcKU8fjKj0KhJLvAo2CTqI8fRQg4acaaoQbayQ2ujuowgL1Y2gFYDcLMu/1Y1VtnQzFd7
yVsWggBQoqtCPzaabG938VU0eQ6B2Q7PzsSEvsCl/4WBZxY5gPTvCnjKHrsVkwKPuUUS1CIFtOJy
geMfyBeluIlnEPXATL8cH4u45J4O3CIJ0jQf897OD7PT8gK9WhgHKWxdnOFCdQN0xlgCBpVRydV8
jkxCfzy9JXG1MaPpr570nNZOaD+m+/Bxn4/2fDHYws6Vv6JQDESawPrsh7RmD4JbuKEzgtE9+Dm6
BiTHkO/QzCVd5ssFxn4ISPe42zuU/EH9Fg6+zf89NA9FyHTqhqUNVTHC4lXV+Vt5d6Vlx62ZMZdU
indKyIezsmdajkQnplFjbfYIPXhNKL4FKPPhmVY4BcUR+qw6ev5rF4hdkZlUfPgOYIokRuyM2zSu
NvXB/RIjMVPV6iIfqMoAVXuhWc2paS+yh/K6XelCVwosCl1uQTlkeV/6tF1Ga77bzBfI11zHCrPn
AsbNI/jkw83llnHmIjQC1Z5EvoaYZpubaStdyyx4rWeu3cGitoeL/r6hmiPdz2BRVkOmr33kef91
LxtJjb0V+TnwDKG0OwpC/DCfrFLAOoairJNGeftudj5uTHZ8qI7K9ajC27jtWpHonfov5gntMsD2
LaeEtBlrjJye/T/6ZHi9yXqZX/wxLiFVNR+NHjm4/k0eNtd2nDVjmjkLe4pVJ/EfPdBlV/CxmF4e
bvvM+UsqsFjlZ1dd0Dcodr5VxUApnaJl/TLMYBr8J8XMcmj9T4/6mLIFSaFDhcGSDQj++D99FPpo
uRD9C4DNBhhyqGf7s1akN2yFEZtm20O+b0VccC99uHgNLgs3RqYHoBfpUDMfYGUuicIRA9lh8TWH
eA+wYZGBTL3GYKuPlLYOLeMX3BZOEsTcoUdS0sk41nfV22NMJ7T/CKoGJemSacfCR4KUtZo+ZFql
qXCRWHFBA7C1mJp16hCt19uGDDh8KP83mZm5RIXvifxjxz5xATt7YL+rvztqzQZKOfdna/8IbKe9
8S7IrwXk0qHxlRxFwWDrrQBTFQbyj2N76QQjodtdtnUykshJNOg+ag8Tsr0Zo4ZEej0wbzM5xT/S
iZwurp1QoglMX8yuOXAmstdqxU70OO2wh4AqJiykMSmbE+5auYoqZKUElXv0+qxuV2X30Gv/Q6xq
f+U5Fbn0bVlUagtStM6Z3TOBoEHdmXeqviNMaf9w34ALqLlkJDxBkJDz2GO8EMSj8jYAxXgZ0ZXj
28nE0LFmgqwANfw4AX8jn4n2M01WSB+MBEp+XqUaAzBTgSMIFT1DqUbjeAaujIFzsK/LX6ggIGZ9
YeGC9vF87NpHzJ5A66q7C0H6ZamwjXAKR8EzG/wg0vVSLcDEGzb/KfH3kC1KmOsqR71rwGO7eGWe
bDyJSOAt/1kpO9VG26MsYIJZzhoO/vGK2y3DqQ6avCHtKbk2U1U96FK86CeHD8HEvMtcaRfyBF1A
9XRqi82HjgU7H9fslfL4h20LFn94Ll3Qh0d1DPqtyxfFKd547gQ+HG4Mf1yawx2rTq5h5grKt1qs
UmaDIrDyfJH8aC5LtfzAJhmCpXWCMnGTBadg4uIbziB+/rK6VINojOQQAykII2SYtMWGNs3JJ9Ej
tb/kVO1m5qUiTGbxGxG6tw++g3WE0N2iuj+flqxvr3uDgSzUbhMslOLXUVz1teSjgvSsOZw0EQD/
302thyMgXXKQzAW9aBe0yE3mLhi6crLN64wJweTREeXd3RPQscSV/GxX0iS9/6Dv12QWJ2vL5R2a
wgqsYEJkyx4jG8jbJ6fihJnkO//4J5I4VvWpRqvDgJ7qjctiez6Ya4zwWCKuU9zqdGjeda4RKlyz
+0cdIzAfB3SKUbOv75qxTeIoPTGenKF99o3ihf+mYoRYDNj4nq4bE+4eDxc1RIZot/OJfTYjtmzG
eE7ZCndWWuTSdOSqGDMj78sNOxNuGSyYN5dyPpq8l8u0FXJgxp3GWML6acBm51BPbc2vKWu+Lt9U
l4GJIYVm58XvjrkZptk1phDAeqEbSyWcrDsp8X75tv3GRbA5yhvYxCbft6xJguaAnPb3KNDURAkK
9WvUjYFk7QOqM/3SJhgfGDYycQYr7ZXMr1hZ68M9HZphxpgywvUN9WDZxyiE0EWOCKFxqhU0ChAb
FxT+zXlJoSpeO2jnFN3/bDVe1xwQGoJj6OJlj7KpnPGEJ9STsXj53maivMPJxwE7XIn3NiBe8BdI
5szc7N9Co5AagoaCsRQ7MG8sgM4y47emPbDNX5obCvyy9+mp2+D3MZNPK+gKrVjLgpyD85hdsIzN
ekcKt/O30MXP6UPY5ew/+0n1Wyo8OE5MmhpZ9Y1Z0GBEBBH9EaZmGUnv3I6DZxUQXsXJYXBCnWqh
KX7zfZgmzLkJRF0PguA1oL9la3em/jSI+CosxHJ9LK6yPvazyM7mnYU+viQnv95g+YpxfIg/hGuo
6EyWX6iK0wbkoiffs+vZNmkwxrvnIqKAv1a0Hz9N5VPtW5o3tl14btdlHcat/AvYEfqcWGcRUQry
CSe01r/H5kOoEljSkyZHCDKK/RZrCIa05KNMn4c1W1q09wwVCgTCF7fTJO/lXF4lcABhI4dWdd/Y
xdUKsZvGxR7SadmIuTuAT//VjLXAHzGasIh1ychCQO4WaxErt6zI6oCTKKai6TtIZe458lmkCdqO
CShaSpvcGIINrwhD7+GCLwLzOfDAq9TAfZZtj+rq8PiL1HO4E1LP0WG39p8C3vsNL2rW7clSOm0g
KkAAhT5ix+6fFilNYz3jk+RK0BvXw6IBI4DIqSK+EqeYe7qlBp+KdIBp83GT3UnFV4o7lQHE6oDl
05U2WEwrGZkrsHCKB1eKVeFi8bl3Jsu/40934jmFVfRS2UsGJ7S6eWZwIZVhrVgTn1dsPe44DWCr
9iFykj09zDDdyQLOxU8FbwYQlTgmZmARdCQ1Hh6e1zyKSJ6HDuD7w9JhZ746w/5DIoyb0ZkxUph+
RY0HD5HmUiGfW9Rxomi5I7ez6L5K3EcAmLxMlJUwmRVPERBI8YsSdZ1IqTeyhV5YFRSJKaZ1U+qH
ZQ09Oi1g1BpErRmVgKEoIQiMk3tebZSKhbcvAFVLTSua3XhUwayz8SyvHARXxZbXGjgbz8pExghg
fvsPwFvWffrtB4rxqk2yhJZtotmdntcTqaK2dnzop8TNmMjBA7lJCwqrjeEnkB2bEUfwwkhYbt6k
XmDTap9qf+vV7cJCyT9JNmuqLDSSqpEDj0cH5Yi1B3LQpK2Msdwyhe2R89vN1NcAoaAcaYXYwRxe
HsGcrN1le9dxwBnmg+awVkQy6dgvL/dRc2dpxU6pEcXSYNZDbB5F+PsseJvyj3VTkj/0P06pzH+G
crv005lg2GE5YAqLsaHCJ1EA6ixDRib9VWOSo4uzVIOtNnBIb4s5IFB13rBT6WOJlPrB/ddJJPsY
K9EyhuaA2o/7xLic1BLuf3+zXDdN/WdiibtHIRISzANt0mB8lhQJ5kMoX1VxLQ2kSCgkVsH6sp7F
JnkndIILeAo4Wld9UHdObfJIoWoE9Hx3DTHKQrseqqTTokmTcdiCyY5p9xfijfwQT+pnbVJnPGeQ
xtD/UII4/Lo1LEy+42SFvVRLCigDz74dm9r32Ilm57Bl8Dyxo5VTDX4jlCsJnE+iom8CSntpRB+q
L3U6d2h5JaNqbxWllGwhzvaehCDUYuuWY917OL+iXeFzGWLFvvGyFKQ4CyWg0LWV/sgky4xTyJzc
zPidPUlvifkFNbSeYyYCfbIjHFaZIqTUMTo+eeV/uCTNCIpXQnyNqCO7dyA7pQXC2AGBysgC+LZl
3BZQLEpombLUfiYQivttKgqHtrz3aZvc37qzJD6ZYzf2j+YPfZOtdbsp31Rh9fVynAimyrI88INc
Wi9/FGuXNQBTLCgCsJzou3wg8g4dJLvP9UVyus8WcUCMmyZTZDCSdqGQ4p4P1d4oRrgpwMeqgCRJ
P87ijbSed6jNT4vhQWwd9nXR8k3nEsogee50zFT4b3dqRSz9uDEiH73+SEXm5QSCAgwkyPVhTdf7
w1uqr9B21JeTkGHy4q4mAvlBvCy+5GtvSlT4DfWmN9jzCt97+cKaMr1qfWRCBDmTk3U2OjgZ+ggD
2gZJrOyE2UouB+RVGjBwmWKnzowoqlalOu5LknbZFvwvl4/1vshwztsecE3wAzWL3D8Df2yezs3Z
sznnttp5xqs9QcvpHbajKQCOUKyOOTjhgJ9fHPX13wDI5Or/+UFAXl6ALTNSEwqMwUSQJ4xrNUfS
5roZHTzbHHR6f7pCJlYRlgLbQNi7pWq8zO6r/474GRc9w9GgcwrLoYRGtlVkvp0XJzO/fhhN3HJh
1PQmUiUe+NCILY3jana8tbzZ/ivvhKOU7dxVIfLeHc2z2yTJHq5FfJKZD++Gv9UjeBAseCVlcuTk
yx2dW7w/Tya8wcJ0vWNIWFzDoXRZZznj1wxqY7vS7VO/ds4YK17/B5DZGCVQrz/+6/OAVTruMAtK
57mT8GeuF6RDE734cHbewhlHxZo0aqaGCH2f+9g3L7mN7zDe3JhajVSXwodDs6iUSbQEMVHqZgld
jo87kiafskMtPEbyW+rOf0PFHD++6B09BzUwa7wwXj+0FV+apZd603STs01nl7Sy82P2lt4zKHjL
hqRfyV6w7JWKtXnP7xGtDjPQqf5Vp+eyKZ+327GD/n6Q8KW/PS5EsAxzsOzmLqFtINDyf6jIN1Fh
vdCEReDAZGU4RaC+RK3WRM+/WuqS5itJtUTkq8UJNshefrtVltlaKfWIgHKxLHF3FCJsfCVRskfs
4MVBhc5Fpl9purgnCLxRZF4iF3LbrtrK4kqTnx8PZV2xEDRh2n85UJaLvmi7mM2ot0YWZH4wflhy
PUayy+PYOxeFJkiWq+yBg3SqngA8iNrGNVhBVWyYbhqjIBJYs14+HtX2L8kil/0gBLEk4wJNFtj/
zyuktvp8Xq092uWP6hoeBYgnvC99+6pI2b/kJxHW+KIOPlQb9JKep7BwNF8A/Icrz22RmEuYu7/J
+MxUPh4deqvbPo//hTqHJUD6MJTemu+P9z6K/joXW8k4N4UqrkYnl2zM9OB2y5lyxSOrUdL+G3Do
miX8EDbNF6GsesdCPkeAN/JyemVhKgXdRUaFHpE7cLAqYPRSW3g9GB0g3KyO02yU2bM74JhnCoXy
iupVP8ZMbU5GeKGdNLEGrFJPoCf8pJCFYqqPRz4d9Ut//jZfBGCeRl+ybJe1BO1D4pUVczcvsZti
REvSf4V6IHVd3p+Ti6bRBCrZ9jUSH5GRJn7ZMn0TQSRaAPOeKaPJCcUdMbikHs7FGZPUCoDU+6Yp
YtZRbGGP3zKY9gE1kB25djGMhiIvTaE3Lfrzg2nlp11BkHQkqad0utGjOQd+cOlj0GQkVX2l/O9v
GpwNmcdfKe7c4XxVhfZEKWia2vullY3Z5LTXPi+/OvLyDf6Jz38n9UoA82cgc11CuMf63I3uRVqn
V0MUcNXc4JbpGbAGJHchDFxXZXgO0+Rr1cXybcPcBWCHHzVt6iv8O06nubnWlg4gRDhGFsfXrnUU
272qzeJyOg73LwQ+r3xnNagpWtWouRJUvgbOx2mFafLWDE4tGb1AOx2mIJ1Tmcn3mgSKE3sjNH8j
vqEzh/Hj2kdsB36K4Kxa6HxNAJ2a+bDJvAi7BS4FVWrRu2wJXP9eU8qumlVjI8hfU28qKULr3Zwp
+hlHQwkkSez6ETG1x6uhH6Xg1Gdbh86i0yZtsqNX++cHiUAPF8oP3nRzTFgjkLpWM8VnS47pmxXC
mXm2OBkErwh9Al/sAKsgmMrSWiFQMsxc+QNXPIhMCGgsjzCDYE1q+GUo10/aLRBtWTVDOVuBBO5P
cks3kqwXvIFwE243MRZk4nHeIxeCn+h2a2BcJnk7rsxX7KGvuwuhlVBD8oAF4TgZNVKhvYNwrsI5
9AhH6SzpaNLein+syusvYA1sM8M7y5Bw70wHrfqloMPm12SIFaOi2wKWU+I6yG2I0l2VpB4aO24o
X5Jtq3NVwsUzc43nE9vHIt5XnD6r/YMX3lRI0W6Ug7aBKU8qMWo96u7860qo/uS0U21l/kQgKKTP
yRjHer/XCKSYqnIdbcKJWtVWvBeGJJJAQtlv5piIoBi9EBNoOMomFRTwMhKo6GzbRalrUqtpwgub
EpHcx1lkd9jI7/1YOWWkcSSVUt9sWD49SlT0skqPDNm+p4P3tnA+JwAeSK9CqUD6pLaUo7OR2jIR
c1vDFvszuz3QPepZZvWfHGFehf20BJ3tWB9OyzXBwCCu3jh7HJn9+wOPY9bnrYbBjvc67j6HK2it
bv1BGM4R8Gl2BUVnfXcGzOUlBKBxDzkIuxvpdoCsx6qO0hRIKB9eZusf/D53U5ri8p6dSklpsARj
ZXM/X87sighYE9F6Na5GvDx0pozLdrtCj9AgVcZLiCRvmuhWVyw0Fa35ZhfW1FmyC3tgReSF3Nb4
j6gFYCkXpwtagV6MK6chaxA1aSE4XMZ3/gR3oMl8m4ky8dn7hZY598BPWrRlQrPReAnqenUOu3hj
tXBUK/AC/y5ygR8EeTb61aGYzeef2GQ1qpTZf6tBNfqVVfsshCPhh8s4UAH1RHgsVQI9uBDTvO74
feDMTN1qvYg817YAjxl2V4W+Uczm9Z7DJNf2nItEYjB7NtCpOFqMe+nJsyc7jOY3dgnqPbqLR7G9
8S/g/iilt5I8R8BXie3AmravMdLkss68KNDOBOP3dTFZzFwj4bd3kVnwiBK1x5U7CUkemqkCoXm6
8GhPUG049EK4/crezeAFNpbi1E/wP03kZCEK8GbofBzeH6UVftvE+p41yoRab6dAjErtqU6iL4Rj
Ocy9NtPnJ3ab6IXonhi3ZbBbapcXPDsmArQoiSakGJ+8VEVjXPcci7KEyVdJaEJebdhH/j1Svhaq
VV4pt6PWOX096w+kI8pG7aB7wwparYsmtXZZMPkagBEDxBM3w0D9JJMl/UGqf8Ud8hPjBhbuVcD9
vDtCTOZUywZLr/+TdR8u/GKjb49VHMmQFQ0O7cwgaoQY7OIMKQ4Qhyz1pdz+c18ohGUuyRrp6KmD
GTEz32P67JQEZUBSQhjPcD8eNQti+qeZDsvxu97nqwDvyla9WHtVsROSybJ9uWIcrSODLcHBNfdi
fWx0f/7O+d3Nw3UIhB+ASP1PdZhoxrjpTZ7RcGCNWqASCKMPGLR2TqmrmZdIhcX6rmO6UtVrq2AD
WJR2wUzhvRk7gV5a+0PP/GSLN7d4+oJDMf/YxnzeG5MEqwdm6/tYSjUdiR1ip1IybTm0LUeih+Td
ypnrZtK8TO2c+upUS4v9bnL8gcbCertp6zpaPOoPkDCFG2ks4QULzr+lQmYE/GZPRrPBEp10veKJ
l9K3coGk63vTHl8am/tJ+eACKj8ckPph8JAb079++zDfjhf/hrhgVhojKDpWRmV7aRlW1wwPSEf2
6j48HrxLEZJvqxlg9bniUvPVoYaqLLlYUZE/WwYvKkfz1sspVSh+I+36g9mlQF/mM7v07ijdtLfT
L9c4Fi7IStKvWayh7x6PQFox99G3IfcGfwhy7HoYydXIPfXTrpiM6FJhq2hBohREBoPm2aF1l4IP
ahA3vVG1cWgYZInZwUK3nOtXTgFJlCBjjNUZoDFvQi75Lf2KjAr9kATw1Y84XgUGDLXLIJc7sI7y
e1Ar7gagEMkqZ7w+zq5BWkJtr7ImCys0b+s3Iur4dyIMkSpDjuIQOpSl6u6s4Ujfvxx9unvA4uGv
g4nes+qjMtH+7BeE6bWq7ATxQzkm4L6mdhQlk28LiS4XrHdq8h7eQCdEVMcahNom1MtPA+GRsSmT
bZCp+pHQxLo47IhAqZwDRjH6QedFC3JvPWIZWz5yzQYM7i0JaBuQASf6gUvAFe8atOtROgVjgJxH
GtnPwYtwjrj2Fc3+3rJ9rENZ6/K3vIxU4utdN+T0hhaQfcvHKuUIsCq2Se2UPGWs3RQTOsKYqPJW
yH23fcLTjb9wUvXpzJTjG9GrdpuQqj5KPlV0VdOejkG2m1qJHnljGOIIiKvzIAS+zEgebiDqCreA
cw+1dROdBCwe4DWgM7nmnUcqkaw8hWZpRkSWno24AmrCGlGz8roYIkFOWefT2t0rwyNY33Yvl7V2
TrjgbY/AZgG9QuZIgSeNa1esogUBrxi6Hqs3+om2IJhcwwyUuDWWnangdHWvN0ir8fFAX5K/Tb1s
9hEga6CXYqNGrtD5m06frjxsUKkmA5Z2/QNBLNP8798kf3aM1vxX0tndyxdd7UQ/dzzePr1Zo9xc
qNXbTYi/94726UcJsVqSbhc1DbT751aDKB5HZwABs0ynH8OvttICJ2N06ygjXmpXKAdM6ZjedC83
Gh9GAsh1tOWh/cojIxu1uq6+8IWg4CI7thYKYl9i4oFYl4TOGExrpdX81gpQAb0Z6S/YLCjKoR5+
p/C77/x7K9o8MlhH6gYO5RG9VvzH+SoukZysrUA5ZBzbyqivbWtZ7AcAnw8xNFWuo9K15GyBTfwK
lMov96vjs5q1yIB9Sk6PoJrMQ0mAg33m5IbZ7eny9JKzyuet8nWF8fe8dRcjnOCXKc6erI7WF4pX
dNabCMLj+npFOaxSSQ1L01UlKf4ZmA3YGsRxZzCRS2IuQ88j3XZxoPsg0pHvnWWpeIwPSNZ5ToFr
ClYRwNDg8yHfj6iwafoUAM8eoMuZzfFz3eH9SAvY05o5xzx+3ewr02D03hj95f8fjLJAeoGomoaa
H9ooe3/HS5+DgdGFia+2SJ6H/vB+HwVitbx2kfUO9ZgiuS3WbHbItusqKMaqdPGbr3JxGpqjRoy+
wPq8rdCt5z38F1olfv15GToEMDUUFbw0/X59h+6eIqFaCe8E3P7nx6ClI0hbzaHrBUis117GM98A
FIuOmuq5JCyCwRqECPe1rt1wU5TjoaILMFBcCWlSED0FbwdAvCrjA2TbCCJAopY4sUyVcg6m9sMI
kJqYWYzhPUZEF1VZHTUhci/TOX+FIZsnzATr87vxJjMXxGqZxlDxP4uQ/V1/qglf538MtuxzeDOW
5xyer88BadPlDCibgwgCgnfjgMNeXMGcH8Lz2gy3PCtHUuj6XgbuU/LJzaNnjrwKHiwqcx+EgGM+
kD2NH2Ck9GgfdV7S5OLjVmeHMlMv/GACeIO/0AAbdKS6yc0W6PODYzA5GQdXRyqpeN9x2JWFhTTW
zhT3h0aSIzKD7Tcs8QDuIAZ2HM3R84L/C/GN1CZNM97x5x4gaKCB0I7HqOW21rM/EsmShGcegicS
i6zziwuzvPWsGU9XtoGEVbF3bdXZiVQbBTaPo6ez0xnhGMW5KNCLGobrA1XbL3WIAN1oVa7JdJup
C8ruGcKHsLu0o9iSvoTu8OgZEeD0HVBXoRSAUC0drxbHyCrezZndf9Qix+TjQlv4+g8cVx1YTqeF
NHHeo2fesOghFiSwNBHKP9F5H2OJGo9BnsNZKD8xJVk1thKTeG/F+mTiN8BKrun+qTXg199MFGNp
uxb5vvt/H0B0rFrhRkEBwp3BucaKeVizTgNhhso3a0yvZWgA6Le7AyW7C9mIfKAECj5dd26OxpOB
PjB8yUWVlRb5cVMU6HUJu0VevO22Ar+oeK2Y06Cr7aRZ1LjyAttfP8fwEJTqJlB8F6T7QL1lFnFM
n9X8qVL1mLizpdGAqgAgFj8DvrZOerwYDRd0A75+tN2BfaZTCpIaAqs6LfCcn8xXn+sAV6ok5hHq
lFPElK1Mn22VRqEmuKPuuTPI6P7McOktz5aVebCZ3hycuuUOlKm6zBdCWEVeWCoEhqfL/dV5YGom
L89HiRB3f9Jo4Oi+3BTnLXHzhNTBTzQbQEc4ctHp2ZjlAD08zn0vfWvI20sTSSQPx6OPb/de1dNK
SIMZsRyGnHHCG4PEC1pP0CZYt65p/zeLgm0r0ZjMM0m7KQKwR9oZylrJYIpzc7qRJspypocAQ9lw
RiYpiQffrZs+S6yeERT+PkZm1mZxQ4KoG0Yv7RYy0+yEysFo5sSXmNibyKep+/nB7YbyD4KpcPi+
Cmg+mUYKTXzumX2ORRzvePfxtfKFnlLExp1ao9MVIJA026M8DWsJsoUAQlEHiiqBkZ36w8kx7+8m
7ToV6A76IPFq5Jlajn0XF6MHDXMXwwnk9V6gx56VgXYfF/cCJpGdzNNM2eaPLUmlleVeXQyHo/QQ
/9wMTvT8o/3qDQZHW4dXN0kT+8TZbE/VH1n4qjN2SMK7fKwxaf0HeXexXyLeGEMQc1+T2l3oa4da
A9tmwVCVdtzSBAwkDJUup9+ywXl5D1Su7NbFJL0+nC46q8hl2W4o+RVCmJ83vlbOytoBoyCTIvu2
A65oeESDaay60pADZSEBFDgkmcsc0y6AadLCVaeoERap12TeRi4lrGVPiNq0X/mCHqFN+ZBR+Yls
HwiqHExcRvlDQVHYs8ZdjWA3xejzpzX5MyQAsXwSl6nJvwL8i1tqaL5iMZLFY/mu9RnV1zry2DB9
uOdycplJhJeOD05h1UTBnTcGr1lTg4UVsZLuZWQcYCPenRZJbdnLOFvUPQJxDk5lg6FD+o+G3hwp
e9NURigx5Z0qT2l+T20UwQiIYQdB+mfRsxz5HVAUpnSu7ozC5gfTCZCbH7kujnulrYkhqlNHUfLp
DzHiczp8JG7xK5EP+dp1yUSq9PIqdDMhj63Clum5NW+iEtSgeqhR8ZI7Hvxx7KngRdAYuh4GPMrN
ubTR8ITWW/Y2hoUZ7WQXW3wJ/FJgZgJCuzXInLlxaUDRXOJX5yhPaf9VKV5bGpPtnRLJdg3P2cry
HzmHydqkHfu49KmNDJajhxCt3Ilz7nxbFXpI+Q6zNdUalhRllA7locpZR7NTxoU+NyBKD4nDSk2e
bSpvzjD+LC5fjQ6Enmv5CBWTu3Q8yOhgjGLmAKhZu7i5JMYIWT0Z5vCOqO2/k6nhz2uPDSuhfACh
ASb6vafVJDIYw2npmqvCdMfqxRl7h1YM+aIWIZqd+nholv3dbmjdR8fReCSLtG6MXWvQDBG4qeEp
+l9rsYlPzNzoz/YkqJYw6ZVInyINvov5Do1SC9v2yzimcJ/uODPZKlLu6YqCQPGTJ2N33k01oOGt
OJC/7oFKixRbLS8e/8BvjRqdGh5J7LMKKpF0mx8K6LU6tHDL9jHmkg59uGRhq3Bkn/E5Khp7c8Nm
Di0RMmfOxl1ihzdZ1yrEPdtHkyFfb2viAJ3N+aUEijK319hAu6ygwB5CMbs/1+vFiMvKGxnTkV5S
jT5oCE0YjMPlwGb9pgm5aw45KAToK60ElnmHC0K7Jz7wt1o+1eovwDdD3gPflPVKEqdWiIdx3Eqa
vfcX8rwGbLLrbNEkvK7cg28pmTAFa4Iqr9nTGaHE5um+JXae5LVTiqvvmog6pFfPCfQ3+AWgiGwK
K3k0l+wZgw5xJ136A+tapgvDhxtawaHIR5cMy9NSqXLr9qYs+b4bCa3HB0WpPjwMCuBDNEjluj0O
x8Y6HtNqBDLVYGFh0doXvPh5vX/fIWZi2FSDr7t3Zm8QdJJa5LFwEjhwujHXGVuTru7DP3K8dD/s
3/xBPQoQKyZpCkJU7LpTlj2na5gl2V4vYwoX+JP3bHxAgCViOyvkm+R5+wOC1tO5h/bup0JquEq2
T0+OhOHr0e457hqfAdJXKaOSBLG6P0DcnAwdDbP2cF5dhr5v779KNuz7COT0Tw245FyhcMnKw1gm
QhLq/NcMdZUeBbSx4RBWshlIgCpBYNQmqeWylmGME0z44gu//+zQAJ53rj0kBf1zeRjqnJ+MxdHm
jpBk2KS74Y3X8e6/MJyfB61uDpV45YjeLoK1Sl4ABm3RMPYqD7DjJCbLJC/YwFaMU9yE7VxKxmdB
XRv7Jq/OQ6S12KKQACTmVE5M5IynZbcQAowTap6m7eM6t1F+IFLy+X7ttTy9dgKgarCf+cmhIaTR
C8A0/ZZW+s3bBpVs3Oeb+xxhkGTD0LquSp3sRd+AOJBVgwrY89susvkGzqpsEr3bIXtRI92py9oU
Wm5I3SLWHtTJJeOqVB/m5GbTiStnDJjl+2qi3E3dIUZoUf7RVwzaoFkF/hNvBiTrGPUQkvzzcKvh
9jxR7LaHoBWg0TZDQNV1FTNww0XAex1xX81bJwRWIaIRdPL3cnBlPf+nFq9lhdM3M13IEHbntHQY
t7fnQFKZT4M+w2q0QH4/Bhk0VfMUwpIFOhm736U+8aaQCuV1qQN0jZ/b+7vwFGJb5gO9toMm4SjQ
oNiiogeRZntwQ4DkQxVLxniL+fTvCi36wwlxaP0v1vo+5yIa7dZuHOn8ocHQOCA/maZWkKt/c9Jw
zVWeQXds4X6+eKV56Vl2tNGz4Wb3S1RvebVzSE+GDfgUktqWeT2LeBViHsguczRQluWKcyicc+YZ
KBGBlCQ+MlyK1eeS+VqOcXEx3cTU1dCBg4N/Ynwd8GFVJtET5CbEWfVAXJTbcnIFGppUzgQyungi
aPYJmOKQQws0Spf1MgPLLbY52KCpUgZGlVBNrMgv8sYMZ0pztEQ9CC7a7cly6xffOBN+bsEjAtkk
nATPSBU5jW5ImtUcvKOCm4Mux5ur8cQGos6Ru1n19rgksR9sTHndni9OXEwjUkgVF4rpNAVrmO/P
pwcLyfjnMVq5cj0SLO4YBIsChF7eg3zC9cTPtSDS3KBQLR7jxJ10sFtxpIlcNTQqts9lDs3WF7Fo
B4Xm1IUPRNKcCfhMPOt2Z+x4iPYahBfsQ6FERiUhzPHxlnMKdJGq2zn4MkUrAXeAvkjl6/2sPTSy
/d2to159c/s7tsPB9wLvEqUEQh+3IeOhOJ8uYIjUzvxexaFjc4bTtA6ChO2M8hcTCiZt5FRWLTd2
12F0dh7yh9+jWpY8evN9FDPqsw0+/0Sfl3Z7ValwrqpZEXJS0pJZvBX56Hb/QzT0HYw1UYbgjxSX
tu6t1etgz1Em9tCS5142J/RyB1WMtYo0AdTqVGlaYaAah/HU6tvZMax+HAP8XhH0dnawViQt4qum
q3HWC7maMn6SAj0DfyL7XumrSr/hCLgnpoH5cAllgJy912HaEBXtLa+1m/rR2ZiZQogFsGIWfbOc
8P/uK+kVoCYzERmBFXxmspqVtOowN3JW/H1wi9Fd6Hqwl4eirNjiXvRPZvvNMz4aXGo9YL97r9vY
kQF0XhszS4waRCnriBRNA3wk4Y7Q8/w7fjhXFBhQClmSSr9z3y5Cmf9q3xahkS67T+lUcs05pJ4F
OMslZSbIp1q26EYM3+ZnSLZ4oGK+Ryz7/o5Ju4QDVXvGy9oHp6x33u0OskxAalRjSAS5ouaAp2gj
jQbrVw5Iih11Q2MGK+NZMA1fzRX2lLmjComPTQVEqoows6k9Qrk7i4k0OsE4Npe8sQkqFl2PYPm1
/4slTmEuWpt0s0YZmBsY2cQf6i3/JobbHxqxzGnPRX8UShe94UgqK/2KAANd16sfG2xVeeZa4nUF
e0jwILmEINRCelCibUIsKCzt1mGOtCy7/1KMa0RdDbB9ZkjVXh69VKu/hRKUbvu0kt/Dk4kVZdpH
OIj6qyWdW5rhDArNOjBdW9MJ22c3w9rW7gggXTybHxi0OVcxuxv+XkPbatqAcrdY0siApkqJXDEm
ORrzYB7MvfTLFA5jU02P45GUBszieEoMY2688JlsxsRRJxp3Uc3mqCnqiapJlgrFggaKHPX4cU10
MlY11H/MYxHlakyE5Xu5woGTy1Ip3BDNyIMknNaOq7nx7UWTThJOhGwNBICX47clbXfdOdpCd+Yr
ZaVhk972+GS1MSVZoIJ1fuf5w12CQUrc9A13gCwO4bfhLjjQRUrkEQzhUfbtfbWrrYLWQAhUhVH0
fToafbDahZt32euCa7/4q+PDlh/YxT5g+fPHZr4MNLOe7VtO5UWyvczCkwrA9udMkZ++Zj1ZqMxH
VxPrxb+0kgald2BhaVQldIIOFUU/hi1dPdT9+haN7ybkq/lXQKJC7NvLffAdEJRC13UPS9Nq+7Tp
Q4VXwtuJIMgi/a0aGC7mHyYBIurYA1MN6fu5qYYZROb+DhhzK4xLFggblDK6gx60c7Z809o18u2/
7ZrMkcl7l3a7+Zy+Y+rZAQ57pjasm4W22Ei1MdN1cuzNCqrJsxk4oVNvrNO4BrJOglMJ7NDlCgSp
bQxZisOdZgU7CdoC7zIwdjwwqDahDA9eUaCLxHGKRzu9VNzP8btd3jDpq/34U+L8g8fIAeh0RyHJ
6IR72s6c6m1QDaCRgcImspZM7+Ap6TTUEWgxif2d3kgdWNurTbJxmCkBO2Da44lpsnNL9ftfRsaZ
pnALVWXvqoZjIKID6yfVYPelekHecRZfdQO12p0yOqJeEgzQhU2lNDRcP9Q0+txVuCeTAWIqlure
qaGjZrMgXrbvq/+1JHaQ5vWBH74DkvR97Ireh7Z3/HH4x4sOk0aSHskVhqn7+CMzBe8pKIY+Fx4O
ZwpZSSpuV4FHKQcSf8cXsxI8pNNO1uXEyY9dRlzc3sP4SSgfqovqvmPw7jfMNZjhiweQ+qXyFtrS
Mo0LzgHYK/BXxAoTFGo+AZGTnyQAR/gE2BaOgkwXk+g04VDfTjjyzaAInYk3608vxasbtK5czsm+
ev10uNFFrJsnYqTQXC6mkK/femZcZCMtiOo+b4gAB1OgB0r6lrRIqsT4nC2XA8Ql8OQG4G6YyGQR
yhVqdFoqL8xi2z9avDwiHOsWx0tkLJaXIiLGJRl/HwqiG343zFFQUP/EPUr+8txR5nCJZWY89oT1
4PpqxZDkTFoQqsM3scBSUuE2/dmguv9/BFg4uGkWTFq/zciyxckubqv4mccoDj2sNaw3f/YB9lVT
jsfANVdgLDMeBV2wTqjYToYpLW5D2ojr/Gp+trlJykirEHIL106Qalwsqa3jDIrWz+TRtFprak0+
Oh7ejMNObYB4aK3WPfiWSES8CVRkzfLHHNN1eqmhveMjShWUbFubPiWfyBhI920u1ELm5Wu21izf
KgPdjlchluqEBty+/N4loXMrHbIC9bSj8/DQdFwlHkUEkaDlKyQaGc38+23rQTKKFCyF4CIxPOzz
89kBjg5SOKetYfzZZEWnhnEPiW6Cs2wx6Emza+pvSyQdVW/d8EZXmn/Ly89PdpLY/5WvR1/eLhtA
TtAWHTJS4J8tqx4FKbBf4ai++uwzGFG6RJGqKxxR+iIcjjRBLDGkTBQbkjD8LufTh7QA+uc0HEVa
AnfnTAPAG9/ByR8uhhBABU+bmEMFSvDWx2A/GUOJEQKO2Z6cNGLl7dIszzkgKcIyV2CyJjIfK8dE
iU7tBm2ZzK293yx0zYOvRmtW/dLhyyXuz23aEG4Wz0mNB5ffnuYysvzBUuQeXmC29ectc/e1nG1Y
flxrO2prWmZSQsA3+3tGV66EkFQsxQB1rvPzZT3Uqsz4RTAklZfg7naaZ5v9+MnL9+qBdkC5YmAK
o5/Mpal7YUXt3HXHjCUooK5lb211bLRA1s0FhCCmqXW1T9uq/eSzN3XsQjH1nvA8cLZOaKefHzLc
38bYysBZbHl5OJuyv8Hg+oll12qvgkiBOaYTq5erO8QVaXEBeCIVSjnKMof1dA6qwRIctHNCkver
NYr9GJBOWfr/aRWwXLPnuBDVjKsWji5khfSbvoXMKN63z4e1tJvXR28qvCvObe0j3JaWevcunGEW
rPbWqgB+1mwQNNKbdigWjUS55jHYrhsXaE4LeW6XC7xz37CWU4ZPiZ5KdIUgH/H2CtBtc5/PeBls
2+8oYyOEKE2TbNb+V/5HKgbAYulOKUgUerr2RRNjJ2hXREn4POMlLN+Auu/zTFqiyxrFcsXZPg5V
VuLn8PbO1kQrauf5ryqT2AGCmRz0YzUjIldydECVB4tKsx3yARUmuiwFGNDdaxfXR/+8Ww1VUQDV
rkkDam7YSH6zG1zzR/6GW/X7aPplu9iwf7MaBoJDMk7A82pqZHlttoDepBvdXiIwf0CtHDjY8V+3
r+6AZGe7c4Rg2tR4hhH4BLAAqyYI/CwoqnGX8mFOS3jHfBzlkq2GmP8yr8azxJNrx8nxfYf1I2dv
QXNJvLyL4IQbCjmi8kjn7b4O5/WTZjRvR+cW8DXpC2we/j5jKMnSorx5MEuyH6HJeAxRUZM0l2Cs
2wpx6iTqedNKKV4zOmxHzxp5XyOO+BP8ku+B+1MdlQ8LtyPtHQony0eVzu9gVAvYsWc87vjANztY
j7nkWgg2fMGLlubUhUJ8FHyZhIGPYk7U5FXRLcs36MFlmRJdwrULyfka+vxW8Q2KAPQ8dnlBss3q
LC/tS+l30ZIsI3/MLCXhGHJEOeQAzPwQQWFTARYcyDDS772EnpdtF0IGL2VgxW1hCHBBHFm5U/Ja
hLC4hDBSJiJzMhqOT5Ln0O1ZYUF7VB+R/QhGhExJhCtnOrpFcU/1SY+5MkfApQYv/T+0P7rJ63qZ
x2wXcCbZIHji6pssZsr8KlvideinJhC2hPnCR+1Uen7iKq8nB6OHDOD/LjLYeeAYThcZ1LXBTUIo
md68kSBFHpzK1jpFimmr6CSPcE/6jLbI1On0t3S/yjLNiuvOaYYRI7UtvzSAN1CyaP0++oObKoEa
63cPJFOMYY23s8rRZQCJTf1Miin+ZTHH1Hgxl/c6pH2b/E3uxKUmh0wL+D+epYa2xJfPw/9RJVni
HzQtAR59vKbwNQl/n9dwIgxdAaBKF09KZv5yazKq4RqPjIBkjgmDNPnr41WUJsSb28/b0v6rol57
znvCSGZl0Qm7QbV7jZjo084sYDQxkhmaw4qz0zU84NMkGio+C3eTE+A/ItgFK4V9Ia0xpwHZRd03
GEply3Q3h3tkGoKlOX8tw62kyupYiUWjfLRmZH6Cb3N+qCS5Yi72EXsKewS14mAdT/K+Sfoa3F2D
ev7BZ8PKyT/3IrvfmeX6hfb9FXCvRBkWuW5eqyNBqex4ryhq2gc5wXXywnUXLNHKb6ASplWpMiZI
z8mJy+hQ76NttW7lWK7zHSoYQB6IuC/dMbAAKTbZ67AaDFiwnixIdj1DyaIz0DjuCP4cZYaT557v
rZK60gprv64D+AyDQSzccwvg86TjHtwERdtNz+VOqJkBy5nwMv+wqYkTBge2L4ap7nclTMWlp+Vn
lKn/h2lkZ/w7KoyrZtPUExGaDS+Tq4JFEtIz0R2Uda7dPN9HhaskRW53+bki42MsGBZ1MvrZipcf
bzgQMYnOxFBMM0BKCOUHutMk7goAQ3qEJMHiIHTTZUBENNlGoTNVyzaVElK52vQ0I8DdAwJJXZYq
hdsDoCYP/6FL6AI8KN7tQdjBPoT8X7UJmX7KoWmJtBTSwwf3BK+lE0Kt2BXS7Dz5X0/msydKAii8
sz1DXXZ7MYCV/yFHRDeTf2WrNYRmdb2LKOuAY1ArT4aVdGCughC/oapnvx1YLPMKauwRJSWxou7J
ePhdb8DXgetmDWvHzPs3eK1bEKm55zylK2Pjj8SJ8v3faiIwPNtXEu3fmtFXW9l3Hxywrhmdypx6
r3vZTaL4iInIj+rm7YWmlUsfAvMZAE7IdqwRm35lT9DuGFN06NmM7jGR793IcqXzvJmyLdXWN+lv
MC+NpeqmKBHYKN/yllze0PlrD9fH2hVBLjoePrX4NBgkbu2e3QK73IjDSMgKpMsOlTbiFmg7C/kX
wmGkFpzfBH5TDuliYS0Dmf8uS9fiVAvOruzQaEggyOy7zC4jF35KD/y1DS3kRYqhWYdwI5Y3VyXe
n5m6bD1Sip+fssPFH9Z6+0F36qwUxlJq+SL6bitQgLBQTHXgvgwebAVxhuyWPX5U3V10gtabmh4T
+K+lg/dZ2NQV4w/OUJP3lWSLlsXmC7MaMaVTSqbnvTCCyZTqByqZdczy2eJnOCpovbCyDMq05GEk
sOPDQQ2qh2ouj5gmcKNwXa3QUKjPnIZ1LVjYF+3kTXNByO3E0w7ZtgvK7WANiSum5+8XdlAqKVHP
L/Oml+Ofp1F7gZA0r+8QOXlZm5MJT23G+wUYpmC5y1ETHlZ90mZn3IrtTr9jnrqPAN3zyAViUQyq
ZnfKfTXXieGB7HMmMKmzT71GtgC3M9bQKfKN/wAskPWHadZJ5pojyrEJo22REwBs6ttjiyZFb00L
LEhTNY7FXqQbiiVOmU1x7DhPJZ6y0Ygt26bjJeZJWUaJnz5jKE+sllNtHegEZr3THJpneSzllKOH
QaquiqK5Gqz5pvb8zz1GcbXgTkevzabKdPY7IIeynn0Da0/I5XJzPrEzG5iWhzpQxwIywV0AWQEh
agB7CjZGoCNGTrzEW7wrQCbMQEz79v/gVguQRDiHXSmJF1euXTdX0JJNDwaeOC4CLJl8l4Jl0tz4
oySkHk4tZ+wbsXrgYYvBx46Yq/Jlly6WSZ4YaXRNsITEl/cF8Fv6gNLbpLhpv0QtHNbYxDILcK3C
WcYlqcLLxwZhszdUowAVcjV6y3pKwbD2Bdk/sPceWbDSS+GaBZ7WHpO4rU2iuj3K8PC8H543CXh5
uVtuIk19MfvFko9GlUsiRdAMBuJ4zEEFewu9CRkr0vL5Iet4HWFZ4P59sZoB47kK6K6TLJ8nzU3u
NIx9BhNbTmu0rT/6d/LyPhdZRZypd+yF0Fa6MHTormI5+E8G2BP/49zK1/3KEnrJ67HFpVOnbaud
/mWpKwjj7Mo2oVpjYpWObThkf/7eft5l5GKBO10gAG1/otf6dHovvxxlwf3T+DM4PTfSgRFxForW
cuOOZ0+fN0R0QLCZt90p4DRINbraWBEYNJqBAB1kluWb2HePiKzE2f7CyajQS0N60h4I6MrJt6Vd
lq+T5No8rghA5YZdc3xZv1gMQrCT2tVzJjYiHkbOSpVEU1kdBdG20ALKPdVsEe7GgHqLltzLkkCi
JlvujOLTigz7jsjNpOoz6eNfpOZlFGOI8wGIYu2NO/oPrB7ZoZXE4/O5+GNLR1SiiNHNEBAUcddJ
J42ETBFojDIEZdD/cjtQlAIf2U2U/q/VKq8IcPuF8f2H7oDfXH41FBQM9mE0E7s65PSsdGubxrxa
KJWjWwRLOLr6UWSq0e46iETtoTO4PpJdqD/r45OzBqO4o1zejlJP7uMJG7fI+/PyBRheYtPx6LL1
IHptpJZU0nIEIDjiumAN2qJLGwpwDjpiBR69dnXHKlKbjegsLLIORoVeTmapICNQw4Vj+QXNzxZP
jfeaugXSWEmghv5Ii0EnrI1et0VTVX76E2xgISVigspqi/wO/ref0PpKFMSANFH3kAHWUmjFwms2
8vqO7wDAJMt3e1jUeFcGugOj8SHZ1mYoAPGIu0+r/fkQX4Mgp3Lgg540VqNmmGbO5Ez3VI2i+qp1
OjcQn9CL+5KCX2No+sqpDzPN00wa1EasJfNK/+MHrW4Q8j9z6c4KqA6AyKiUZEDCNowpj6xpo6mR
OpxAR4bOhdQcSa3XtpvBKiIarksmEp/hR8+75/6wkeF1hOn1zmhNrE6KHVK6r9Pg3kOqFMBbSYfY
4Pmz4IHaoQf9nIqZw7y+WeN7HKa3rhUVzt+51Zozd4kASTWKC/6WR7JIx91StSzJa8+Xy8JSioMz
O2qFUmIYltYnBxWoyeiuhgO1aAUcI5l8EBrouiwrjIjGJL/2Kjr5NuASEcKvzGlfxXl+fWAxFlCM
UvtMolunK5zJuBnJZTAD4MPiK/AL81GWM24NXKMj96puWS3Uo6/hNBTsJmqcI49r1sUXThqTrsHa
0FQb81NRl5uB/2laIyeWwfaI6IsVmiyj6VeV1GdjVoukepfS9oQR/KhnEvVpNvmElQNpnMUGINe4
B30a+v6+JmRBa/z5VbbYd9RGOcz4xJQm7tXiy2RdZYM26zCF8OMTGY3xC2CJ8p1s08QLhW8jnEaK
wUi/6vl8NBkGUHchnlS0011RDkJTC2a7MtLYnB6RAOHnpl4Br25CYSEKi8E7edRNt1q5NaazVten
7wAax9SMCV8+69Nx4vKqq3qXOrWRpFrnDbhFkgc75IeUYX+g121rSbYx1rsIsBVwQY6oeRuVqqWT
dhBmzaWDjw9kQyayZwp32XCslfxz8ZrKJW7oB4PZMZpSMpwa5kcpE2SxdVBGsL9rlcLDVPzQsznV
2uHQ2ZBV+GMR4u88B5RPlsmD0t/OsTB48wnc+FcImjUKbuW34Qsh9gabBlZ1B0YQA8cgqkcKQeqK
9vjBykJjvkHBXP+IXsQ9khFVlHOIcpC0/kgN5jIMloJhMgSVrwVydN3D79JqgIz5OMtZ9LnCL8r7
ZyRVlSTv3B9f7aD/UeDmqRUzorsS8jPy2SIjv+vlFp/gnmsKGkaLY838twRvwPdSKKBeVQdlyU1E
NCshG4xlwkyFaHYQRBd0LioJvbCi0/WsLdoDz829yWefshx27hDni4/yFA/uXiZa9qMUc8LGPdtZ
iCqPDqMUIzn1du/nPZJiZHKo1PilyTYeMTl0SGtAdnxIK5S4RMKu7ZY3Icdo/4h1T3hn+wpHNZhZ
rdS2+UtlVe6EqcqLZxPuHT7onMyPmTNBI4nwytfx9cGz5yrEiKcNpGYbNKavkB0NnXG/8tWpnp8P
hplS4v4rEcAjsZyt6xzG136oo7PGi65Ht3nmSNw5S4CN/JzzF+Zuwu7Y6XI3MAqZ21rVHtQzMCLd
R/f0PSIvLjQVCqRecp2c2mDm5XpUBh4FiTIZhR9sWF0QGxWi5+B0WBW36hByQQ4b3RRhxKTuwRG7
XfGgUMS5wIPoKz7EyVlRfhTAh/4fv76Dsvl0Zqghq0ZUNRnmEKBOAFuNwacC6+ZrtODVJa6bVBWT
cmdsxJpIOXgPk06dyecOUL4KC+rBFsSjgaNqFmhfnYO5/LLulICpxulJxnx8/fl/gA5liaKO0kkg
JDno+eVCa58Jrskei8ohvTEMmSkNfJE30a0bg0cJ24p/QJDEN7sAjYC5Wxvz450LlZg1kttwnYk2
9rtNQRKbFchSed1x+DRjSDGjtBoeukbat14ODNauVCqwepvQTw13ZF+ALF+4iRFrzCBNX0xm6oSY
WP0dM4jmt9KLw9hyVhnuHdTzGqQaa03/kN2TEUR5/Ek7oMK4OKdY/JIr4U/MdGjgkj/X5pZcmM6g
eb4HC/bLiiIV8/W3Luzb1ZApiU4rz2naCEGBNiJRFHbvXXFlHMeWxSfIQv/VTAvlRLqjzUISbKJz
bqqgtGxuL7pJP9mSpGENpWlWf7Vz0TxhP0n7YjdvZZm1jTDgIY62jahlqP6KA1Uad2UYbEQxzK5g
wtBnXzt1ssrJbsYbacSYdVr1fCwJJtbcVDVKm3pPd6+2EWs6EGV/fSmntLIGi220vjfd7XREbpiY
DK3Hcrxp4Nk4x9MbrOTZBYl/VS0VcYJEcsZFzPjFKDsoEPeWBevVKMR1TaHoTV9oVUGxEVuGGq7u
a7vqc0cG/wjUj49kzwCi53X5N4NML0ab/iGQek9T3xmNeJLHGczYvKix/9L0AOJOPLII7K3J8OZP
yuy+oXD1MeVx6Wyizf1v17BQ/AgkKLn9qOvXcYZfDSn+Cr9GaSL0hzvhSvA+XkkjnCnFzWI88Eih
8RG1rFtRVrBxc28dl0VAwH4sZ1F3OKHsSt+7+hHmJvcIon1TGyn+Gq3W4bgllfW4E+tRZVpBY0nE
cNVlQH5vF5E8EZVJg1VSr8uLKLYY4eWnm6E6puVSz3jrUIL0iOnSqQXt0z91hzINqRFZc/mvO7mz
ZhIYC2IQAAT87ihJ7Z5CT+117yQg/BM34brxrlZF5u79kIMENt4GyTYfDn0aOdoYkdC8o4byvNuP
rHy+Vx+iMkQNKsBrVXhC0/EaSO1/3JyBBQ8peRGFwfae2/qEil4Wv0iqM9/9sQs+1xo9dvY/zxRO
hBfe6gp3l8NlUUkO4mvaqXNtQMsd7ngM8z8L1WtxKrWqH75ahg7v1J85xkK+HZwv/MX4jeHkRKLZ
rsf8j8aYpYeay0n1SUReUrSM8ekX4KaAOtQirI5H8AFVOn1JvsfAjLHAU9Ystnqa/74haofnGFW1
OC/D6hAmvUS+BbPtjzxPno3X+vXapcb8HFW7uSPFt4iZ3rtFj+bCqyb0md7D63IpJUMywbCQJx1Y
ZQKB3WHqK7pjAB/RKo+YccEXy1vJ0zaMLUu11f33JsMjSawoIlzcOP9+zris87DHGowY2pxGgMj4
GsG0XpqYzzrhx1UBVB3bUPyQ17tYPbUoIgLEQ4uKtdQkhlcGYwdVVVr43wZ21Cbn+eSnbJvdrtLB
ZzGNA5AwhVb628Ou3Jf263ejuSBD9PCAGn4C2eOSXzk/ajMaftupmpf1Y78YS/Cb3HGPSd1Y3D2k
NzobO1jV84fEl2x2NkELXQrdv3T5zKx1JtsJAXd08Kuhx1U0q7rbAweoaW3f/aMkOYGuMg9crA0v
Ih3WStAQB8Oqs2pvHB0McnbtU0Accm7HZo5n2SjZhEgnOVzlOpfMSHq6pup6f3nWkpB5DYSBLuEi
eC26afwNgxJrmC8zYyGFb4EHOSDw7XOWKfBxh+bAKGhLBFMiOOOWKhpmWbyFUlxiUdPWwC3HGZKX
qkaJ1DfrrLOIDbWZeeUCIXETpsmGx7P0Pq9u/OzIyKiUzFiFPc0/Jt7s7JFsHv/83JbDwzxrPFHN
cwVWsvXzp7TNHp0+YVLbvzf2cHB+yt03S8D6r21BzafKSyDlbJQBx4rid8oqYD42qvEMnG3oUzN8
7g3JdhRbJu4bRoLrQNXYCi9+w8fGezbn1dS3D4pRgp0XwKfkIaWO2dU8pp1ZnlXQe6cjj34dMQrQ
TsvFZvbMRZCFliNNx9fzyfBR7qLqSolfjbOaa5cydfOFThq7xtOCTRK86zeDTCbaJKCKMO6ctX9y
NSTsnDJanrNJRPahTCAT4QksurMXfbSxrQyJKTstKfD7JDZlPdO0Xz2ywkI37yhQSH/V0aHIx+KH
NgBuE6fw3uyPSSiK5tZe+W/06afWIDrjM2ZgkJBfe/gEmRDBWvqgBRBoinNsj3MpCxDlpoc3k6AK
2+weJOX16WcFLdYZ0VkfVc4hVey1A/WDL2Cc4bH/qm2G05yfGc14CC59GBNy3lHYa3KCBjRreKfD
1X/wf+RpdEH8Ov/PpYSXzt4+YAxjBcmGSVVp8Z6pz57GlwrStXC0pwtfqWEP3ujF5kpGTImTFZIS
q24ptrnrgh77r0E+9X23lrbrEQm4/bdpv5PQPo5sx7c20A6wDkZROtpm3PDUNB67+WcC7lnGckYK
J7O8tNGTcEcU+HIjPZ2zEWdBKuNl1m5tYB3X7rbhxqPrcjlV5F+5csTksoDimlf5HzqqB83ughru
1qvMOWorrZxno4kd51WVb/nMKuxU1c2pOm6JMrfEwbnEL/6UR4jvlpSbUzFT1piC+28tp2SRpSws
l+ZwJOizIkXOuJBdM8NJq9dNBRwWFkWPoPrbAt1ondUFdmyf4fwjqxYqui/PzScYmLLCyEUM5XIa
mStaCvWIq19fGpOASBjZbSWzT6JZhTjvQ25Azyvbcv1jHPvWJ9Ca3aw9TrbNLwdbOo+qltYhZuvx
oPLWtWmd4YGxoK+M63pVd6YEG4UwoTHeaO9QNJ/qNjliNpeco17ogOWdK3EafPek1HhZKvl8x4+l
lsfongunVGqz23Ls0PCIWJ3ZCPlcudZOg/CD5LLrueRhGmqBW+gJLVIuOpIQWvDuQ5zYnwtff3+q
3wgRPk2rCbVJaHMjbieTiUktVMz/Hj5ovcOTXrIjouJaNsdwTcUHRrb6NMJAdn8IorTaYVZjUwJ2
5RlhddsVjD9drfLA6UkZ6GxE3psI6eZ5Qme3ghkSRNAa27fG5Lcu05ugCJEjxXVio6tIw1P4F4D0
Ib+RTW99XKuFYj7DjRAYmk83ReHfgb4DasR3sFpz+0/jz78FeagsbLPoPWCpObs9kvKhce5ePvMp
u9Z3N8XAom+btMjuRyUgMG04pkHv6PVNPYLwyDXrW85KI06/7tAdV3G5OZ/gujTApqXSZqIknY7x
kOIY/tgETMILt0affArLE2LwYHWV/p91eLyGatdu/1bkgqxSAaknH7Y5u9qlByc1njDKYSv3B2Jz
sQlQKdLhtAEnu37/18VUIssxrObVcJWGdOGtUa4mLCzErMcZWUKF7rxreoO9ReePRZUbPZMQhN63
3mJz9Kig43HddJLMdvS7pDgFwYqcBkldpD6+HvvpISO+6uML2wKgntgWU9o1gmOQHrKM7UyjGCZj
lvavPFPrKvfqlTGW+gXA/er4u1LU5YfkB0abRaU6i4TDSGtWOfLIPFHoCz2pbA34ZY2I809PmFUz
uvZT0doe12en93NEi1/SBfHLUVxjdpPDPK+uIR1+Ytb8ovqG8OdH5HZKKLUl7ooMKtXOAqSQeNyL
mxLtZq86bpoquBgvQVGj7SEz6w/VCP28ztfbCJxSuSlElWRMHNxXBgsZbtxjU2+mR+fjXUKps7CJ
8/4zT5ZuRYr+tRMeJ61UjuH79fD16/I8pj0O2Wt9QEcCCcUxfZlplnhlZr/Eg65hBT+LJv1pabRd
Dy7qsRrBkQEhiXMW0PPvoIBYFhblPoSOZ/cQiRLsAbY0Ob1m70y69yd723NxB5O0z5NLR9vGOnwy
i3WL+GDLG0CK7dKnrlpZnBpQasLY4UvZBehHjEb2GmtmnBGZSLU5HBG5oEHiFMoVh/9rBLzK3w9v
x0a0hrH23uRFC0T5F3cDlQEAGvMu4T0RnmLtkflT/9jhtYZvSoW/JMOjxJybRSdApXcONNPgzri7
+QnY7iQMjMMWUVXJrB59N52btA+97nAxCg11fgnuD0sO0oQh6qlrYjPNg7mDQZbyU2t5gK4K1Rnm
80omHXR/ZlNngvDAmal3WFQ9EMA5LpXAx/uokz0XIeicG8X736SgybUrsKrC7Yl4/yqBQiX19o3h
gOve7TQevRDQlW79OW6htIAeqqvwMkMBJA7xSE+tj/q55cSWuh6Oz09VfZm2+OwHHVxMMCRI4xMG
Z4aBcp35ZU9gRFfbLE37jegqlNcgdVFuqDAg7wLR6QxeU80NuOZ/Ka4M1YoQhyHTAwpmR6eoVALh
w7HvqE1z4tDFVt3oINAc6d4op5/oUrL0zo5ndBe2o6cGqvLTxPl6wCV/FZqfum1Cba9s0FqZyHFz
srwpbV7wymOr2DT04CcQLfySX5///tfxD6ty5fpFdfE9536vuzi5HgT7wDYLbE8SQ6U6TfNaai1P
qR3KayZtpILx26wmZGtOLhnk8uNkkA60IK9z817oYOEou0z/OyBk9M9h+MFHi5EJ7lk1d8viUn52
Kse2UEYptV8pZ3ec6Izmg9mZFACp09H9+XyltPRTuwgWGZZCxjxgWydgklCBVrRAOjPVQgxjSrNH
F9SQySGfRbFFxaREnKOXAQ365KUTg8T+1ApoUwHr8YO3T9yMK8ImItD0nGLgEKB3MtOeVWZ5/23b
1QS4/jdOWRMovnkyI91g559vC7zJOculYiKcXuU00XagiPG1EYiKbRJ/WiXZ91JbWFOIzDcc9zjI
YR1XwFSiw+/bqBb1J38mqFxB7MY8OK/J//K9h0ZLbtJEUq4RSTeNBp9OsiD6XIObfNenIpFDBY5B
MNG+egjZyKdYMv1e/dkKnWU6kE8PeCLjFFk8u3ZgRkGlkmfJeY4S0XueZpUaEcdDjTSO3ubL5f5W
bWTqJ3ZWK+B1QalRxzedlmrUr/tMkPG0I3Su2qlB03xWTWiz7DKyjITcz+hwBtB9qzEbzhmhXLjR
6I75cZwWF/dH3f86NQEN2Y6ll22XznWKYdi3cV5CffkullWhAlWx2chEHkT8uKx3oEt0yPUhpRWq
mD/nIWcnoMSM8K3tEKLyVNipYgFT1PW7mPgcIsSrZAwF4zgej1kxBlycgvYtJ/dxC2w1MBnPXrvi
qUGDIwlQrM7hLjSdvQDCqGfEWV0+DCB4CX1kTXHdVllcLsyNRXtKECJLhdOJO+b7bppWGOi98+Ah
IZvKU+nLuswIAfiMCqvujhrTNACdzlW7WflqqYQ+Xk2Alw6Kay4hGX9NbF4nrZ84af5wcrbDMl/R
IN/LUaXt2j27imPd1+z8zn+oFGJbVGh+aU5cbiIf1X6OafqhFd/WT/kFgNfgXujkxSEbm4RRB+tr
P2pTY5leC/IuIkO1ZTFOWj0yPzz/N5BlYT9r5VNRCsk+g0GpYR+7oh8OyIFr4N/OWFDeQypkPvIJ
ZT9q9oDd5o2YaHafXWFJPnMFj9f921F61UBOkFH6cU4F0pjZPH3/hMN8QEe36KsynwT3GwhPGgdO
lMyd3cgzAyW+TXMLig4+5JaC3B20nOXD85QPqcN6CGzNrq6R7wbn+6mwd2tOhWwkUHk6aE527bXC
EM3m2+z1lYPmgQts9yF5rEZxz2bgdYEISZvhYPpDftmhNSKnpcE5LZS4sIwJDPUOYNOGEP5AWOhI
1zGVTvID2Qc34sU+VZuvIKAStALX/uBUm6PGHcQ2zR0PaXPVssZS9BbA6JKzulLENOBN0XksDYmR
hnETw/qDvDtvRjLdJqRDISqWwl/8mQLjgKpXLwK5gJwqM0NgQAvbjAGVJFoW6YQPn8WTljUqyiRa
V0V2uTgjuL2xIvrV2rmuqjyuvohVIJs0l8VfNofTgA2mh517WzwN1XimGx2gGNYRxm5WA6DsoYy1
pWqHYm2lTYwfqJCIJJEACOPl8l4XJWzrSVn4HGV6EMN6/R5Ur2zamFtzmfPVMIKG6NqxvlWU9ifd
/IjyWctgEF2ae8yx1VStkPRkhOT3FWY0dBENvjJFLSuwPaAPrYZN61i5Zf/A04T3eZ243LsI07ZK
+qqX2lpw6PuplQS46spyZ/30iZmRipLw5WIie7VAh6uNaXYTvEF0rQlPMspFMteGr/r2RFcPKL7T
ERoJeUr/ZBoMwKGddWha6yVQz+6inwC6n2v6CU+w3l2Ni5rAKQhFthzHGv6VvtcpAyEx5CMwWWYQ
94sqWH1Mkaxmt3pwIyBJ7+AtfT3+qVb5cF2EYLj9QyBRhw1o4tyzlOysLEqOr47xUWGicEJrrMdH
eP7LbExisRj6o8NDnLheaGNSg4W+nM8QhbfbzA4UN+AwD4Of2r0lrNNHV2OH1f5yUR0hgIdOeG4y
mfnZmRRbYS9z8pBEW43a15rRqSihVg2nbWvEyGGlQZRzJr3QVym0wCG7f7i07vjMqJ1mKrQj2ZMv
8WMQqzW4HUJuLTPcAxmDmvFmpysobNdCEZvgCXjvJio0nzjjfiLhkSgUgXsy0lh/Mv136DN/zapr
SKHiqPSxcKwKfiem0L3Pg8Df8a+w2VgfCvWrfXU/r+JdvvQxc18Wi6q5BZwdwNkj2YcnKER02lF3
jnqSF+gHWZefyv2ZoULC05fP8sgSWOKFhYhuKZ1fOOk7tElXPyiz/mBvm+xOFxFnj1tvIvzwOwZt
my1JuPhmmxqLAAo/+IlhVbAzI6fPf5M2iMffIOT1hvroifwkvZUVV8WrSUFr5ot1UjZkp/wO5PLY
6eD6jlGHgCXIXMfMZlUOYOWtivU9jJLGxnZlX3eqCBZu4JvIHMF27vU2AbfIvcHXRqRadYczjgdw
6T+VZQjHQjKq685911cl7aTw6A37LjF55G+FgwFe/AggTcDj9HDQ5u8dliBQc4R2zCAZXZlLnu4E
FkK5GUQZunJT/wOLe2VdwBsuKMVslllaVdPGIh77Nf45LRchHSY4OzGiBW6/1h9dWfhRl2HPa5+z
unECQBN2waUPOltS4iXUlzl0utbGlwFMYS6KRKd1gyoIwBUEw89N8LJeqmbPfGnzNBSLzL4LADmY
D9cyYrKkWITBc8aCSW3ypqt9IqkBBJSAd54GjNtLLaug94uc4sY+zSJiOsufEelo9euWUQO9wnm5
cdpUEg04ufybygYVmpPS5f/bcpcTPZvUE4USf3oOXTDBeStVlKCy+67DMjUlNHdA4Dix9w5RmFYr
L4wpqNYsBskiWIl40oUpZ4UvzDo6JlxWcYUfzZjRlnhZCBvYWevwcImpMdlSOGbZYuJV2SQMSzXq
bQNLoS4L5UFI6LoMy2KfrQwG/CH1R4HO1mxgfxBizsEx11uJCH24ytV7t55bbuEIQpfgynmmLqpu
pZV9TUZaFaeUZG9CaWPZUsfveYEU6DeYxnXgULrBcKcl96wxsivIxjnenr8m4+60xygOE5LOFXJz
o/ki+M0R2YDihVXFI4+1WOE17tkWGIHRok+GYF5/t2iEgWfA/4ADvl7KrkFctAItQQtdGGyvE+fN
5sxBUbzolJFUSzISSQ9sqbjQO3QCwfdCqvhazJivX9fPegAcbwi9ZROtpzF6nQd+FwMXXm6hbI+f
XMJHeJGbR820rbV4r/POgbYGE0+NDBJpip/nb1hUWNYZSVOUHyTf7GTu7dKCpqAPVsH7IANwG+OD
+23+aV3itUBDp5Vwaon38MNWMY5r9ma9pwEeQIvLWObkBDD+9Cy1H/R6UKwN32OLwz6xcEkYeUh/
YjfZqJK8jmS9JHAaPTPfJ5ltwflCMKmzzNq73Z7q3aPN//cAo0JALrSXp0Qa64P7xRZk5l6qwSfN
WWZkDI5ooPFs1KNooopbTPMXMIuZYWy9Fak71NnhDux3XWiTXYQ/FWLJw5n/fdWbxQbVVQ0/rHjJ
6I0byr7wi4rF0XWy1qFy+0Qr9zj9i6yMIVZZ/3VEDBy3eozIFUHlsXkSpJiT1X1oXTXqvqOak577
N36XWkZgFu6d+Fqun/e9YH+crLvLyYxlpfR8se1ypWas1TMyG4fM6lwUb89fWS4FHzKQZuzUelZS
kDQbbls38Ck9bZZLNoV9iu3DVr5cWcbwjTBUzAOuodCtft1DEvbLEEJNsrPz/fXgChYvdNsLzpSZ
mcrMCy9EmNxLKS70OveVE4t/lTONIbkcSTkCyWw8mhIBYss1o7lOHtjVY0xvWoyB/KhFXs/3aINR
4Sb+pmrMLpZ5q7EXruJuiAjGoikuNNK9ui9D62DZXnPinwe3Gt2Dwu0Ke+/CyLv3EAXSOuPw6cvF
SefbD6lp8tSGz/VOuRFXjSpEvH6mBr7C3RPCrNQNspsM58G/8e+Ek5Pjd2w2Endxf2CVcPu2ICF/
mfjdcH6iZJzyiTt+FElndKXAihy4pk+etMyKLOFLuSEs1ZjrIBnd8DWckLxTvk+zmnaYIsAmXbef
3+SKbUErv0UWgbFDLa7VYRtyyEn2umg+G+GYuldRnwOhBCXWiScfazRb1SRtfdaKK8+D60sLQnDt
Qg2Qeoz2uAt5U1KI9RY7QU6hlRcN77ivJzePiZk4IHbZfawXO6a09eGfvXfqNUgohfQuvkWpoz+v
QXeGIL35QBtUSNKl99AsU0PLdG9yVCwNecVON5ZADS+wvCvcPGegcXbWbHRJIKVff764lmArqWaS
wglIIDVGSKsmo1BrIvjJPalix6+XYb3Ib46QVYAojvaMxPsdDbjNVaDk9n4UR0jrsmhljCHS7JQ0
iqzJ5lPiz6vea3uCxA3y8U85wFclK7LdHcuhdeeLUG4tNmRJPImYr+wFjZ5VlM8q4oMp8uuQ8ene
+27zPLibMFmNh7w6+ylXGT0P7KtPktCTQZ8wDI7qDJrL2pJ/BPV5V2BE6titgAKuEdjjtD0iBKVO
QfOHJrtbiE14HssdrfJXfv45mI2Gn67kRg0q4jBW+4eSozRFljfH+QH4zmwdmbcz+lFZapNZt7Fb
IcMNAGr5y7KWGuoNjZjvOAtGL2GDNaS/+Un1BlcIfjEGgbzI/XFQrZlDshcXCkUjaNn2i66NYA1E
8k6p5PObpI+ZulXihgwin5BsFnbrsbpH0ygtG9ZVC3S8pjQlrWpTLY/Z0P/Mvo7eYIoskQ4M66or
S8/ZiXGBnd5GQUNXhAwfJ9T/ripgAFA+jGHtJ6efhvKTWt2htbvaJCEC4wamrFdkZ2/pu/HsVR0u
5IJImnOhetABaoS2YU62RiJ2T5yhUMGvp0cUSso2n+/UfZddIHB270QSlDH/ddHCy4fFurM/zlHT
MAHeviWdAPK0pQ9BGzumuUq8yKAtR+Sv62TUB7Oet7f2pjO4xKvm5TFsDctVk3D5mFJKfBV8dLdy
a5u4WwUJZoOlmvfb5BdhYs+05j4B7RyQVYwwA6sqFh6rLr5EakAmXSvUWmZzwfCORCX5nLEoGS2z
1J+Q1o5YbLquxxK52yo8G0iIRARd60sqZIcuGZ3O0rkPtTZhY00cjgxWT1QQ0l1D5EqZmS3tGdBz
5hXF969+rnc0E6rnnrLYtvzWZKkHcYQnOD76nb0VHydzfnnQBt90Cvc5uUpf/HRxHgFJn5638b7a
N75Vdwob65ogUv+4Pw7GZTwOsvym3H2JU7midjH9lbyWNSWTgxSDouPXovklQLeTCuAqk2aqXKal
NuB5j3k8tLYNUvhTqNxM/jtskqLDd7z8TEs+HAOIADvw74rnQ6LUNf2mbTljXXeTGmxug/QNTudS
0D+PJDb3HXDtO54tYKnabYgbKlNE5h9RhiitT+Gx+lnkH0KxfA1ow2piTJgHNlzO17q0qwWinCTD
ymCYEBew51DJZWOZ8x3DOIkpw3CxBXwNeN2T55E++KwFzpECi0lCU15iUjCVutkkplOPPjO7+4f3
WW+7yF/OEXRz6cET6MkJKumC6eDV/jQ1XxA+Ony/DbPM9kesSd6Qy870Xgae3tQv64zGJeWcIi6o
zSvpbvBDVXD3IgErELen8ZeRLxYsypmk34Eu5zeZ9uMTLFBm3lIvqHabSkxysiWzRJ3t55QZNqO3
vDsHb4WaPqcW3YkbfVjds5q5RwvjkspT7c6XJOdZIVnvlDwTtW/yfhmqnGKUf2xPRYw5smYgJAma
0OVb/QYApbH80WUYNp4cMUtfcNwhbfXe9xB5bOtgG60FDMqSiIxsgoHUY9jRiwz9wto+3n5Al4oe
tXp+bc0qPaNF7TVbhe/pzMCn2N2Ak+ACr7mWwTXjMtbK778Dl5egOynA5NFMJuEcHI90GdCDF5z4
etBEYXStoBhk34XZggnEHdarT0EP6eBxPJE+8nggn2fnjYlDe7n68EGCQiXo50D9q9FDOKp5RLgc
tZ0VtxauDm6mmzEHGTXfyDKuDTUOTPWGCaltLMmaFqT5nO8POxYdmIlNwcbfXk0wt5ns1BTt62VB
hF1c2vTfZaiNX6F+mlp+IvoEOiRqD2rcgwGfn+zOmvVVVo1a0tiS/lREMpHjbuJuxytZCs+zu5AK
AiiWRCjE0ysLBbMcnO2KyTEyRnO/iATfqMVa18ZMJNGoHahLjlz9r++4oQ3bAlK9fDJr8tT8L4JV
h2MwAABeJ3vVmZLdaJC6Ach9wZ52bjrJErVfVmlxyp1MIkYGmlRpetKYYHztF72gtUfJ0T/AkWQM
k8FDdSWhbQhIoA3KJte4mD+PLc0/Zr6uEAVmCIGtcff184sosLgItCUOYkx3nsehGkmgsWPBr56u
EU3lzckNxMmi6CXv0Fbo3dty4lDh+QkyXJau8qCrc0SGoBP3NdxHKeH+Rd7Yl3wFQ5BBTKzEuFZT
WxL8VmWHZWZSTxOZz5ZOnntUleitJ8f2B7yXNfpM4Ln6IF2PLiOR89qeBxW9SFQzRM+Q4GAPpS+Z
Gjq8ALL50oadZ/bJlOJ1XdSZCh5hPE4cXXJv08/7bAq6wkwzBoSQP7rrpf79FV/zsoXhMO/fxVFz
8GmlKhQs/LKSahSPVE3htM0ixXanxKHZJkGCfs06QuJ+RWBFw5jHQK0UmWrgQdS1ln2jB5SwlQax
u1czhUYMvbsuqWFwYECV77IahjLrvX/alxfcz4PkoyEg7AxWQacyXrsANCKdMMXcBZsAQJmbDpsj
AJBhKCt1ciK8FwIlhmFRo93l7tlr7eiDXuGqsQwOlkg+aOBVOjMBXuZ1EEKT83jETG23iQzNM6SE
IsSJNTPW5SzDIuACJYnXdH3fcBVXUtGgzOykWjgi/BF51A/HTuyaSyydIqZ2prZ0bGoVOEtsDzpR
H15Vq2NuGnMd/vvT2PACha6EmeGKJLGvlTQRyHOEANBh1C2mGsuT13CopZ8EnAEyfZ7jSZmhpHRH
oIkcccLRTSYy1zNFVbppTWXQ2ijjRxFnhQ1eQu7xeMiElxoR36buXie8U6LkX3nEWde+plKz6diA
1bfyTjSJBS2zru25DG58NFcxEG40N3jpWxujk0cq3pm4IjqZ75ORjQL0hGrYhLUfCGcMC9O2rj7i
eb3F8gmhTpPHwUevd/WblbBxDnMQbT39ivpI4jPi5Us3QjZpK6s4XC6YvLKd1KG7AYXCHm/9OStt
5UUClKJrzebwixVaGS/slrJ52FTP2g5ZnY3VsaUm0l4YiWDGd0/65fFAmZapJ2Z1xWytpc2nI/02
cE7UDQdsooytcOmLpkwGRGbEPgI6iCeaKLezBzXIwD+1ryPntaxAUYO6rIaLPv2Ew6gPJfYcxN7J
xSLsnRVJoPjTMQ8j1o+pQdKPyuNl2cIoyWg7kxr4oim5kxvjWahJalScWRPiZPKfhpIHKgs70c2+
mDh4D6/ccEXOj42HbcsIaHQnDGD6tBAo6S7DOSu9WRevd60pbma4YNtuKYUFzHe/eE5UMRJC/xV1
l+Wk9oUDwZ+E5fDMT4GaPOfSOHYAegNQPUNJZ2tE6YTfddkoSH+Olv+xgAtKXpfCKRgmgwsN3pNo
ggOK+r0nzBAXUg5wn5nIcdWPnSV9oDsjeNMXYbs6LdxhwD5VTjDomHNn5T+gVTIcPttzQlT2Xu3T
okqv/U3JRxzhcy9Ih/P1rdLPqXw6VHMeyK1LrvmS14RlLBE+HmmfuYdLUT2OfpWTR63Vf5JuI4Yz
q2puxV7dUMA+/GRGGxrbxG8/2Sjf3xjbf3h20GEgD8CsNSBnUEMRxiRjQlocSyKJscLZKO0vXk7r
za5fQ+VcE9VAKeI03GNQr58+tqC+rHjg3DySfW+21WWFmdy74iEIb0M+DHWHYq8u0UUWMaUh5dmV
TXg52jR1WK7bb5HNJlyE0byFYP8V1WldRyFTdMROxbgQTc64q/1G/OscWhluZ78SIT9YRnI+nCOH
0lBHrfd3XXw55IjutzB34v88jzUxoHHIK+RQi7uLd/pktWG8mSw8Xkub8ROJoxJrAhXu085O2ded
WhdVaCiit9y1iT/RerpN/3oyMnE6q0lcbK4zXw/1me1JVBhxVLhSd7TzH6Sp/0NBH0PwuNTS9mNM
oxOxKXisVghAqW3j5BwBbqVSuq1a81Ykc8z2PAyJyStEyu32DVDSU2ZEidc5lY07Z+sz+z33EPtO
mAtbdsaTC/27j2qU9HArrnpIKLTxMjHNDLqyNhz5V14Moz5mAoLsZRM2vb5C6pYuY0fvFkCFRR6g
OCqlhtOIF7jXhr5a+JEN1n2eAPv82K/JU1s9ykATcBMiAyWq1npnebUH7xhyZzv3VFZnqRJ/7Z/+
RfR/7NhBnlRmfrsn8l4CXfQbmKMqeSUoKS1R4LUdb3cbP3SkCAwnqg/a8Y32vU6tTSUTWdHMkDZF
LGQH0NYoqMX2LfPTXfgWd1YPKe+ddkwqgr6XF0/yd6Gtkypc7jI7/6Acx9rPA/Zc6D3JPpSe88Vx
YFu+aWxJpb5gu6cM8YbeJfVva5NXXso2DZ9G4xHhvb279ZZgxTP/7YES3Tkj42fone+rWMEeSDVs
vZ8w4/lXr5O2wiMZfLk1Hfb8tmZXNvPM94Ug1JT6jwCdnrP8LsMscN0qkyakniYLEyre7iGecDZD
X4W/VtbVzkbsfLicLBKp420LOyu66z4YRv54udnPSEwBwauHpWAQZLlJvyTBUKQP7OxZNMiAbOro
l4U1yhshGSwHrDtVjYdCI3txDHSSimRhFqDbL8zZTjq602hzvW4+IR2yLjuGHdAkEkRTfAIk98M9
V/duuHk2T6h3JqBz+OylOubRBQlu7/lecF802Jy6SLn+ftDa0Bxl9f1Oz5qSKfTtZcQXTQ5Ojv5P
U3RcSBBIrVVDnLHNya5S0+3sEVrJlWR+2jk4JMTAIOaJEFUYqEL3c6ivMuakUIi92Ri32aSbdop3
7PfVPokwNQkX71gejGWFNzsYVngYGrrsnGlh96aJmCWrcTKiQzJEcUdZTajxAFqnsTacyO8tL78l
X1eVZSZdCoDq9Wqoa+uCnutn+pzTANhjtImUeHljb0kupiiakdIwZ92uxiqIttaaNzmbkHJSdFKK
CZ6TkooZTSy4bv95xBb9FL6I/AfqUWXLXarqhDXgdxwrv6m0ZoA8Q4qlwNqnhGzT1+kQT5+qmtFQ
1Fto6pug1jgCUvBC2x/eo6efmp1po4xZAEZdmemUU3nAXFiaIro389CxPZeInkMp/w5dqQ1OsRPE
YSx7Uhs8MYpVso7EetqhavdPkR6/KuG9O5TnygrF+mu26D2gMU13ZgEy8rzKjnsGqP5Khv411aMA
CugOs9c3H27vQT8k/+gWZOulyseeKSxwJb7C+cwqh70mCkKxVgDTENVZhJc0JF6M58wlKBA4bmug
mD0emyhNmLLVKQWj814um/jOm/e66CUBaSa0wF8hckBEblENlFEjrF4JaOmHScU9eB40EDbQMql1
LXyg/bFjc6D1q3tTumEEwzTGbVHqryCAoGaWhybl1cXLpGS5nUTA4Bznn5oqWSCjeIrS2J0cjFFP
FGcH6FDHcTxwxFYGCVE4Dgb9Bc5TOqcWGkcWPIR4SLE+TLXYrGRbFn5ZuqeVh4udAJW9Icdg179y
BetjLE0MtAQyWdAMbNVAOLOlKpqSjfsLOn/aFNqdIpWa793vimn97DJnhlUhhvi9aKC0YmEE+cfM
VDse/IRtCnKqJkdXaOQvxR2LM6ZYxK5zr1DkTQEy8fHf6df9xMZL49wTH/EPk8Rwt4WSvM8qqWLq
dXZYBZDfvMSjFTzgxFiWcOjU/JyvREHjVh8NKhGb7EBpm4LQADr8hcZ4PyXKDUmCgulu6H1B7v3l
rWXRXiVh/YzxnDOiXfXNiYS9TNGi3h6ylDKXs3jHS00aAMhan1epxFeetJ6sBX7J2+nFXBvj6P8b
Ne3PZe7q6ArH/DmzJEEUdDuGVsgm4I/9b0n1TyWDZ8A5/toX4eA6syCoaWfl3TR2lVAFh6hJUNSn
EtXjMSoCtP8Awfklk0yH3nMggXXPtG0RVbh6MCdLhXiVgQ1IacyLo6/NCioJGa5W67L77DE7nSnH
XXLKp2dlwCVig4Ptv8qhQ+vwCAI93ANOI8wrhhl1JA3Py/v1YR7miu4qbkBj0kLiVHd3rplKf3Sn
80OFDtFHCSam2JQmgH598Grkf73OzFwpTWqVWOsdtGss+ZvDEozKu47C1HONIViNT8Lm5qqtC+bW
K7qB89VldgWISRq3BLBgbjtXahZg0BZuIXUoltVMnWHot+PoNR6eX0KrrHGee4xIvUiTXVxlNgSF
P9NifXdlBy9QsPC+SL7KqcsQDYlFzN8nWWZ8URfvaAWGjCJjosOlc8Y8K0iQvUk02aiJCId3K491
jYVtPG9eDzmw9jjrxGIEageS6SmUWMpXAD4OtfM9xJg+AMwB/cK9FNDk2kuLASr/PUVWY0QPRuu1
8kK7IlnfxiekWc5iUnQfoO02Pk+OoC9cmRhiGTClYTtmVG/vheVnUdf/g7LPjdbWOWmqSPdDPo8x
8ja54KhXa6HcOAYZGnRvlBPtB52ofYIAtjJcv58xBGBh9DGZtLTXC4gdtwqtoN66tkox2+Ha9yN0
sBSskyEFeVG4uOgj7ZHMylEUBLyYkNN33YbvFWyhCYBQARRnO0kBXMW2W+tnlU92eAyEuIqtbYCX
kJI/Dzz96bmw99m+HtG8vGGK7Pm2mpmV+HlGIxjghZI/ohOx7STvCZLvC5pBtFDtAasJvBJty0uY
ZCQBOm3d1A+/lUp0PJt+Tc6/DybneUwGAn7ybCbaa17Y+KOguvT8Lip5g2IePAXcAKVQKBcjLwi+
dYaFChcYYcXk0qJAVSyROWvA+eMKVST9V/2n23+TZmUhmMoc7wvUg4FurfMRgzTZ50slRbQH2kD1
wFpLMVqwlCRQJeXWuQfkh9weDgcN3uPL/3f+Kufv06ohCt9q5dNZiNlD3kZgDabcCcdwRBuBxyrL
9kdMabn6Us9g+yPXg29nMHpaH9rY5mvzzAq1IA+OLjYcJk7Y9J94Gm/Qv2YdHiAZVXnFCaQjlJhp
J5NKiIvA2ATo1rppfZmiaYFVyniyI1lMLKU4OKwlI2e/DlHznDydfSYZgrpTZqk/GN/l2LhSo2RH
tWraY6ibtTP85MDWvQUEu79LcrpDblRlPYskigF6xinpKzQ5uQoDAztlODRddUTnEpBLQWXGNsvL
tXyoQACp8BoWRGS653fb6UZh91q+AQDUntqg8PVKtgxFg2N0DVLYxbiSZvl0yQzxMNFUKgMousCB
+LEQb4Z7DHFkKSD+PXU9mpYWHp5NNbqG0Ulx6UVnWPlCEdwH5ubuVEpu0hkCbZRVeA1VV6LFr+V8
d5DhEivvSiJXOueQu1UIzel6CSnwKXXKu5TxvzU8eO6+xCkbsa+8NoBkFAFtir/7xDqdo+49v08K
+CboDrq+lvVmfSRgPoava3fULi3FglsJEPPHR9rN1CbpNF3s/mOAI64n3Nk48JdqN19bUx5R/XJQ
Ddj7SgnUqdVFu7W0QtbsphJkofhtBPnxFTzmRIYSsAII1Dhu9MjIgbpA3vwV/4eR7/fwfw20QuJX
Jf5KrMatDIK5Hi3orOkR+Sgt4I6FGWcr+de3S27BjBl1FHai4f6HdEmgtGn1YkKq1pNPP7O4BhnY
cMBBKpcpXYEq28JuS8wLSThHEjZzJmMj94/N2NrRoaW6cBMPzLewNcETHcxHjMhuLmuJo1n4R+4w
qvL44kazPBa7z9MFtJ6ohAG1moMgMxiFJHL8CrcKT2p0vNJp7rxr0z6wEXlzyUrSwXky9DrbjShT
wBqXrfMzkvskrv0X4tUC2BVvfpkYfQbctpr5Kkgx7uDymclTo90zjLiWwCfdBTq2VnwxeFHhILw7
FrtH/Y4HakrcbLKnSXLohr0E4t8rQNdLavyssdHCgiVc873FNAnoQBwSM3PGST1F6lSeA28HUn9H
REhcsm9rmhunUw+3qdL3lCOeb2ggyP3Wun/HMHSuT27OF/tSyCXilhje2x4kj1fj+88l8jtCtnzo
Xh7OnzPmOddNR+sofEQN4B1PfiGs8INP2zUjHtprE4n910LQFAjLHTK4bTdAMDcISqGt8Fw57vUm
UFEBgPROBlYLNX5kyJZzZp9R6kANUeSsB3iB0GadirlXuuezVIyqwsqNnQZTYobkngD8vm3wn5Mj
pA1x1RTbp0OITXabk/vURZi4Wti+gGlH8lRkimjKsBTFyonNyhzLnfmK9uZmY/zIXGGgmb5zLBPy
S+p8tfLKRNa/w/qg3ijSiBDY6yaK7lq8zKGNkvIrBIaqtVLxfPlKZRntEk27ouPNfJPBGxqaxo54
Ey/v+z7Hyx6fzC7nk2arWTQGTka4Bp0GAJKI2eLxoEnJ5yyCzl7wNETf/zIoqZr74H/pG2+sk43G
g+9Ev6tjcb6yy8r+1j8U3ugwRqonc2FKIT1xnB7cHDTgxU2KqrRi7ZPEv1A4Iej1lD4pR6fViA0H
1hciDBHxCEUzUlwpPYxITd0r1KotcGSVRYOJJZ9ia+mOkq4sRlIyiQiiQFKr2vM0lwq4x/MS0LVv
ahw9hI0PgWFO7lk/GMt/Aftn305qACmQjvvZIU+OeT8w6trM6Ltbi2AfJrRrVfqvRbzCIHgu2YGm
rbwOamRJJNBWn0JGQySRNe20VviNkWeidvF9VCMtFFwPYSmPzCJcR9xdQ634aYVbamFY6MAcbXuh
D3K/ozYt8yCxaQn3fVHhwZMJP5VAJW+mkWhZjMVknJpuruevxpS43YIpx1MeHfW1ZUUESOYvkE5l
G+CljL6LkWacLmmFbeJI1jRQniYHcaG3OjMGU5yWwFFBkJniu8qgEHKFYu4/rNGGy4bUHVMYUVFA
+MUf5zwf9e1zOyxDL0+13xzp/nNUNqIS3djjTyRa2PHo5XGLkEUTtZdMl90jeN3nW4aHLKuxOI+K
9ZTw+IbYeWRwisemK8QLB9hcs6TEfyDl1kQeL9urcLy2akmzQ1acKxUoOCngoN9NLP+Gv21HnlJF
R3A/qParDvAEnhZ5l+3h+96bgNOTPTA9rK8U1J9XVp8F5mBXflMRgXJVd4N13flHkE4XTNBKq8ym
mbrX+f1o+1EjvpQmSpW/62lBG6gF4E+cCuc645T/uyfmlUKf3Tb2wMUqVLXBNcLpCSmV5D54uJmN
DE6Th/pqgruabj5w0h17XymCrwWBPGgB4/taY9NC60ogLqIEiQAG0fsj0xF97faKhH3KPYLx2A9T
tMk3Pbb3M0fmNhQqOdA2TwConD3weuStOILpuzJVjSNhPa+KSSGfnzTNs/vD7+Zo5lRg4pCxuGIG
aP21f+Wl4ZsalxS/HXIya/jYrI8LzW5HvufHY1ecJ51SpyACO+7C9TNXrTp+9O/qm5p2iVEzF8n0
T5UZdZmao+TKnoCbQHFInXOmFKM9iLbTJP2zxd2izG0tNQl7dwE9lkyfJ5Wsz0eHgGEjr1jm7p5V
LQTXFNwFVnXF7yBPVby/C+/X37aa94Rn9GczC9WzqO/o/78mv5fPGboqJFaLJO08q20X3+OteYnr
lkWF3+2NMUs4gSfqHdvNf0EkE73FdLhOlQaDggFqR/7kESfyVMi4NJJ6/mF/aTBPnivzWdYkDs9A
XP8sKRy+kB2w7iYRJKhKLuZL3nZVwjgePTOUK+Rg+7hYMT/j2cG0dBxNk2HX25ccLMhX35ZWMYAS
bVPFWMhdnuKKxy3cujl8t7LNkRqif/VG98i+bCTPxkrWZJKhylF7uX7x86h7YnXS6KvGt7CVIct9
pHtgsa8+RbXZRVT8a+bvKA8Wsb65fqssZp7rfZUTH8xAoK6mU/nk3dMSIZUre1TONL4rNdJR8AQj
1AejjTj4ESiBT40UX+9Wl3F/ywLCGKAy23P/rztk+FaW59+iOBLa+ODSxzitbFQGCq3WvbxLw+O3
ZqCcL7YnWo8GQ/gbul1/bjRVDbN9AVuGzbXN2EpgaL9dr6RtHGucgunoZ/WUJ8T2GZKgsWDoEG9S
Xs6QLjh3XhYt8fUQAGKYEtjGrde6RDrU25TOTXSCHUs7x5zBqbMDatXmbxvwlGtJN5CjgMVPuAXh
5SgZ2CneEUVF7m5xtrQ0RlPT84zP8RWrSglzPN4CEuK6VYxWrU8886yMKFlc03MVltK5SJUGsrsx
lxonvqWrxdYrB9cbPPdTpt6OqHqbXW6scEY8fMmbwf2xRGI3iDGWh0d2QNXGb65awejgkLpr6RKz
H/9r/o3DQgZYcnJbQM/Cliw5GmPk8/Q26C4yvjG2D8X3qKzuKttBXKsmOgku7JgYCQFT6EilorN0
ooM3S9l4n1JPMqKj2SIiEoXsJSdYfDYMlq/g7+hpiT2IcoCRo6HHXeGINbNT5Z6oX/C4kA69mEbd
wHyAkVkzfKL5WBPLwa9nX+jxIgR6akJUqenDqhHweq/gv8vAsq91GOLUy/kpj5UsW3wZix/1HJ/1
l7iPa71BU0Uo4BWeoK6YGf7JJOcQX3F/VRbD5namoFB21g6zuHmeDZi9myDgKj2/P6xpHzEk/lV8
75Xuxy3pF7okBGt1tSa718UuNXtEs2RYJqYUOYo9QKeAFdZMeNxe3gyaLTeX3zVxDFPLiDtgJql+
pvvA2yRvP5VUMLsT4iak/M3ukUxSHmYnPtU9tYx7T2CnvvhH1mQOa5dehcuwISYgXQJ9hxjoO/0B
Za2SXI18OPeD3V/UgDAwypHf7y50kiFB5D/j86c/m5v2iO/I8nL4Gam616pGpKgc+NTCqWDHlNiJ
UKAS7/lg+WhjzERZqvqDFMdIMsgWrgrIB0QZumB2ezO98aiUPAlOB14q8GOT5AWWcIUJnRPo13oO
RcmNc7TlkRVlCa0PQEd4c+UWAX8YVHE5RbIGDDeHQQJr3guBFQlg4t8N4mT/UtbGY+QfDvHxm1ek
CVeU8813RRg8xS+zrzMn6RMAjH/poTOLEvKNheV1xty41OVOzB/K1Cd9nasI/LhRoAmKYPTnImhl
nJUNV7CcNlyOTMxRumli7YUzudfgumsP7yxSEuOYFGx1mrppFlm3gYqUHCZn199Rs64YpzP9C4J1
JB+LG5cJa5rLPhQOKS26FeYgs73ErawqOQgjE/hbaUy7adpTrUU6YHouuAjX7jH5EZw0xHNkRZda
QTemfGGyQekn7nEsw1x8acapkBP9tIXXy8cHnFmfJgWxk65tCBpwgEfJdIuWahmJF74h2d9KU6yo
9ihM4ku8vkbXy/g4rGc+tJkEOrSU0QMlx+kx2V15oL/cR+cqMYC8HyxifZ5lbfwTRDY/q9sI4cE5
oFMLWmjyxARPi9h8HMj9RAr0C38IqE+zMXdrQnBGjt8/l5O+FFSsinaFoUt7F3qEO51Zb25bveVt
hq6kQhqFHSQFeUTnOoSB7j+N6fbyDRPcr2H6C2rcqVIj7Z5OuAZff8UL49U1xYUK1MvI8VxzzQFN
LV/CH7Q45SDAVAVF8HzsEW2e12HK7nJljdEDCCHi6jn+ozspWlLS9ln/1QdI5CTGpwF3Z5Nvpncp
pLL6Egr62T6Aglwp8ZAfNGtFRssi1k5P/NCiSKdPzbu1m4dylUt6dGzSeuRL8+6EAoYCgABvcW5I
ER+1El22OpIWbG00FU/kOktbN85CMLhOEJ+L4OpVvEzsSTIbbE5yW2myoi34GVmvEGmOvT00AFCG
E8u3dMEe0Pqkh5RGdvT6+vCa/qD4uJiFN73lCykmujq0Whw7ljBC4jX9uWKeHfJQLHyDZoEcodvb
G16Y9Uy/H+Ay5y3dKOKk/U4VIzN8iiqeJA/2k0MXwRMinmXoaD/Ba/3oyuq6NJbIT/JpdobK45yy
LKF13c5Vm56o5auhy0QUwinrvAoe4HW3o5wcOC2EAVqFjxeKoH6axKNwiHJ6A7bp9Qy+3KyLmv4R
+yhYkWFIx6LqVLY+kNg4bIBT+Qdn4ccGyn308ytKbmoF9B+T5tge1zIJPJHuJ0AZBnIrUQzdWMJ6
sQdIkXuciuHmmsnwLmBkYtW/i1Zst/AVot6BzSQhMQzKggKz4eBDCmCNcl0Ep87R2SfblJl4w4sL
gX6S0t1xMf/LzDsCGFo/jxxmRgsv8NZByMEJHkLNO1F6G1doMWBcJCMUoz6WuHUlm/sAayf9FkHI
9NocoXjsZuzafYI9weY4RQPGJoisG3AlEm3Rd/9msTyHfuuidvF3nxogveLs+DB3mptwb/dsPFUo
APLJMMRbuPS3wto6qa+c4UiY3CRC6xW3Bne+LE6B+YT8eCRNQo2j8XB+ktgkDmaUej/gA2bbKM83
TbPmdxKO5HtEPD0DN7KDgXTQdYWPG5HRDtxw9y4gL3suEaFRdWF12EsEuRFRqML4lN7OsXlMi2Jn
PZ4kbN2hdMa8fOM7ihVZQIYDJOndM3c/Es8Pr03TtXnbMAkbdstC/mU8UxbTZqmnLolhTdWXLTBF
Q2k59bC5g1NzW4zMf6zVaM8f69smHccu1/GZ/5i2tvQeAz3vLrwPKt8rY9NsT8ZbM0jnfdB1L++9
bq+J02FSVN1fa7BOl9atwttzwzDzyIaxDwrgbbHHNTvrVJnjkdLb09VdeTUDqGVK8T4YGdoNXx+B
xZHOeN31ZJCwD9Vi9e8YTzjsaY2njakI8YLmfOCqj6OV8zo5sZlYfsygqff+YkL4/9S5pDTcf4Ni
MUSWdGYsafxyjAGk6Rsedjg2YKzX1UoHElLZ93J5lvjSCQZRZqT5HFkxrJQXWK+B5sEHp3mW5bWO
qg5xJu/TTgAYpQCGG4rHHGwibhlMrITyazqK9ZEOssyHfEQVECOdQXKdLlW3y/xlLYpFee6Wksya
05ifSgtG5zsnfBje13YsVFaZEwpaM32Om5+hpYQ2Qbn2VYEpZYoc9+roVhSBOXneKc+eLS9VNlVw
jesrSGj+LqhiKhejUfTqbLLLsHqbKGzQoHKkQaHWmmhqdwIek8dIM/BqxtebMlRzXWERJaC8kzrJ
1DiX94Bp46PxfkCODqi355AWU0C2E5IITQMkomwqii7rxiphlOegaa+q4iBmO3WKnz4P+Njta7tr
rUYZ5BsrMctIkp7plRCoT/9wXdkpEcjIgYbGfg7s1SpCEl37UQXT7E0g1El12tdz5Z+HzVAvO4hK
4do8941BXPDqzNl1v1j+GUTw0Mce/74xus2lCIrYmdZSP6/xRmi76b1adN/rmWf8++OipMlQ5TAO
Blrn67kb/NCaWPWYOXsyXFIdqQTXn8FxZmjE/pm9b7ug5ldKMwGTXY2kqixzMrqnjOt0orR4ouZl
Tpn7Rbnovbl0ZFyyB9t6SxtRVlhyz/VjH42lmchHgbpafpenRvKqZ8Ot3i9afzsfr4lng8J70jRs
EV4iP/h46G0rEVQIX69k94HMy0pKlDASwZOgL8XoJZCY7wuffr9W26TtqGYZ6XaMSh4wePJzh8oI
NmgW9sRy/HsZgmx6ldyauPHSTlMWcX832x4d2CFUL5PuFla/moxnocxTk4GIEqzdNYmlQZs/UaJS
vMfW4fpSGOMyZNEZXklpuOa9MEDMRskkllDMmt49KDPtuWq5vlA9vgVr6BymNKAr/u23Q5+yTBWM
Y1iGCMsXo9PGiRfODZPIEiKKgu4dxqGmTgQAfM84cngAygxx7XRGJ4CaeVuW+RO41pszAWbcTGtH
lI08QyhgyAYxhkAvPIfnpLLjXQ/QdBXpt3Lp5Rw1qF6lamyPVEYap85Dtb9Gsm5mNvFt7VTOiU9e
KVbogqWMywXmjUFWvRuMslyiFCmwP7DFqdoqC8r8vJZbKK3xlYAmBrJBmZzQ1Tb5kdAQpyNBK7LD
b2+M6L1Xtr/9XgtawmRmpaSiGERJfH1q06PtcP/5SsNOxE0tp7iw7RKRHFzka6ZAiOQSzJX5k6Ls
+bkxLWWLJ3M8sNL2T8HqwP7yARFliZxeiui7nq1HGHGEdJUYPKcP9YZL5ekf0MWawuBwivji2YZy
tAWfBookd/ZZK/FfJ+A+f61b97tmh/8AtZBs8HoPmBEGDaBPNB/H+TWpUhvLgr0SPvU2FI0G4HqW
HutY+a90DQovVOIpI560dsobu47bJCuuYCNyFBKMols90At2FvQ3Vt5HjHJeLHrjZE2W9GMRzHtz
WW/1TaHRS89Im8PiWenCqp8dnvS5YJ+uriIoa1fnsDBg4Wpg2yyT8VmZfK8r3jlasp3w8cInEHn6
3iez4yy0x6NFJ5+UKlhYIB5kHe78yjEwnDdcAD/BPhRyfs4cbRL1Oa4bK9vTa2IgjK00EKWrHO1Z
xpm12cfpVmQ2djtLTbv8wra3iudhE0y8Pxp2i1/nWpKfyYcR43z8ZNzToZDdO+CQsfoBzzxI6QEX
Ia84nagfK5EgcYX3APVJ8a5HoPVmG772rV73Y/6/+/l1FnA4INv5YoJTh1tHwGCLPKJ6NiiPf0Z5
hstFJIpg76pZ3OCZu7/ERLf/roy/n/uAO4VB70cVPfPdNrzAIaK2xtiRS7m6aO7vZvZh7Nb59Avv
EWltOKOdlgVb5jYSMXTwB5e3atFKmHNQJdujEbokliOkTRMfgL9AQGEI+a2KEJqkAQ8McDQFkclX
9TG0a9rKJ4WdAdM8pMtbHyzdZo0x0k3Nl/PrQky+kHDdD+licDIm3OT5fz65DU+JW0uGzgHYJuXz
cqWzFueCh2E3MCWxbEFtf2hQaJYUyHrn6P9DUdhrBA3MNradTVGNB5bB6BiOaGsc5jkbaGsD7WZF
iOf1md0IgSmuzPpSqf2UFvgeO+Ixvyf7Y3ftzsdks1c7mARs1kOnLZu4KRzuNM+cTdiAoEMnZu6D
lTrlWMcLsGCKXJpWPzT/FJPhTBh4UT0h5+qsN7fYMjAiTdcKzbT/7q/T29y/4ldWFWsLl9V4tt8V
4oDN1Uu02mkvCH/fZwIRQSKISM6M6dwfiYXi3ABnW3OiFKSX+ksJMU75PLriJFtam/yqeKYxkhSX
XeWqdtR9PqPMOTckPVz1twUt0zaPxTOifa7G8UtN3df5glrTfwCw76PE0lC0Ep7T21a+HsXSff6c
I4yPD8hMkS11FKEGonXp0VmkbwUFLQicnX6QJjCUBZCrsK5PcbToB3dRQz5UbyqLILx1Kgubc9Xg
/Bev0azZin/TjtoHn1u1aKdM787v1jODmRP0tmvwWqJfrvilL4NRrUW/YYi4QjXuJMhgZaH/wPsH
QVoSj/prrFe0uK1wsqBivPwtqpLynFwxUwlz9RyKPc96fxJ8Pb1dUzEvP7n35DRb3id2m/3QoThl
7GhJ1teC8/XwlJpLVjdNK+n3dqS1GJDvbQ/IJnt3zlBihBK+G1c8SguewYZwTcC/dn6afdZ37/Q7
SnyakMLS/eFh3h02O/Pz99h5/tYAskEEzDkIWt3ZuLWg564YXRUyEwBgmIoveSaruJXRgDXtlagD
B+Q76+2SBKkOH1QoruuVbInKJXcsLOM4qS4PfTqAJfWNQF1/Uhaml5cBTmHEIv6nnD1aThzke9Sy
SULHpErWgN4owNRH6AZ53RaGkKG4VD53z0THsSO3SVUHRZjLGUGO0yg3yg4yiS92rQmKyYJsIzko
rsOZAREEEzQ9OyNizQ6pphSPP8Z5vImMOH/z6R+mov3xAIveI7DCb4juED4SDhSYXYhYpd3NoVy9
VEKrSwuYN5ZNYF2VLCZ+MOkxwQyH/8gBrwkgdyiwzEh0qa3pX7ew4U6ljTltj1QHxeogHpbWfsA9
jfMXGNhB+zzrFPIfpj3nh6mNZvtmFHb57D57p0fIaxGAKV+tUaC3u+m3MO0QdFELnQosh4xeh7Mq
pOwcHyzssEOTE+pb9jo7WxUyjASoCThNDGst2JK7mPzud7C02lJOrd8eQb7cXei0uJGZOrpfJQZb
CeIqE5Wn4mB5VIHPoR3rg2qpke7gxMllAgOA079ecyaYh43N1Nqs304dCtjFmE5lGcOTllKCCkJW
XN3WZmQ2iNU83Opm6eUcStGmVQ2l2LQrXSZ/tpL9YME58w/kUkJgdt217bimh+TWwETbJdmSX+hB
N6fOYzk2Nt0+xnhc6fxoovkcLY55q2IbetRvaYuzXect73BmBOVBDXeSSiZmdmqNsTj82u4YF/kH
UnNWcu0V10g+Q2Va0M3/7YpLsnpCvLylzAzCoRvktZtxj/ZuE3u6EXB9t+zbAGkCg0ZHcx/kjfQe
BpRQqa4pcOd4bW3VmsAX2LrrmxTbnljoNS92nkfBHObTPGQ4PVcxJyLTtIIYUJDtW8qkxrQbwU3G
S+CmO+z3ZE12CoHjunY/o0Uw9BQ84S4lA8jI9RyDwrbEDw5+lyp5d0f8HVpxHBATYti1Tj971IM3
Jz2DtoymogY+PEI5rLYn4ORXhTl7brgOmlGwHBkf0NvJxv1Sp8jIMnIFAH02Z1es0V4S7wEy9F6j
guk6KxofAh/wjl6DMmVtAko3DYMITq7FNS3h0XJnyHmTClaLC0lzaWsp/yijA4IhnCmzFQrgRRjV
+vcPNA/VExzDU3mby31D3zU7tAZDg/zjoA4lst0SoRgtig2c0PJ40lsNFrsEi7KIpvdU1tgYyRl5
8qUqgr6uFrN0aCvT9o1pDpJkPsptS36G3Zm6bZxgjwDLN0eM/BF5iKhbyCYyzKK8hqsmz1lJLqu9
3Li9XvnaDbJBBvvllSKpvdaGMBRqNLBhj0xUAwSAwIO2mXZmtoUbc//JL5YnxVjuZ420FliF8k24
8hiayxZ/HrwJoHeubSuJmE9lPsLmq5PsVEohtVwb+Wmi5d+B/DFDBcbe+QxVJrbHJKEqpwQzc2wm
YQT7dKZlPZwrIb+10m+aLXCi3HejU2reopyJKFyiTIwJMyAYSxF7lSfuI+bRdfqQueHOVLrVZMS+
BaAUwfUJWSDyA50hlKKl2gCbswG+ZJ7sTkgkjOMw5HKhCoOGDC8TeU82GDrtDRn/TJGM1H2BPx3G
8vQUCpFCW+Krh8cxWQzAc5JyCjLDlDvHfvQUZrvO8PlOHkYsvcq+FvU7KkRv4Z0VJkJjwK5SLzPm
ISDUpwvzrZ34i2QhNvPz5nD3cEOWMi4bvbZGpJXE8K8dcfGa7qsyaTxVCsCHQ3wIPcrNTK6klliA
fWF7SsXucxvOl4H7C/54dQ81dNYJOzGT0ReLSW/ismntbDpgvCHYoUUQ5CNeY71L5sPc/HfEoGK4
ljqiLQuae/LAxNLTWNeBBk7yfNfEl0dqB+aT0EYKqNH0qgWGCxrbNkX+P7OqNKTd9J6LqyohyFfy
C9M4mDOmTlgAhAh5ZIl5ct9DElTaB/iVrYTKzkWgknISUzrpHpD/8QOlnDdtaFe8/mL4tWQfh9+X
F/MXYlaswojc7YXQWY+3EGHxu13dWoNoWgDwjFXEE7ZCI3uOsy6pSH1+LQ0FeNJ8/aX2Mq4ozx9Z
6FK70MPlmLINg7y4K9Ys6zLUeuYfEC31tfPVnn6F/yA6C+kHB2aV87UZqPFLnDMli0RpQ4SpT06j
4nphnKJLRdE/ecocG79g9JFlDJPq7siri7q74UYA5VYLW0HzT6Zpzuz1jkRjvpctmfsTTcmRAa3Y
62OniQ5k2fN8CrYmzgy5b9RlFOnjvqMI2WVGrW0XTZCqYXaNOFFVD/wafB6U0u9FRqSM7p5UHd/c
ikDBAFSWEI1ggmdIFV8ECcSCCwJSu84WQiJnRc9sk0ikHOYT1Hs9mfrT6lDi96F4IjpzGiSAqnyX
/RCP4F9r2vaqB5odVKV1/Ga5LB3jdd3uvqHt1CTmWXr9QDJvvK6y8hUBG2KkXQE2QXjgFEt+LZec
1ecQVWAoyF/k/2ByDo+HuxvRmtgumANicpPEnc8imTEWXFvtifI6o0XUKtO9S073PLhS7/qWAceh
IyKmDfLf5vQ9U7yxalkrn/AfesbDCOnVG6FyDXfggNm2rbdvNMZuqgFtJg8yZowTXsAA5ICoN3ec
Q28wjhJff0V08X9rgDVylMHKwnGSj2eeO+udYnWoAyDmB6eWp4gXgvEaVSKWI2e9V7U3N+DF2+SL
5/q+NncSNFCc5eXcG68wOWDLjvCMyvNtIY7M/wo80qAdlTlJINo5V//X9cibOBbH6qJE2Y9IdBFw
illZ6Ko0BxMFIg85WO0z1JptDHKSazPX7ORVzkKXwFF7xHH8CUbjhD7r7Avt061kM1kSz/5qLQ3U
8sYNso6r+y+l7L3sZddyuvLRd2S0sMurpA1fgYKdipDvrRAQtcnLXwJvSsmkR8/LJPkc5ucswi0y
J9klzxTY3B7gSsN3li5rdoRe3AP6nD0g60kI5XF3DzEMZ4e4v1DmJqR2q9l2gKaCAxSAdpPVmDJE
+S45NzztdhGn0sThkFrTz/1zoBzdUpbD9brpi44Aza6pm6x28Qv8/uYCMLcYVJVZUj2iFBfuu3Nn
pGLZcTnlfm5AAMoXi1wHvq2PCgLaQ3SIU4a0JF6UWkoP6dlRTXwettB7V//GF1igJfTy6FERikBP
pXBe+zVADKR3X0Xyq/deEmsho6BAn4tR6WTN55FUAYm3k+sO/L/Gko5zbiR6gU6GJnZabWH6PLXj
VE+ea98qmGh8BcPBQCI3j1v2em7KbOvxeVbsaYcCxhgsO+m30D66g522cF8XS2Ua8cj55B05lZIt
JGNImjIsf0w7ffRFGIXYfP2tTPpL7K0IKC6blcX+/0p59v5G+zFJy0mpgWO44HUiF8GIaA0ewj3f
c2L8eCWTGnPsWXotc28USWuoeq5+Nuq1ZzAM1DhmU/ra60PwKS5dgGe09dmMoapmidIGFK/pO0LB
4lPTfB5orzASdmSi8sY5sJMRj8i+QVjSCHhYuVHMJ5C2Z1F0miiH8qhNPTV3xczRi08OdwXXy7GF
ZPGqxV1GGwxnXcJ18dsoaW+hleFoHEL6y1v3YPp+b6tfdRMFhZL+yZgNcsQcaXNGeLD5TmzCrFe0
HhA6JtKOKueK9GgqToil/IIY1KTI0sqSsNTEKtIEwED4am5A9ZdMmfjjX+ELdoH5VIJ1hzfdDFHW
z4gCefDKmROoAm0Txb3ZEbTfIlDJ1rGirchKALRsf+0j/6w+Q7LQvjSglcaBqYsB8+v/OtqWStGN
wM6ENAB5EPe8T5DXN+cM28IfdT4NTs8+qRZ4cW5MLRG6RznFVZ8P+zDTUroX5M6VmaiVvxR3Qyay
R0/kPUPiiTVdNe2T0rWxivUdz6iqrn8PB5/6YvgDnm/QOLxKxpaB8JM5IkN7q6UZ75lBtYkpsY0A
AfbbgWGvGrjjbl0la4z6oHd+XOQXdpKmQQ0gM5JMG/GaBe/2fSbOP7ehxYqR97ShrbJRXl6N4xek
P06UvsAyFvMuS9Lgkk1jXsVuw4fynr5sCs59LaPR/fpt0ftQXz9+SBYsIDxKqqWHR3d3VQF0BrH9
yScyiGokLswpnhbO5P7cJdKZTiHZZd69o8wNWtGr5H3BTIWv2t4eZzAbSYx6D/Vmz2upRlYNBnua
92e//Lm9iVyswfyGfyclfwe+zkfZzqVbgMOa9amh5hg5BTNwJmkOb8eg8bC9wPLAmOHwYAFZKV0H
nh6Yc3sGV7nQxQPnXUp0FyfOVMmLw3ghDb9YIMxhPdIVvyAXM0rOAHchNc3zNgb1vj6WV7m/GUm0
R7oivRFStCpuHA5GJStw+t5fnGDa1IvyKmiIXFOS1/PGFbr/r5JXqplXL0mkGx2JiViqQEiLqMfT
RCkjxam6564oJ+b1rp2/5Ovk5v9zG6uHE0zxQzprKPM1xs10y/EQeiceXutZhYtRYlNgY9aMUUeW
TUi3XdTcebizVocYgVMrVghLuaOrVxIrdSJzfr/nr84dTPThPlacWmS11zxZabj1Eo2T9XUdu3EA
SAbO3dFk95g73Soe2r+eHNz8rUDErzxjlSLvLoM8r8s+5Y8VK72pxd7OKUBUgZ4wRza70qm5Tb3f
jNYa+sMt5HwpVPByIH/gpb5Rl7sDpTh7TMfyjfIPrDwRBCHSiIesZXecO/XGVqbVTgSLFfInjxB2
NfkvBMd0Uzt9L7KvbuW6VWGO8So7iNP8pKSpF+Obk/p67xEnKPzV6191WHhFO4T88mtTe31ahc+I
i8Rp5u1Ukdge1hKK74gjjriOobnnK04wJV/XaiLR1AuzVeIgG84QISb4VM2Cd4kYwPr0H/8CPRQB
vmgXqDxQTAJvgl04kyqLKg+UbXDIvyzxPzEP6fH/Mndt0KxWLnShKoS6OCRkH+HWUZNfgyMq4O+7
rhSEsHV7KaG9XLID6x2WMAuPIo4WnS/RhTeOlUqtjNOQDfrtHu5zXznjE7XuMfEEPIkzkfHlg33P
hiWyKRGUIlvaY7DNkLZS5SzDS6gsMfJe/gGwT2IUnSYJ7vt8MordMPAHgUEBYfd2bhQVrXRvBBoZ
jxYqiKOefrBA3mg7Eqkcr9t4sQFpAx7hHvQF/+R3cxMIuWR5UBH6hmPGBErK2urMhvJHCLBaEqR3
A/jb8Qgb5MXfbGWNUIbFOEUyGPiDrVl0F5fapcFL8z1hcPcG7FWpesoO9ha4VYJfpcDs2BA1CV3/
NojhPrw3mW3BD9Tn8s8MQr98iC6ZhrB8NA16JaBVNLcYHsfa5hYRiFrA9H+2wiOBsPCiIttvOotP
QHKjP9ImT2Gs4NgU59aNCnluedfzrL1/nloq3GhFTfgW5PcE9hmkv7NpyXcAQH373bpfwwyHl8oG
KwkwEBnsr+olt9srr78l/7ZR2Qq3WLFsG5EsqUP1jWjlMvvm/j80hznWhjhl/THMFqjEmgoYty3K
GYhlq9WYPtqBsXlD6JD7UKo6tJJTX01ICN0AAClFDFN/opHnTd8Pvljd8vcrBfDX7QlSZ6lWuaXG
rUnQkLaDVlctOC4gn7Y4d7FOD387H22yu70Np9P53kJeirZ4zgYqZPHWJyoUXSe8+PRwCLnNii48
yWwBas4qHOUtfv5ELchBNDFy3CkD9QGyA0XiMJaFB8gDfadHZNx2QwHNlFWE0ZTLEPRJyIfYeNtF
4PImCj2nhocspoohfowfO+Piqld3oVbF483RUgQI2Wa5SBWioSVbDgnGjdww2S2677WLpJtJJ7yC
cCvwE2xO4zhvpyZDNTr5ye8QUTwZUkk94QYlxZ+diCJ4F6HduYpM5yFFyjH5v1UvPJzEdRMYsSE0
uu82o4EZ9wv1YamDrqr4N5exXCq5iyhBL7i/Y9wPa2Cb09EAoScRnSdritxf13ZeWKKoT9wj2dp/
BFB9W0+R9HDzW0MNEtpTS/nLwSdKbicUSnfGxT8M2AP5TZpde+8opBsxcINobZblFOkG5r0/5797
a2TFtWag3xfUs6szi4u89Ud53VEYAWrGVILzYjs16eQuqvs6H5ddc9L3zepdgNeNyjl+PMmoy6zO
TykH4ezoG4+tETylzz3mjVqPoFXMvB75Q6JN422N6IJx5jtoS1/M4kUjtcQX8rh+KuIAY7zHN6gc
mZOfFTkG07fS8u9OeSiuCK/sHxqFJvONYXmzSDqqMyCn8W8maO3tx3A35YY5i0SpXND5lLQmbcCh
B9dsAF93VbbimPuL69KKMmlQ6xowMOOfV5DYHM/EJ4svtvgMZQZI1/aIMkkzGMRN0L50ZtuyXhY9
K8QWvlIb02cOAgb9JG1Cqj2EW8aquwfObMS8EbRIge+50YjzIArfG/1jlSeDkuZWsWeErj1Jth7M
X/SGZ7YXfFjgT6N+yGlqdWFd38E500LS5FF7+/xl1JoFKK5Znz5WWM+VhS/QSiMPAdA75pb3kcyA
OPx77UcItadmPZgzvIjtdTAWHNjGApPLI311QE+UigZ4VHaMS30gU5ttFzK6PHRBOr3sEDfOSX1z
RRh0x6VNsfdRMRPtiA4L3E42dmUv32L6CxRevi1ephYWxGfMqeu2XHXUxdp0O+JxBl054vYsgfV7
C0bJWL9TLjG2WyV1Jz7y+3xJnwolcua9zUzqBXzzUR0KjkNjqVncsJFANcpHfKhy82LCpkToKQ/b
YP2K3dc7rCGFxaVQw4Ck3MGJBTXgWHYx+RpasqiFmW/VBGNZ6x5C7D//MimlaGV0L+w1YBW3aHIf
cNIDsisFaHtQ3k4/IgwuQwOA+TcWobQMkBr84PYfMkxs+LmHCNZvsloFaa2eTXBXjcLk5blVBJrE
3QEkC0bWH7lsy/iUsXrr9yTGdXIiTMLjuntly4+oroyDjXR44s3Uw7oZ0nt/1M0jXxhqFVfLRdog
DOOAvACakMN1QP1M2w59Ci3IGtKahMRbxyJ62iexTDyunqUD1oNDrpMFps8djmr/dplp36xZ9orY
Ac/KbJSplhWHNA728JKomKmaOkRg5vfQGfwLHTla+yQU72m1+B4Ti1UW9ko2xXw/5Pkw7vR/d92D
Kk3PKTLbZ+r2+knD5YBCbC2ariVk7iRc0DGPzMkslOqDUtSP/YfCT79dEGU7Emgg8FSMelq7OzQ0
SOrgNX5Ztbux+lB+n18koHN6vkB1eyNTtg3j/DvrK4eCbIVWJ8mNZhVhgET5KjC5T5E2c+vGrTmr
IBEO3ZCoyJYx14lHc1T9M9ztz1pKsXTpdW5cHVWpBcfLRBI9ngTSz2fTTU293pflY8BCz8Vh9Ts9
wgmwLMzCFMeBI74u9OX/vqFhYSaDBBAqjvsdndDiIjVLSvQVrX0yHFTosfJWUm8wEEeKzls6OliA
EL5h+A1o5vDxzKBy3wtShHGGye95zCP8jnfGvXcSuBXu0rvQ6t2lDo0gaJeQND5V0kHAsUu0BKfN
nCRWWuHfT5IHcjE6I6ntQtYpq8F5tajkzfmsjCI6nR8po+/5TkVVcQJUP9PoXreb6/aEuVooJ8Hu
iDwmyin0DvmPU5iFTzOsjvhUCKm2UiwFMIWhyOiE8KKQUvpy9FBEwPTfZ/Yzbz6luH9SuQgsEQm1
7XCr9JyNZL9HhsgnG2hIxFMHrkXwbMEIcWlJwwSOMB4ITnDcWfzks3Iac24aU9NYLJ7wMLTOQruE
setctvBJwBj4WfcBFOcTV5D/W0pRQdT+8es7d9IIw/hcR4nnW0KES7EpjHivWvUkfUGbMFBFcVOC
aWOsuO31kOUaV0JWvyYUu1hhg6LyCRs7sYdF9/4s2OxBrbVgEaaqnYOn/aGmGQntHR3Na3DOBLPC
Ej6cj95OX5KmZ+mwWEsw2o36xCp8IIe1QybXjdBrxX9peD+YjrnOze05LAO4Ruau2pI671r+bXFU
Wp/Ix0D7xQFxbFRfjCnpZY2EvVYjzf0LpN3X0maDzQ333w2GiFdBJgI82J7jOySjyk5iVQ3FGFks
i4VVepugatkmPqwpOmINnM4VmOKX7czYW3yIn+CrvDSfc1EUtLJYcgjHnqat9/ZCYS2uiFzW902h
a8VyXT/tMM92RTdbzuAvUaAH9xY/T32NCxTGbxYNLsAoNgtQhhdps3xg41TVHOEy6A9NFPAOiZCc
lOH0mTsqsvKFIU3eJfnYTITPdiDe/dVvZlofiqLDlcIyOMh3DRS1FzZ0CjIPR0dd8gVDsvoZxYU2
caTngMSv0LFlzEeYy9TjhbNxy+sweVbGYh7XNzdBOGl6nYPdFznrYiGGg1EcNyMDPsgUGw9sGgHS
835o6vhLAUhKPwKPcieQMq8LC0bMc6gZIezsdHxuyIu2vwVNMyXJk2ntdrU58pde8CEnJ5y7MZOa
w829STYSQxdM+MvNFsc15iBN4oy4XnpaLy0VrnmdAcPziD1MieOfzKcmhAId97YQ6Q5Ac7IdTTOk
tLqSE6Zlw15hOEdy7lewElSo5gabYtz0MC0wze1cBtZeQISSkHW5ccfzMWhAv5wPAtozMbEiBBw0
ay/9Wml5RT0HPn4NDvNKEY1R0sCESjM0iELml1TFhNDibNSS8HlS9IcFEX4Qaa/3lpCq3F6KUKut
SNpLMZ9Bln6FPUJBk62FQYDJ/cx3l1xHWEu4pqST7cXWqEFn9uzGxRiWJKznWG+grxH+iP4x6asV
KwTz3joap1AHJiI3C5NDxJX3+gXRIQdze1N2r65hYCpXyodrov89tkvyKC5afmyQFUb+a+0KJA5b
pd10fHYvh5jY1dPQk8XKiGvL4Aqv6oQNWB34oHg/g1eLrjlUQKVNFu3DgIj2VhoccsbjIcVwDuzf
6sHG11N+gzqpSN0zArqPe45iPUkbYTYaxa/XYN5oezR9kAUuYDZz4WnPlqzQQmpI0pLVhTkgsRGL
AubFREW7UBSDEvkz0y8+tBxDatlUMSnqHgj+FiOjClS6s0SY28pjiGF2Goz1GJ7dZdqCRITabaw3
9f1+EtC7wKjZF4tG49NUIyFChPeXs21e03LmClMGC/lEYpYx7kKYEbgpjzdWKZNlVAFKQLD770td
5rZ7NV0BUnw14gHVoUkilqytyjdqjWh15e/dDSjlLFubWpcZYay4Mvi0eekMghYQuAnXdaLIAIW+
dsyb9uvo7/XgjlF5KNM1Qyn+8Xd5OVQozbjZFMZnko/GOJdNRlFnoDg9fi/MtrZIEw0T0ST+gZJP
45uKBCLaR4PfXQwr5ypsBKCK5riJCd6A7klps/YubxjB39lPNv+B5t5zSFovS9n8kGUrazxp7zRQ
1Ig24tqifAPdU/N4VZVaeQjq11E2cahIk/RoTTphYx5o/oKI0f6uFuUD79U3iVy0c8FdeRKA7ihN
P8zqPo9ItaLLHOFfhzQ/yd9pZ62oq40p2PjrQgCD3tj73kOkV/3SfebSynVU4tPjA6DjyiNC82Df
0hCn1F1Cpr6sCii5fIFOXq4RLpzf9w/z6iRQlLoCTKXakHUEgP9G27o1E4vmOrss0f5+DJRYdAr8
X8DCHHvkxCEAdiU9EfmrSUTYyTVPAib6IYG4LUDJHknQ9wFSECz2xuFCRfaSffEn+5cl+VBNideC
8KBhlPO0yLG6xCVokJnQz8PPmUhhTBwIfbjgx7qH4vr7IY3ZM7ZG9D5S9ccexvhkb5ltNavqP4Rt
WpYc8ry0vD37XXB8DEuV1egnYu24vQCiZu+13heUg3Es8sQP8jWCQIaSbo+2K/nXPhTSz6AjyN8G
V0A6evzoiaPm3cU1U5EvZ2cIuvJ87rDGUhEHia3lvR31gQ4tnxKInVPtrNCEVCN+7F8F5FBI73is
WmkdecnmXdPagnAYBSENJbVZEetdfMcJIxLwxZYAqC0xnTdyoVbPwRIGzGil3dhVk9hOwaqSvUST
IR46RWDrrIcqjrS+Wj6NHUzydDpH7FafgBUnWQVzfuz7cuYlNroAAr3hEa1bz8w9lZ5RImwXIVSj
c29Mt6rkOf2nWTYlHNHwcE0NnrrSfIx+zkDWJhJZm5QBRn1AScojYw7xCmllQEsB4DpY9msWySoL
rYp1nYFjIn6TFD10cl90AnY+gFJDKmGv3AoQHUhPRr4APaboGXrhOlzgu72622m1tU4sgS3plTvk
zg5hafrTmBxqYh0ZgMs2fuSHeh6t1kHKrPy60xZYDqtMAAjowhkO0TALRHIXCl7tWRvanGyXp58l
YGGvrRtZAA7324pdky+nbLolHTH7Xz4qG+In+uCnaRfRS2Cs7XC3NBBHGfsj6Jv1UHED+gpLr43v
krfSvyIx8NmjAwyH/7e6fkVcIsDTSTKOAgGO2nc1fYrzM1Wi8iIniKLmpoJRGv0NthUQSo4SoqFq
FsMNXlFwhuIfQnZCN2cQjiR7DbYTFuxmr0Cfkb85CTMpHtIkpdtwkIw/ibUTQGaoohg69JlO1K4M
szoLrIblBocEmBQT6p46D9qIe0cYJCelM1QbqrPnN093t5YB7NsAQ+I5sMEwd1qnHsR4l7YC0fuq
zAjQdWpJgF03H+Pcc9EL+hldERtnAchI3IszXe8jDOhjsfpnD6HUjYPNwpx4fn1l8DOhhRsXBe5J
3zOyOmU9X/ck/0bmDEmMaovihwchjdIK06aSwkAADUF2HCbc4Oozw9469xeOTVUBRgfZ5eiGtMga
rYNw2ZpVqZreLivkgzA5ZF7Ngeli8V/E1IzVNVagWX6GQjzD2XoPttWFJ2jPYXAbq8EnljezZ7g/
wa/fHcV1VKKq26Y9ksw5okNxOrQesfEzZqsZtlA2MlEgTKOBqEuzR6LOS9h1QszzHlVsRjxs5GpS
k/HT2UcbQG4URM2VcTKNsYPrPw91oCZ7LD65DP97gh4tZzUDljKtAItP+gFsGkpN2Zxxd59lG9oF
Z+EG6LnN6dZuFTDT+rvm2ljTws6PHDkq/Otwn1avwk3IPOKfQIp7bUIM0+oAg8+kViYn7VjY7kLl
bkLfXO/Hm9/G6aBzdM1AQUZf8drEb0b1MPHGOpk1gyKi6j8jZVnF8RXMIuqAd/lkab6d3Doa4rck
m/6ukLzh2cpA43BzsAYHGipQP07vNTkWHiU7k2d/yftt0M1EqEYYSJr/dtjFNhPCg+lcluJyrfyA
3436JTlBghZDOVenPH0ItsSc47sXLsOnFgbN6KyKDCEvf+fywuOy/s7OxoHn4nBICtVX7viLuobZ
21GVW8Eo4MGGjzw2XTuE65o8aqts8CCboCDa3g1TDqVNXgdfdZnJx+spNYzwdTbR0A04SPwQ/h7s
khQ4Q61K2aRpBOYx18JXjxNpFnq7bpfjH9hoOdzAFLYF8OMzA9/HaIcBjjm5S+z3y0Mlzw/oEOyD
PchwONamnceXdssrs+1+Q4O/ptBwXTzsGI4ZSgHwohYSrgVTUcxiGfSTxrlDFT5k7y8pNudbuT55
7daR1nHlD8DDcfqjXge9bQTaymaJphOaKbGxNvZXyUHVR4Gg9mk33GopDhXziLMVar8sMn7bfU1r
ock0wrkPAXzCEpiIKpjCp/+8Ye6dGQ+YVcqgEqrKAl6U0KBgVS7kDVXKnRY78QDuNKFq7t4WOM2V
PTrYGtfDCSe/2B2gCt6Aa3VEFHhUuxyoOok/DeCJ5M/yKoFZXM/b5h06CBvL27JvyucUHvwv+mNX
6w1c3fyet89A1T9GnVXoge+h/UNV20bInf0q7OHZ8P2u/CRPWiSx8JWmLDX+E5GQM2p0Ye/Q8vD1
Vr/nEeWglkgkxKquEXgx92ADpp8IROwYDFcg3MBBzyzv1NfEdAVy0JY22m+h5HkRLg3YSceAlmOs
Oyzec7ETYKjlan164I2WcMLLYzbHsDljzsvbi8emZQja1YNNLoMhh0/zL9SOL67KQ2QT34hWTZ3T
vJ0xo14lrcn2z9Y2tX4utdob1/lQXFWB76QcU76duTs498J7B/+AWQJn0n87uHcvtEp27WKhbqim
6xg/hHjPce2z9SMdh61wuwYEB5guNmaS3e9SFBaQ1JCHP7eta1ciIrKH5o0aJQu0nGFBZhd0ICqY
KMfahd5bYa8t9FwmPePcCfLe12J1YWdQvOuyrSFASsEztbfjF8Z7jOxrYTVBUbUlwekh3P4PRruu
vlAoB7AvSGBr8VLpF4xeSWfe2ScmByE3iuxhJPnp61G4iCpi40GeSemR/T405Wt+vghpP3gPhQZq
NiK+gdcnBNg9cu1aflYpmA4VLPnI4sVZU8MUdg2YVggVAjXeJz74XpD5ykexYKUGIgJsRmd1JkTC
mtu1RaAwHPkMINtSnz1Uw6qR3sFn140aEGC7wPB7hAyr4a+gS9f/QAy4Q9ViHkRAnKh0Jzg2E2fN
t1CmzGOv8+DqVRfOZrT4TMCUP4Zk9I40A4LCQs5/l5ZZ9OJoSg4KzJhS7SHPs8wo6P29zx0ZYMtA
xUsqbCIgN+7tyLslcyNCADaU/TgoWzesDVkAlYFFIXD9afKC4ftTYKHnCoqzJWtTS9nSJaIE13HE
DdXlSjYyAWh9gHhQsIO5fb3StOxafwrqrvBBy7dywHIZsheXTXCl6i62FkGS3bYoqojk0IuVwWGU
awMy7/Cp81OlIBVm6gFIzO0vfj/+ZKFTuSunaTBkVTfbEGxiId3Id7lmRQiYWrm7T0GUW9OKPeG5
4QLI3ZG8ZO4uZmA1PLkohj+JHBJEOq2nB0TBOFmocjoF0CdgmGgxlNgcS3dLP+N8gug/X5Wb/YJU
pTeF/NbZaeQcGft4xo2fea/g0oTClVw1vcnNI6EC3UJGF7Xdfu4Vf8N7gehFh7OQWhksotIJimAE
f7No1D/STz8dLJc5u7aXzSdJ3YxhzwNf4L6aKCAfMbPgWy1EqQs5LGtmoOdAWN/Px8xqQ8gmf1rD
dneD6Gc3S3BaUe9113Nr3muBrvIGZmorZOHpqEFfltoABN8rPPXYy1bdaQ2v612mLDklqxT33+60
zDcNTFn02LcRBxpac3CurjBBiJ7C8AxMN5DV6iQiMtGO8iBA/f+tUdkVx0M8u0QPH9RC0kN2jJFX
U4md4MeJCAi1grW89uHgwA9YyZoJOJKV+hQGdiW0qoo2YVXK47HV5OVEQ0eaRljGfnkO1u7s+M6h
qDJ93IzlKVlzQ0k/eUQcfFKYYf5JbK0729x8/m6iFWGFfQiKcdD2xvmip4B1m7EZIqLa7CNB4QHY
geiiIhZ1Mbn/+IwFMPT5HlzBEvkyPwzn5+GjzSOGoXD91GdtDsv5PKAluBna+2X1RmJcW6UeMyph
5wmWxSEnuyvvD2S3SRaRCqJbFjzghruafvmasgtnMm3NBD8TbWCGyHx97XIReZoKShIPG2jGU3wK
R4DRp8kN8+fSk0AvVeResp4KA0JHsA6IV4/85NA17tiqqnt/h5MX23O/Jaz5aav4qJqo9vx1r496
w0QxeSmR3APMiCdFWi+J0/vDlQXHqTfezkMG3rfiYD+oKjH71eOJ+LPwVKp1AmfUf4Wbha13JwsQ
JhKyKEwN4dw9+Gvjh+jqKrqCVwE27f//nQ9VH8u2RACC66dAZMQCcHOcnEIe5IaCnTlKWm8VC6A9
5wAWJjBtVyaZTb01/xYwY04QXS/oyx9thVjJ6ewOD0MsNdmo/Bsqupgge6TbvXxnK8+Xo/OcPfUm
71qgbG/g9bTFsBYQp/frp+a8ze55laYYm/F8/k7Wu9U4Jr9kDzInN5W61SCzdYvPD9Oz9SHZ4ydF
PFg7m3lc0pDyCPtFSYONQaOyrhXpdWxiEvCrtzWcho4AlfRVrdsuHiwl+jZUZf60KYe6eBhKwXBT
QB68LxUVCXCWRcmS3WNJQHG044VRU2chh8SBPNCJdVgC95RWqoPf9+z5bKDnX++S/Dc1uC3zlJ7e
fvz5NVpqGizcZsZaKTEj05NbtRrX3K8eYGu9Q1gTeq6qzCw0H5zgGeQRi0hZwL+ga92AXm9HLwjo
G4ytBfvEh4PBL8B1gmqXUDzUNUena6CxbLm9l2bBw6FV3OAV6OyALtbxg6kPyklrGldwNaOG+JRQ
Aps+5ZWrY2XVZWSZjs451tetrBbmDE0/Zeekx13Z/bt2jmBf2tiNogCZsKwzklHg4bQrN4ECRzHm
1e1pMvccXnH3AIG7Ls8VzqKC/8IIGvlzkrUDXFv2OkqIfO7siXy0t16zscOKKQRyu2kbfPWGcgKH
TcAvsuReoebo9RjRwcx2lj2Tn6C/R198lNYbH05yZtFklht46aUfTL1cmkxWwRAB6tLXbB/oHsje
MEhtIPvq/wjDMe1lG7Wg64a3ocPkBK56B6n5Aqr2yzF1GtCkKlJY9L2bcAkKsZA5x4YFcortq9+t
e9AVTuZgvQim7R0e6jsM1qnBni7/J8eAOm1xSDjrOwfA4qduJlPwtYcBvFHx7V8bF4cm6kv3gLyC
DKM43WGwRda9fg8pwIGewA+gC7EShU8OXbGEtrsGDiekHCHyqAY5GPyTE5lCdM7ixQ6LjKTi01sS
I+FJUJNyKxEFucrCTuXExSZrgpzQnmCDJhxs45JyK7NuvdEBrubhZAyB6kX5lFJ4yVVGUe28dK8u
1fgbM+4wHDlmgHy7OqbSlYzy2o+V1fZQboi4GvDIEXlt51TIJJNOIqNj1dW9fMeng3vr2ownptGF
n/QbXbDOXNLs5Cs3b4AfYS848skmcvGGgFq9DTncrNph+yofnrt2ih2NUWQvZYHeqMaAaR90IMhO
L/4WkKYQftGvhGNNQEkBzxrHw5sz/igYFETdkXwrPfhb7tHYD8qKSoPiJL+wfBR6bOxva7jSM0Kq
NPxSNbMbzJsChQrykQ3Cwamoy89o4BMaAMFfTmm7Z+slGW0oNUFQbHkZCEz77AAP9D6YJOuFXqkk
mLpvSS0wKt91fi547ufkkH+cK+6KFZuMt0qyLlFL7hvl0ToUKxPFGDrLXM5kjS7NBim6IJPeEkaO
EfLq23mDZwNFZDxihsrROrks2zwIPKqRirINAO2Hjl3Y00UFuVSsz+jywUsJzRhAkoBqxy7iqh9t
ZVQvTfy0/m7y6xLjghoNsNH5PDR4XuImwgfqjyKznZ3gx8VZFH1uLWCHFC3NrqyaGeqgybo9E8Yr
1jQgzh2UjS/9UCBLtJMgrlBYks+QgA8SGFPY/YHCe1ns9o7FuyJPkl+AFDlrMRS+HKrLelbhlE1F
MEDap49nE76XLZ8rJ6u65P70J0EsVyXzsJnwYrmQB13uKQ7kdiZYThj5cq+yXcMOBv4SmTErso5E
CJZhomVmkpdJ5nF+DYlzGL19tjEzK1GAaYMkYMjbKXeyYkn5kKBLlBmDhsROUHxGWGGS4f0vPkIp
jB4UVVFjlKhPUQ7sLAwCyHKnRzsUJObClKiGh8SVVz9MnpaTXnJW4fhSzfdE/uflMYMaGNCDMgkF
LFqs0XhQwAjnnPVMRvMC2rQqaKa9qOPB93j5v6+Mmz0axAWOiEW3MSFavLeDmbj59lxy2cwVuaZr
6QWL7gXakpi6MNjSo198psO0qyIJiBJns0l2pZAvlJPjJp1vgqojenr9R8+TJoNaaQCVvSpG5w8K
y/nrUe7rMNzPMc7O54DEw79cy+tlWH5/hoi5ZXMgNu1Lu0odWNqZ5VxigLgUBJsUXbVqiBu/FP9F
syHtPjH2NBfuLgvrVUM+zaAPhkfRWt59t747MdpD29gpQCyzKha6MLhB87B09OKoBm/9qwmVq0XL
rsv+n/JSZZ4sjHySaGtD54NbUSZhwAQOphRGMFpiRQHm3D8vOpmJLukcHl4jzSiZctW5TOnGXvmi
ex2FhuHxxKvut6lbEa2uqL6o2QOoFjhHBwhe4BnvJCVUjFwjk6sdMDqyerNod8r5Sabu6wmmzcLY
kE3Xsh/zQkjy1PNcnsvAICLQ42Pio6S13UweXMM/zCPxDR9bmzfo4QXoX7NkyAueq0oyHiq1dkvJ
OGMknitQOlRiOJnxdmx9D9jFIo3hzq31lvx6QjoYAytJUl7j3TF/cwAlyMDzIXVrfjAogdvmzfuj
xkeWbmjc7rv/fQAy93itAyPLHxvyaFQVFvIPEHhwKDgv8ag2pW/ZRsx6U5WICceioawyYjD5t6Iv
71KgWpY1fisi6jQlbzToDMaibYSWUJQtUliMhwOGgYiprpxXsWWM1g6r/5PJajpcglNyJg+/QvxV
6qaLFY6UyMP4JXYNde16Iv74e4OoRqhxZN5y8/ynnajqZKd+BjSLFqk+RM4aurRskXKtz5/4I9Vv
LZoBr+aGMkTp3PLQsX0VRei9nFd+naUMVJp0hGQoPKoLyOSdHya/1oCGB7fmtCUrbROUX8n8RsvW
uslwQ6sAUcDk34hID/hC3IAWUC94I3Tz7Z4msB/7uttp0BVt7dolT/Accn5VXXah3kt1lDAhZBGh
gRRD5islfbD+8NM89ZuHVrBkiK8zUBcNz4kr59HNIyl4pcNjOvaG1EAmDPjB5pls5c68VrvCc5xP
ohqsss6sa3U92/eg6hyT8ZLpYgpCMCaw5JGT81pSZFIXieKV5y6ejDx3icV/4RsjZt7Sm2xMdc4k
o9bBrSJXCCGkzq81hbi6eVRcSaWouswKoG001vAIBVegBTJrfNrefXGenCWZG524Szm5xwxZntSC
UtYA17tlI9FVNQavLpUsYX+nDqFZI/JvrRhmUkRr+jR0u65AGkgzDw6JTWRDWQXFYg1Cw2e/Qj3S
Z3ibK1vVY/0HAw7IzSJivsWYQDNU3LG7C981QHEAO9MEQ/8nZAdVHTUuvox+DuZFW+EkUXKRlWJ6
bnRV8jiVEbBR4A5WapRvEuzf92fBjGDMBfofO8gzogF57URDzvZYnEYI+Ek99MBZ13uQ/aFT89x7
ByBAP73eg7WaJeUSPTzF4llJwtg1bjQ2s2s5Fxm3KET0epK3SES5UrswbKIH/BU8LGcc7paR6OnX
RChmHC1Zqy3WEBQf4KFI+Ss6eV00C2BOmUssAws/m+dpOxlK4bSpNECs2HkmeSHQwfM2nJODxcRa
V+TltoEVnAkrK1FUjcmSAhRY4gOj+GS4nNqtEBCG+coRQ8HMr1xw612B8G9y7t/LkwJE0Gw5/xe3
FvL1WxId210X9dSp+8BP5RgTEw1saT6QvQDoz6khC8dw3srAKcYCnaVypEv2GTS4X7ZuSdJVyFBQ
GgknF691EiDgOxHgm/IuSLS93+eZGb4TE/NHFcuBg6gDcQQd+8qxv8KGKOZoBSIosgvv+F/l9fco
6n0C9RFrXzZdneJhFFIx5fY/8k7zgxJKzkhLaEsiDu84vpesbLDKL1x8eignQwjRyxrSSVT4dbqk
LpU1fTTE4OK3WBGR1IYSliGugJpI6s6PuQnUuRXMmkWigw+jgQ5388a53wO9pKhg6dVDYxYuvAwI
3GXDrVr4acU+nGlLgVTbEst1BrErWzfQ/C34EvB6X3vYs0o0ws+/JgnenVB0F6WeD4Plqod+C9kQ
G3AGwxa9TJo1d7MO1f7WpVjYevpTLu+k/DKrJBtyX8okZ2pdmlUwfqNKB9+QuUB+NaWXV9yr+rLt
kgGW7Tv7UF67UUndQ7kVYR1458ZpKt7hpc8/U4etGAcPAEfwquf2GQ7TF/YdTyJH+w9rV2mGcVTx
8auAhfPMdy+Kg1OYDHJt1MHy6NTIjCRS/k4iZUr/refjSSsCydy/RJcQS/j//TqH0f97HVD6KrRi
2pBFPf5Ghv38ykruj3Bs/7exuV6kgiX5q86e0vDqKPxryz9lwMnIULxGdyOdQZd4aTdUhlOjpE+F
UfEt1d2+qDKFgtcmlP9av6+28nUQbLs89fZKdCLkDq+L58NtqJtxedjYQCbfY+aJQCGb4bt80bAR
HXDinMWuJp1Lg/6ftCySfcbHW3wUqNJRJHRd2ycb4KrXEuja9vFr6WRAujcXeay+tfr35KYN0WtU
NWzvJ8mCOv/7hZ/GZv8DzrIsqF2aAbnnc6UpH1ZR292VKn5njTh+tYsdIZUYi2Fl6Ag7l5P4lp1o
5NaAtdjZA2+NVESbRJtIBmNVvRrvrei5Onkq6SZ6qsorZHC8YZjantvTV0aEenL4yED3/tj64N55
tqCCy8ERiDz4UTYzcdlThPUIsrpBbuyMDgttmEJFauzj7iBSd2fuqWDhFvryAe45wIu9nwR2Ukp1
SF1jFRf80th5I9VxPgVj0O2ktsAcXUtIEzRvVoQe0+Z06InU3s3SEQFBu9kQyOGjfXrJakTDy8bT
ifLLeAOu5cPSzPYEGEBTkNKHrZ+c8KcQ0k33CRx3AkVA4PvXYD4SeqtaNtCQiKyaeQn02EwBL2CU
f3SNzgd+5n7B+FBz3JddKhNvm5MHJOPEyVvQCW+Rye/lPT2O4mFHCBo9gNVNoedVESreh6QM54zK
fhHG426tIu73McUS9SxEN3CvfwlSMULrijbSCczSKiwq1WXPJ6YhrFfOeuCoQpVaNZ6tN2vpKtPQ
L9LqHxGYXR7cWeSmJsxfsN4W6+BTDWED6xFwFEldKf5j6MdudXrKQtPYeXAm9DvFuU6LD97cOWuB
zYItxDB9/Ssm74Tq9RjTSHkGsykIq4PFXYFWgXz8Ji+ksW1rurYMvIbcZRKcxBjlRgQWDfw6Livh
JmYhdo8GVgeDyZG6KkJR4hqD3PMHhLEHj17aw3llAF5Jx+lCRTdUyctG/VlPz4BHQyduUR3F1a0a
XU0fc02pRsRbg4GvPXVQ0w+Q3T0j3b8qSY8pUGbwL5JS8zkwzzS/G+0uFA71WsgJC+4qACS5Xh0z
/5EbWaNeyGGN73FmxLiiKYK8Q8HWp7ahzaBJbKuprU+6lw6v9bA9Uca4uWPTMcOXjraJYCI0ldT9
vj1RiTrPz+6n9lklGaIuA9TGhNegzsIhnMpO/8PmkYZHzlMQggU/7x2RR7y9rYNvNC6yav4DVM8F
y6k1EWSCjgmep/6IssN7XzQLu0ONl6o6uVZsS9brDMfVT49IgVz+xkeNG848oeTzPbLFuuGXsIX8
2u6UJjQpWEd0jqL2S+NMFx7DJp3dUZ3HQFHNYxkTu6j65vEfcmV1WVyR89R7xjL00ESxtnaGxUbS
u7IbUxKAnXqIsGyh80w/RwDvzkW1UBkiZ2C3ugtyUF9Wk7Ty2KUuwB2tddctl7Cy6aWfafn8ZwjI
LnSLGYPmoLrz5YPgTTYs9dZ7ZFbfHps9yva7UfQIrafIu3pZmwJqvFaWMWLgq1Ta7GshDZh3YtKo
PzxU+3A8JmzdKMgMq9+xHMN7NYCh08tsX55hiqmTfMvPTB1nMvtLjE9y8wSuDRLuFzaA5ADIjAFF
+Mpi9IUc14kQ+lojDne/AEiUvEtG2QNIOFm+aCFTDyv+J22wFsAMneoHTZbo0V2P7ncKxInWLvDU
NWb1kAjIXf2e3mCOcmcM3z4adoidpUFqiwOReZ2+i1o4Bq4W9ReMDrgfCSkczdOwpZEUbvhETX+u
SeUs1LSA2gjwmNff3yVtFMfux+WENFy9MHO78Eve51qfPBcYEA5Ycc1C78J2co8wdLUZOisxucSr
NZ2ew17AFsLhjfV/iXSRb6nqcOT7HmTrCHoo5VNNWTcEb0OoXYsSt/1fu1SazBotMSGlfjhdo8Gf
SF6GCQR3WVSYn4go1T1gpWzpx8leh9sliiu+Weaisw90wuzPIslvejxJZdunz2ucpwLPhP5EmRo2
YqVQUl0mI/NRvr12UqeECDJzoDhDLLoGsWKVd46tNp4TcY1H1i8SkKwNW1jbSvOYy6I024oiZYaT
8FjHNvGlOoOfVlkb0Jqv4w9eMqelMucaD1IGEHGo/eanzSevZrSl81zwNBKDXmiC0/OCZRqPhL1j
E5gIkJD5B/e1pIxe7bb76pmoLMxT7yHFACIc8gSSqpafVVyO7MzZsc2ijAmPj6EfZzPCxQ+Ktasu
Q24h444XKVQw8nLnrKQy2W4imNuFTVa9IsarwnUdVJkLWKgXxIM/hK0nCFetRD4Q0Plnv8eKe0ds
QoFmakm2H0jHN/NTt2FzR6McP2uelX5nqYo9X3RBgjsJQid7/wKyEt+zY0Y3/f2+VoLKBoVKEq+S
5JAcJzqs2zqZa9tvRMdv/yPb4auf9xM+Ny73qjcEmNN9wvY28+4aq9ZXNP6WAJ7K3c8svVsQ7Obo
EDYcCLI37YHwVI6gbdstDH0PYU/2LS0IiPFQkVL3bS0NIcZSjJ6A7AmxH54JsqXicR0RY5YUtqEe
66R7juH5oFwaK5uCjps9UAKpy8MOd9wGcYIP2e0tEmroWyfIDFr5OSUSJ28LOJc1hAnBtiZc3cY4
UjK1lJQC+Oh7L27K1PVuxEDejCsmmIxFuuwCR4IZv+ZE4EgUVJzf7BJpxVUDulDXwtZuemaBqdL3
mIj60OtHyAdgrn9WLKmVScFrippsJm3LpYHuVa1gmWidz2ppESI3nItTe7IWhPdUtHCRojDZFZcM
XWhF0s8QH0ggkpoEMxTHRpt7Vxi29/lbeH0bv93aEW3lgPZmCJ7OqsF/hrCJKubL28k1T50wxIwl
S4rR0sP3KLZbeohUjiYm+pDfliqdas/eUTfQIcX16UQBmIcrSTzQP7psF6fa4gUF1i+ie8XgGVek
yxu/oOQxK2aufpBvuVGZT4mFDgakVyXAkAE0y+9KKePd2juTmEUjGphPIhqJE5k1AzvV2p2kvsJG
6D/D3WHt+6KMi+vciMlA/BtUu2ck9luWF1I8QzJJJ1+gplZ31t6M7LoyDnGEDADB7eGpencBhqRL
x52W/m0pJHHjqtv+IbLQ7kYd2Y8mHPgE1QSOes2Cv64XWGc3bDF8O67a4MwCRehRaB4k0LzOpDQS
dN+Z2z9y4cygn8esgR3q1qsZcOcovC/58uGztjbJBrGMFooF+m7aeCmS2di9I2AXC3+ZdPsUyUlI
/ZMqC05x53NHN3omHfgA+UOIWlHxI7EZdAaPisgdkEq9oAeQQgoxkx/LCDCQMg2pnn8GTx1TvFhm
mciuOnqMCM4WDoku96EXcMecQe3jLjTAyTngAGM1VFl3VdV9ZGxrMIyxNdR60wWdObNCuUMInGgN
uGD4QtorRmGLKnZR1zHffnpkK6F8bTWhck5gijnoFDasJCMHPwmU/lDY3dfJQV+R/EmAdzPO4c3e
Gp04sy4iVjN3KEuJZFqbVF4ZIxkcv42qNuDXuILauAe5mQp5Dh6vj+CMZU2pvwDWgv9LQlsQ9h4g
L/js1IvnrWXnr5l9ia4pGP6bSmO4hEI5T4AdRR1Km1CNNdjJ3+/9QPYyi2ulBqqRVWUphjAOu/VK
NNEqB2NRgYfJWKvQe92MWwibEz5BtllOBP8+Xd2ZkdPriDItvXld1NXz+e/PVkyb89E30cuSJFhp
xKcGtj+1ZE7JQUzp/CmUfvfjwC3qn7MC9z68eM0qXXUHHrwU2CVRpR0h2hEFu7WfyLYAeeCwbnNa
Jzt4X3BF9kxNSwqWbsWCpEWlLX2JXG5wFLrg3pLEMiNedr1afI9FYWAq6eNnO3zjQKg2WXQmkEv+
VIMVqg9FmVaTiJnIEKhObwHXGrAZNie2rTfsEGW5TuYqkhxXleBCn5BYR3qJu74Qq7fQA3KY09Df
xDMQT6e1vuhfL038klOrnr1m1jJGQmbKJqPdCuT/ds9C1ugHqai+bm+qgWgoboXMWYUz+DUlD/Pw
SNdyj/oPrdfpuV3DXLN/nH0yeiMdlO9tIJogPvMLPOYonfCuIakHTjdzVmqisx4Dxkf6VpOxfIYD
j5tSZYYfmVbDGQviei77he7bMFrMuREH8UwKxBuPZao7+NNeS+Vk1H5GKbKQUTWq0k5ZcwIqV/kj
rpsVqomuiT33vUoj+d12DWub0JvhGK0RnfrjVjNDC3736jHfMmkNY8G8cXnZ44Ad/Rc5DjPDEtdo
TFcxNWJgaOlle7aIwzUft5Ln0RsTtcM/8C59jpLgdV075/b/NU2zjH/AUONl6Emtu0HWoxvdX+DU
w0O0lArzdCfllsn2TgpLFSQmeRQFvrUcNj29DqW/DtRVwgIVl5c2n9jRgmRWnwthr60IBZ0AxXHr
Pxpe4BT/OQvWXO8J+lMy/QSc/4qNd1yaQzV3TpvuTQuFAhpct8dYMXHlis7i9TRCsEy4yPEpul+l
GXo3NyyoUqcq9s2hNl6THs4tFmfpzHHEK/vuxtHDNNvbqDBlcixcqaTxYxmKdwWBWqXO6WgPU2J0
RfiXh3iltZ2rZdKQpKAmURvQEYeiwvlMvh2pik1d9OAqBQ6OsQQ0p2pJuvgqM8H/W5Kb0nKtibd1
nO5SxVlpbr0uS1Jz5jj4+RNW7A9wWvZiLUAI3cnbVefMLSYcK3keIaBUZ5Vo2izIfYBR7au9ki/q
eCKP9jSrHLCsItI2vpGyED1g8NP2qV0VYpWZCTGm4Kpn9znVYyaQ0V0atL81lZf7nvAaxLu3BoY8
QM/LYJrcl2kr/XwYuSAOhzjYpceBGIzhEUIzGthRCAZbeosc+SEjVBLMJRQ5n5GZQwLSxafyPtFs
hwdEvwiU82DdFDTYHZ88IadtgEnoldg0vsNAsDQyglE/echmzak/NiB9eqb0DpDeyiNwO+sSmOUN
ucA6pcBIpMm0sqtYaSHqKaAa0paY0JxmR7lQyQ0zcRI4q70mhCEkxhHia2/Ba+lhRu5eoXuaaNSf
Qn0X31KJrSLhS44HJzOTS5qmZ9DnF6NG7T8qL6ODb31yeZqP6PlLb2mtMnUMCiNrvZq22W3d6x61
6giJZGVIWmzDgThbudftuUsdM0lgt+a6+3LFka6ICzH43wDO4V7kA23zAEVKh+//YQxGS14TPd+9
N5FeSwc6EwqmMVyPz4pIGYBy9MdgtL7Y/BQe6l2AwWCEgVUD9A7/jg1F8OrbKa7tA9pkJF+4CwDL
Jn6+LwyaBsPXQqRGAopxbk5FD7ysf3tChV4HPIpLuce4GwGBzGiL9F7etBR6leT1BLeQGZuzy2so
E6u0/PgYxW2mTn79RTYAPYjRG35p7wZMSzsLWCHUr0FCYeM9ORzZEJLaCCaYfBMbnyx0iYQefDsu
Orr5cBK0MflqNlsPC4IXNRoXfeJzsc7xGRcW1dt1GdmaFVDPzER8gvYOEygUTjXI29762rkkA4or
LNiLM/Gjm4l0cswqpciAGowqkOFKw1ASS8OucAYCYC8fiIZM5HeuSDkh6bQtJ8e61fUhpWO5kat0
4b9u5VhH6mT647TkyPJgTBTkAKqqsa2OUkO4pIhbgfXAol40Aq3djBMc6Zlm7rZaOWN4Xvb1GYTt
8Tsbmqj3vxwvLJNlEMMKVoW24y12KmcO5FmqXm+ovYxJ0hnceDnIUyBGNqYxFsTosybVwVXgirYy
fiHXpmljYB4JcCPCWZW0FSZbDY4FQTVhj43AKreBth50aX44nOUeoOoowmkGKnetzBU+8hMk4a1k
82gtivbpflzNMRWgIVscQ6rlMc09uBNiOYpsOJlb8q9xpgLsFflyBWUMI1cpEEYH/RKodIgy/AAP
6ci6JdDiJBWqyXY7mFaYJlYMcIvHJhpV9h56uo9HAXimTd90P9R5P+hU67QokbiQ3FejMUWRpktQ
Ne8nspAhfKBhh9GTgPHkBydUaQzMP38+SGQiE2oUOJ0Q3qQQ190+626NC7y8FP0vZNAtY3v5335j
PNhECJcTqAPIJ3+a+rMv7iXNkiZwIkaXQCEba2jU5K+BlR3Pd506/BMntQdiJXCMGbGHKpGKBJRQ
p5tFwSRT+T5u7NXHTxwzIfoQOSJRuOdtis+tJHmr1hFfy00AhlzQ9/7w4hzI9iDSSK5RXx/HWKvI
sZsuS+mnbWxkD3JnhSjN99qXoqz8jZoqp1wfuehF4Iv41LV5ll65ByJHTpN3QNh1OydTaTMeHUYz
ObuLDPfvb+Q6+dfIzLvzBgPiaypMIjSbmdQe1NSDHI+T1pWGGuokhXViwCBligCgnImaifGXGL95
D6Bumk7qclMFM0WtLxmjwH7yfBIiplh1U4dYCFroeSs+uivTlOwwf1ooSW/BzzpOhK1UafJuiQHC
yv4OgQO52rzFYhIQO0uHpLWTCxifXnPAkLlWyvxRnVFlMAHweag/grwl8jADBKXq/LFt/RtVfK/M
imjPhcuJ4FDA5o7l+mOiWazhFoa2AzcOn/TD69EBXVaNUn7C1H3nW5wLhq7/1ss3RC22na0dfeAb
PEDvaya7ij/76Duy1rCIBf+ZJ1HTt6k7DpHtZT1xxy/B38lDoWDgy0Rt6LiOv+UbtoAwPOm0y/KF
7a/uaHSvyoGeRTQ2Cz2CQN/LuFEWPppEoBZ0+3qbsoXVpFScBkOPXzIwssDwxGMD5b6SRSRoAool
smfA7Jxp3KEwuzKw55Q5jC0i+/l8urrr8NrMS19jsozNcoVxo7nCQE5gTfNIzJDnZeAwPN5xIeni
/qGVoJDOBb6+luS7o4xcSCW8ymRu8CIuYP2RmLi7Fodc4ZQPkQxR6HSIKhFOjzEU+bqNShqoZHjy
DIJPpIH4AZsfQgDADAQi9+cbHo/pa58P845EwpMIPWCOii9xK9uBBI7xXF5/aEPkeoIkMHTxOcd9
qHZhWpXFIMM6EWPeauT8JO6/rYbdkUbpauLwANM47L/Bn47IqJn/mu5HK7kTXc3pr/r75neGUuVU
zyxlqOIQUSVHT9YrRj+3o3AEvgzdqKmUF+X1OkITArQL2bbZ32VT9aSBAjJRuU/70kB0O+OLT80k
ski99L+aSKjK+OIqfzxxxWRgYtdxCOZgaee02T1K5jmLLsSQ6wZvbnMasXt9W0hFcjg8Yq0JX2zp
XffAZSQAk31iLUEM952a9W5LFweFDowz+SWz9y0ScmC5x/wUQ7Vr8i3icaXxEiXyS7TgMRAJGpCJ
WeRZbXSUztMFJ6A1d0TwKTrMCgvkqjj34LJZgVtqJzYP06z1uDmiO4kI7l9jccp7Hasqc3jOCiAD
vKVyR1DueaUEnVVzipIHzPexjiEiBKllKU1W7SUZwwDtJT0hABLDavoyD+t7YBT3FtFBElrdFimZ
8yK3IXphDC0nTPlzj2QrJh5h6dYmhwmB9BTQZ6muErZL9sdpQenSKwhgAwsshTVF5VrKxYXrlFvv
DC8GmSOdw+cymLdZBAJ3EMjG794GBgdVfW4T5CDlEytyb1bl+7sYtHyQeRQKsot8MUM2NXvaTOWx
ujAu4790l6GG9nQHrfG9B9UtugHyf4zUWJ7Iv+7V51UGpIMdVrW8ssocgukGR+R9zBvRecH/nxuh
dN1RXZcSxHdA/MdjMRvHSTW0vU3cwyVQ55xK+lEvgb37/B0HOyljv5oTy4CikTLRBOqfG+Z4zcGs
3cmPBhNJtLt6xabi9hITDzIZlaBKxjL57U7ss44SD/Imo2VUZGDuvMcu/AjI+vlgUeEY8zsqHl4h
LXw4tj1J+gceTxOAPEFOS2Eubd61JHiZLHPD5tcEeUxq2wXDfxj0Cn0Vld+tS3wO+Eg4/N1FvBSM
fkZdpPcddjwSP9RJeo7U4cIN+3Kq60a4zybyltqnm04/QY/McS9BNuDJxh4oZGI01JUg1EbbBQI0
2rF07eoCIuxGnePta7yWqp3O23hi0zUI2R2yozbzUTpAEN2mwVnsxLUWQsE81qcc1dW/lpNjVuZX
2hKcv9c+BVxGwLhVMZ7KkZ70DrETRnMS9hwix2K2Ef04qUr2IDxIqQu/xfDdnf/GbJIAXnFxwxyP
SNhja0O7dmJhLG91SxCHG5CNSS1ZaLJx2cfRz6lXTf/NiWSo192lO24v5ZPW/MGmtuiMFaGDGVaH
4Zvyzfd2agmqWSQd6jt6jUQQ3x99rUklmT7F7VTdH5zR8bHmYDVT3gz2rBRi6WEl2eBszZ2yYprJ
GKjuTQRaKdBKIRip+mkvZsuYbcBNFji6fTRzyZBKWSr1VWpS46BS96WOFoX6hDbJi64ymsatFyRw
JB/xRfUNrw4o6gPeJqAhafzEGRfw0aUBy2MYr5lMBH7ppueAYDDZ/MGAUJ4xtQX3438ELxt22IS1
axXvIEbJ626g81Rvo1IxWvdBJ0l0NUnydIi6USxk5B8IkRlKPhrKGApXB30Oi2p+6+On1Rub1NyA
rucDrReZAyLbbErICOJGZ6DE/hg/Myqo2+1WUk/kuQmP7+SK80nj7z0tIoJEwMOrPBvBjG8HeHFs
fvsVwjYZbwPdFFBEh4cWHcun9v1FJnUYcvjY4y+FHZJwIW8yLHwl4RB/KoVK3fPOaI/2LrDxPcH0
bC5f+mpgDFyhEMUzFAHRL/TuNKuwRXUWE/qqrkmWcCCAVrC/cw19Tf5F/HrcaBfYnc/8oGEz59fB
Z1IjKQHG2JjAsb6UKANIFTAQ7WcvIPgw4dP/J2DFgoJpUuB4DYOkV66eTJoXPgDYpYagmyt0NvrE
B0n5fVzrJvrpBYUIC5MwYoYSQnA6k+6r9Rop9B47jckHiS+neo3oTDVwh/D+ucESLsucc8lrNEt5
BcRIeDwJixYEprSs83d85zKRz953DQhlPIIXfDd1LeiPCk9YBVcItAYhczyCQk6lADXVLzgmCPO5
1SvbTRBad7eh7WRSk+xRltfgs2OiuKyaoH0K5BhW8jLWT6iJqNmNMFtTzFzWjVxys5bj7Of56oEW
VN0euscmtQEFPdNIcBbzUHf1qv5BobGamnZX4CV1ez95SGU2vc7udMsAuxpRfGlPUG6al4o6VX34
B6eLg+Y04ojI+5L68a5LLYZ9epRi0Tz6zNcQgz6j/UGWpFUiGieNHjveAMo/9qYO5dwItC4WniPy
eMzVnZPl+zS8D7UoVqaQm7kV/1pIbnookHA7vH8oCS60V7miWbQOROE7lsCpNfmQjbU3QXHhJeOn
r6xSISYO6WeIb22/Nl7JumL8dmiAKYblnbCgN2q8PWPkiAFLL1FVys6d5BNS+t9S3K/aOL/xzxqY
QLOIsFEjqJn8Nk1yi08fAAAlK+jrOFi2ABikioHUKEpJIbhNSY+38+2pGuar7Ob/U88/+0B1xJUB
kDDSTEU4ynosv24VAW7Tp3bs/4pXULVbKy9hh65iC2yh4ntWZLvcViNJWnPI/57llEzmcgVp3R9j
aPQxMgHK4EE8+PNmOGnKAs+hSKCIygv4c28lDefQey0R1oTRDiyTsf7dtPbbnwI6qnURagdeFmZM
H43ScycMPH8oOoiiZ1NgDNFR7/u3Aa+qZem7UL+GqiXnmGetF2xe8ucWLv9ZyQl1dxaZXbf/SB+6
zgltSkObhq2CyAfh1kS3KdNr7dZdDIKaX+biGVeNHhS/3VwtQs6o4Pvw4/CZto2b4jHE9kD4+iHT
rV4dnhmXsdoa/xGp+pZbj7nRnwYGkNOdCjAXQGMubE0O8Nl6OUkMs0as/mfAruClYBA9rQs5CMeI
taP5ovVQr9Hk35swxlOgX8xb9nkQb0UV4OuaCymFsXcgX8+IaPmifGJ1Zmhy2ThCrJpyftnVfnnq
dL8eDHEPvNk3z6QwKA5VtQy7qiLk9St4MOQ4SST/KrwUs/uiZ/l0KC4l3eeJYysG1qoekVqT/n9C
hb58KARRZHRGyXXfJIt9NfGdOGFydlR2pkZN1LwvxKkvg8pyIoWZbHA6LGyPcBGex4KQ8pYdx/uK
77yF5nsTAqid/fQRqMnzhrrRxxvsUplUsAkyTdJDDaApeZ3SVL7SboozDZ8mgkaP93GTGa+Qbps8
+JGw8kON0IKy6xq0AkLhCAN6PlN32ut99zb/+7bfjQwRmJCnCROUNONAv+KiCGxyTDeWDk0bUury
Nxqy4KdO7EGlsuZSaA37aiTH/+uWZPDY9S7fmoVB0codc4kH7mNjx0NA0KD4PYbckeNU5s1fb+ko
In3Dm5LcNm6sbUoZjgiyS4MAVJUPyHtn7fERrjbHGgdMqLC06Ov1qicL4VciWXUI85BrBsTma4X7
YC6kwftifwIjC1cyY2Jj6jqaV3Md8tJo71lgUdd11cCGyT8X0qeMybnU1WFvtV6/ffIH9H9sPqTR
5IErhoDZRdgUG8JbgAH/uwV/jhNWzzGmvfep1Lt5PyDnEMndcSd89kQjEFoSo0KByyg6yIWOrVmH
ksCx13ctmHul0zlEhL59j8RyvGkh8AI72I90yi3ypL6qYkEtjWF+5fjhLtRrBn4lQa6u/osLf8my
0olMNayOG80GDma5jBbMXg5MFVOq/NhUou6yUT/EWIc7gOhLsVp9+el1UrjSv7IUeW5rwODw1mGx
Pj/JsX2Cf+IhA5FvUKCtyvbkHzDpJNfxu6wOjW4EC/2MHW0rIUazPGaDl5KD9qGVt79F36BI0fYp
LhuF43OyzqeG/OHb1VH4ouJ3sgaEdSoDnz+avJdhqRJ5JmBaK31eyIWYsVgJfJCoWu/ZIl8h8Zk2
19EvOMA1MqLXWrixt7lFwNElnzrq3RUlIYq5sIPZmSyUbCL/tbpULTljZOauC48jm4ek3NyVR+QT
xKUssTtiM+eIIwpCyQFFmGAweq7lGyzVhB63OJ/8tq4/ZKpsg6DWCr7EHCgMx+w2cB9uHiRSUjcG
EFbpgJ95fiflfDDGXu2ZJn+VaSf7iBCiv2BFRokVne8/jR2mkHe4iYwjlRhUKB6wz3IKYAyqsj4l
da57diU0PolOeamUuboQ/tKguOiI2+JZXs/60a7YtoLn3EVKBwfTSSH/WCGgw9uiDm31uJRGiA2S
asykU0jVrVRKwu0//KEKm+KCXweLDoVl75dJy3fFR641Xbzv2+wJquaV8Hqq6cm6ZYiLuXFRFBr5
2pEGJ0u/lgcerS/XZCiZ4Sn3Sbv86y2pTDWj0y8an9tR1XzlwRBDda1YvbrG7xc0uqfQzLJyOA/u
OlKvqqs0fcbjeXgPQWHqPw200/cxSUUqZUlw7sTVfPmKNWrp/oR3f1krQ4CQIakC38sbypqzoLnR
+olX52CKjozq2d8lQhsPUd1nn256weR72XJYyiqd0YKp3w+CXDIGtwClLYyafl/aHczvbMoJ++E3
HfkNqdLcOV/yo25EXKgOQac5L4Jj3SW+FISOooF9RmQsaWrxyCoKcLsFFTfJXsF2UWsd27/g1mv4
RzU2RwhpX5PB+ET8LsO/HXxz/y6CNgrgRrMstOP+OVXqdydSZ4YpM/SZsJWo1VzPsdQ8K4xlD9ov
QP9a7I7CE8KjxEHvxklwDtFyToqfFMYSL4cTxmAPl8FgBRlH8vP+PZYp44g7UtfCk0Buy9+FoLRA
UnXa9aF3EeNlX0+ClHIBre3e7vrmRBY1NO/K802TfIqwWZ6andjWEjhnsgP0g+BmLxMn/yZZCqg6
Mah250WZrI72NlQopamIUxuPCgemGRJRRdbR8sq5Vr0UJNIDbVlIqL22TlWWMeh3/uFaKyvYv1oe
ryHC1HEm2DDLjKiknwKaAo9nOzOeZYAZHdrzXboaCbrKStFj2aNtw+96DFgE+KSKRxNI2WuQ2oai
QZlDQvWPRHAIzrOW5cXLgB039j2KlHOrbX99/9qv53M1nkZIQ+mUs3PfwqwKM47xRHcyGYwAIM/F
rKuFXKBQO3Bf6zbpJshC8JkQyxjaReYXGCm7UsHRHpzbH/HUpF4BSIUmwvRW7C7Sj8keTv3tQLO1
h1lkTW7K1/rfNWqMiVgVnjv8bqgKDcQEps4KVk+pZdRi0TsVgVUiiIlAP1QwQUDzrMmhlnJPQgfL
ul8cjCUJkY9w4Jiryk9chvAib5gFiayXalwKW0Ym6V86hQcao73ANIJsHQ5xw31dna35rPCMcQ+t
UCjLqYsU/Kdql9h4cZTHOd0t2lwq0ULXRE8H/M1S4oizJqijrlKVNGM6H564XC5xztz6zd92FQdX
VYByCGXevN7VrLNryeFF/NW+KkFPow7OLpL1Hhx8+fBD6+cGH215ri1y6aH4zJJa6M+RqCS9QVek
A+Sk7Go8lGAqsKX09yz7ey3vF1f8RWpFOtuL4Yos4x68oZvQughJX6Vbt/Q2p9ZCE408tPl4NEyY
H1f50Bjcdzr1Aonc2HHKu4q4BJUOmK2+OvzavvElDm4QTdisWViVYenGot6rXVlFDyPZuEwRRbJT
YwsIMA3YHiYwaCiIE679gSuOn2jwLTnZ0dj1mW7BSbKm9VPSQSZRim/wwo9a6D063hiPfqGm+Cm6
+r9eu+uFytGW/+diRDcAKHWwsfaMoPtDso9Ps0Fd6+Z6TCkzuyViXXU7NhzuG94UNmMtf1oT79ad
UakAjVIa1/u2jUBGWjxxJz4RgJ4/XJZJaI7R8lfT4tEcbhe1SBaFjPys5vbY8JjO1NcKC7Ex29vg
XLuerbyVd8IllWZ8wND3CVDIPhQzDf0MR5W5BVULhjylR+Udyut0aX0cndnN7UpniQRNqDLjoJEp
nteSwoOguFbyrCdrC/sbqXwuMkUTcS44vsA2q2LS0RnUU3uZMLaAIW5bsG/Blw7+v3hKP2daVrm4
rF2Ri7/XxfcSuNSd3Jx+fs6Lu2LpubUNXS+Gps7fOOdoAQeyVM0m3bRoUb0J3XfnoKRmIutadQnS
Z6s0o4plFbAXYlWxeQmJb4R9jYbAzs3lWkLYd1Oi1FPG5qglRTQX7t7NSqoxaWAWr/O6QVg+Jt+t
wrZpsvvKNf5kXnGy3fO/1jhvzvhcFl2BKBHDpFFDpjQJeZkzkll/qumnBnexR13fDyJLXQZWiAGX
PgXLymzXHgOCtu2jf5fDedUGqznDm56mm1easrWYY6bSPbI2OoctVbDpuvSccn5AjQdXCynq2Y6p
zkom86vC897bA4+5Eq9S7RM1JbP61lmQNzhRBVSQOgffIvEHCPi/fU0GddyWNyJjGJU5zhcFXZuX
llBIWRNJhiHYu2zktr73Gg2oFG9aydA7cZLp6trptVqYvYPpA0vRRh1gcP1JfHo9+l3j7J46Dg4V
i8vrFcY9ZIySzBiGwI8qYaRZTRFl4pUVUVF/8Hv+IBoOW18jfjTrYwKXj3O2jSnNGdhibikywLap
rDmC+fBqJEhs4EgEzy/xo6QtfjgXGtCbIlKeAvDIF6TmRf7qNpvMG4xH6ylxz+XTzh1YThCnP8rY
nZcelPlh9SN05XudChw6SHzVq8rLMK7/HvdVcVe8BsNXfdi7SG8Rj/LSIOA9LztpjU0oWvzBXUak
yFlbXOtW7jGqW9PMxYnZGVWEbWaRpqnTOnp9465udri0BvQXWPnn7pmI/26AL57yzGd8qS3KJt9m
iheBwpbMI/wgzJg4Y44y+GjVDTGVsC+rKv+aGBl046gczmC72GU5KYCKUMaSJmNyNz/ujPf2/Y0C
cmO2pr45OSdjDUDnpI9jTVQjslkLoP3Hh6ihgHNZtSq9MXGz4+IOxsT8ywiywN/TcmrDK3djbARR
XCYchEoqUVSx9bELUS/oreDoBDKHkG7zrTT0fFBKnDsqSbjFGDixbv9aTkZRj5qsuzM8CS4/Hccr
YnBz5z7V+TJkw3v0j3tKrdRiJ22IsLon3+0mxNIRX3s6ztbsto3AH0PupUusHPYNwXQ4uejVEaEX
vhYVmePY6isvHKICR5plaejBgCT9pv711G8cvUkaJW6u+RTShUc7hdQQN5n4+e3Gsick14fdkEtC
vdCuIdvZdooUdgnzbasAJOmSERMXG3lETNDytLmQnJ4yUOuaVldtWwzgSEkldhUospY6QaxHrCCV
ydFAIm2hSF5mnttw9UjMWQeIHPoymg8M49YBOBcys4QpAIcDAsnHy6SnbUF5K9ZNadJiBz9dklYE
yCwQgIe7BC80lA1kl9KXcd1QxmU5yVtXcJ1G8jj2/9RZlCEdGCkZRxen7zwzO13LTyfqi9/QWcmC
otXOedz0v58A9rudQyn427yAQu/hgAXVy9IDWRegsePijRUKo5weJiXNuL3J+YUj0Yj8cp2inW5l
n/aARJwPuuTVDvnAbNfp/RaA+czfVshnuPR3deBy02yJJ9zHk0o+t6VPWiLNDEUNRIYEDqmQCKdV
k+f6Ysl33gYJt6Ri4IyX1Bg695B5/DfwWAdAhr9HQmpi9CETzK2Lbq8gR5+cQS5oFywA6vNrSXTc
6DLwy64wLcFdce2FlOYhNf7m+17P25Gj5ntlIwPgmxomyFB9DAxoQuK2gcf9Tg2lCiLUwZZ13mCj
KgO/sDA2ggqZzaKGAOHPBN8z1orC63l9nWcPoV3oVFO7z/8tKKYAcI675To1UGVk5Y+K2Y9fQARG
2TlC2SdLrY6LtHuSnWWz4dLk2MYoDAPqIJUu3CD81Ty1pkFDfg1/AJMpRkWuzOFPDXqoI3FXyIoO
z8q3IoA41uxPydwtolPvxYlwSA5MCRmGyDvHcWBHAYNe3M83Tm3UMn4mGQZ7UqzBB8INMDc6/7/e
kxrD6L4Qoor9FeNJju9cnlAIW1E/EQ4aTfnL1j6cN1i27+ikNXZ2o5/6mleyBJPCIGf06EeuHqN2
E/i4vHaP8SROaE4tP7IaMOPg2nU8/vapDsr5nvcnUi6NAy/F2YaeByczfXCFgY+C1rgfVeT6qrUr
b7+Li1CLV5oNJQC3zmZtydc27e1xJb3RDdwyIgDEMQ2+7um4HZtHshLDzdHUNxDuhY0p8V05AkeA
neR45xZCrjTR82bd0S8VEoUqOsJoEAdmWhgqzevJ/CLEaoZMy6xtkYfLEFdddnn6lMODzwpaU32V
DFt7TT7UaXg+VVJ0wJ/aSpLLffFAT/jjxh0a4PcjjucK8mglcgIWYACTn0A4uxiKUVf0BPsO5ONj
hqrR41gePmu0Lr00hzjnbob4F1QLlun4cqo5todwizosHiG42zf90x9fP6EW8nnM7yv8SfSBcgH6
yv9fx4ApcxTcvMpbA+TO6GPNlsbFmLQL3v/hQKItByLl5iQ9HUxljiphxSuOUUAApCbp2q3NFMwu
u3IbT1Bexl/DO3SiccD6fKV77yJaOThYjkk+5KxKrnCycWfji2zv6ZtfmlCSA3si0VKX/aKc6WfK
sDz6l/U+2qXfBqPR639zbulow08zgl30GaTKBxYx0cwXYASzQWNhB/Pq21hPU9l6JtxGEkek1tia
kyK0E2Owr259pxj14ce35a6KuaTQy60WoI+SkxNqXT6DSScDq8a8UUdoswpLEreKyYEYYPvHT2vt
H+Hu47lItJOLIjHQFqfby6ES5XYT1HxYF/8Y1o5CdNNCnV+zg42oN4wbktIS7UBgqsTeFy5h3FkF
qWMBthFmUKRTPS3HoL4kdE+UYpD799Mu17TLMarD9sgexFl9ADkHJzNQGuH9l47CrUuw1Br2HkqJ
uwvEnUnpn9qcOz0n+5CRcmMGGdTQfIcvzX6gbwCTVAvCrKwvs8YKffThZzMnahp4dId6amGcQiZ9
Uvf5P1aIv63jSHXSfBJWMEbKJZ3fR8nPwNnXegHsuLrwA8n9voyLJ53sV32OGtu5DIzfoWsQyW4h
lUvxldRT/wjscNMT3RMxQdwp3jDxpRIUZ9lhCxHZeJwqPl9TTrdfCx+kYKRjSLKBBi+Xy5dSFo9I
y2itDbJYLUflPE4zLchuJXFqXbDFANZPyb7dTfZWg6oZNhJJYZ5d4KaQbruUf82If7pShImz7C3d
jPshyXcfEo89NMf4YgVaj1vRISmEJz/80Y64g3GNd/horvcO09BjX4vBDse9DBE1q9eH04vAgtuM
jn4/X6M1oPXj9Z3J3e7tvSorDHLMwClexpeHJGPtVEtX6uMSi1ESMJHWPJ17+hBvocQAk+x/kYo9
wM+zUHxAyVe5RgQUj/Y349n+bJXQ/uqRE9dpRDYMcfpH4IQrgMvQ4tdi7r3zrVLnj17y4oizNJir
Q5Tv/ZBQEpY8DW3CfMopC0asr9Tfyl4gb7x2sZZVjGrwv2ZzNOS3WTK4R3Wwmi8/CFZiFhH5kpDW
sOug3hsMFjGE3ynVLb1hUjWg+BlkKRIArnbqpyxEtr4JKh15Wy94rrOIUaxklnTrcL9mRfDbwvy7
c/L8q4NWzzaXPhc8AtgTZYFq3j5eqFsYMX1s8IJyiQetbR91J+cHLlqDeXKTh15NgX6/xhuGb4ft
kMGtvJ90JFj7QkNyMxPYhRb+cCSr4imKdcquCUXpGjbYWr05pK/LTyaBfrawJenrW290mlypzK3i
zuMVLu+dlBcJwl1EWG5YwAcWmlawJhwhTf9uD1AOmgewtIcKMPEy4D/ThIF+N/Kq4nuMW3Y5tt4w
lQIDOz7LeBOpOxSLheYI+SBKzC3pl9OD+VDWd3vNIlWprVBEqMPqqtoLXdqfbMZbMmpuidoRmlmC
z4Yj4ab8plWLei11um3nWM6sCa+a5DpBMhNY3gBvUOAafHu2NZt/HyP4TunQ3JtaQDu2B99/QYbG
iFUZLjQsZf/+U6ZqjcQda/cw3OgK6bWQyr2sKYttVr8UMGCbqjTAvg35/K1gzOVzsHy5ICWgSPiS
EG7PShr9JU3O54uS0g50JujHuAzT/5ON7CG2ZrVZ+16ePOE+YW2vCqhurD/bIoLxdB65rP7GsExy
2Mm262YUXRoQuzYu8H7XyoTJQJa4RQ97OHev1KLc/ZZziwWwlFVdtDRC1Ob3UDqqFE1ki2BhoAu4
Kyw2Bf0a83VRSv85vUfVm9e7y8EZWfFJb615Njz3WetfOkjsRdJu4KqDiWadcuG2PvME1z11HHNd
MJxLaxqG0FurAQTqqY7CSlhs4CzlkQ+Cc3ca0q72hTpGnONkT5Lv2zTquEcdyrfnmQi5n1mFpGqW
phyucWm+heiP+yHelVGe9RVZJzS4igIAmrlsLZDXp8oM1f4IOxs3015saCfqEfqZsPFIKj9eFtoI
Il/0iFY5uyIEy6I3AwzCG5ODP7TFp4Xjhy4KpG72VJIKKq3PW9bToUh+u31hJpYafj92o3gpHyUd
r3zx+ATXss/0y0VB75/R4qPtdtKinfjA+Zy4EdDxXtZbM7d9n3DpJalsT32P0tquV5vVBWRBUZsO
v1d8ICIdR2f6cOEjNAIoLM8YlZyjvPIqTafYUJ+PiTnFzXn8seL+fWEV+UkESW3rBhZywEtFidCi
ft7Q7OavBPPNMmTGA281bdEMp2FEBTYg+tGI2OVasm4zhM1Ujq1sg41G/g+bGQ+uE8ZtKdfCuSBe
amAYTLZHJdb2Y8Z+ClR7bCVSqJ+ge7OIoD9LSmxJdTNI3yVAvPE+ZN3cErA+pN9nBj7rfp3F+Nlb
76dffhvAmPVKzBqGk80TgplVJoEPz9pfcdv+N/eS5xdjSp4ihfm3GVkEAe99xuxDxwCkmNRhCQTe
wjsmX2Rkm3BYKOaDJr1zvoZXv4M18R5Z2mbhaiRDw5JMOPKxmSpqLtDeJO4n13Cw/OdI3RYrXq6P
yDWb4i4o0JoEpmC+a7Mkf9X3hwmyyalYf+B1P8vze7QaGBUAGkwx8512gvMu3Goo9HTjZmZ7J3As
LDy1OWagWk5ue+IsdciQQlZCdCWyHeCaLkmhHae/GTYwAzH/EU69redF/NkNXuAyqt+qEJMF3+yU
WFmU+mLSg5ugj9CLGVo3q4r7koCNAst+X9W7MD9lqvwarU7kPmFfmpzd2z8zrh1MzUg4paYpUp5g
Ot/8+PkuEBeg2c0INEDeImZGAWioEBikEcNYUvQbgbTyWG9w6RcYSiFCAEHkWBoBipzRfx6aEOmS
dvSPjThdCM/4kH1BTA590n0yRTDbqWdbmneJo4Gv4VWLMfgy95b/lXSf6vUh1uQlRn0cTSUXtqbc
D9Ky0ttaLUR7teSFV+yJRG7CWJpEY8/in3OcWev9e0dQEZozviUSv7bsjDjWREQebWIklTlG0bRw
uXPbO437D0BdmNLDnM9PGpBxSu7vwJ0JXkhmQe/cAhRwt7dFWG0Vy9c1fj+DFpn10c788zkP/xc/
UiFtTGFa6zCzDHp/ZPnyZ/MJPq8FWalSjt7+K9o0erQbKJ1QfF3xRK/5lMXwq5LrtCBcWPHOeqBV
Qi0otwcmARDFyeMi3JFWHKosblMt2pnPThnoyiDfUkaAWKdUem7NwBepIAY+3Y0WKBdQOpPArVE4
vHJ+A18VP82v7gh0WQCTOx+bQ1NPbYpqUpwfqp5pTShI5LZdOt5BOFrbrieGuUsthklLUKlqcLS8
C80+6f/38T2DgnKFcUU4l/zp63B2LJGVUZkRRDpYFZenc/ZNWwC0GP4eMD2qw9MRieu6mlBlozYH
FP7tUTc1dGBEAzh9Ja9i12sD8K07497j+Zyxv+QklvUfRFjZY+BbHx80yzxa/1Bcf+TQiCtnykfR
/saYGXzz8+Od8KNb22BUU1UjPYAhSPVV0a2uWtqWrOBQCm3vdlgHUdbxcSoerfWJw9vCiS+DlbXm
QpMFTO+AGTNZTiI624HvZPxuhEwXQlIVUjqASFMUReOM1msLx2veVa2I0iVNpMwE/Acc/Uu3WE3e
IkAyW7DMkq39YWBSih7AsLnqyD1j7E3UOzgVtY5CmNCCIK77njp3XNFn/TC4OMcA6DqHxtnf1p+d
vfTUZ+IwQpId6QwhDf7Pj/QKpfUs+V4QlI6HQnc/A8cTfoZsCvky0ikb3nCtvvUsd4OtSMRCYuse
TKWUnM1p7SuSm7GhFdknyRT+2rdOwHH5wFDIyNXQPUMB4lSaD7/Y9KxHdZdWzgfh7ZSUZ6qa+qFd
vlBU7mjojSzUreoImqmq76kaVyGYPNCftoxDxY0e2BCL1JQpmPec/x1L4DTJbIWVqVD4ChzLmL4Y
CG6Sh/2ZlgFUAEpcNsvX3UfO5zfhb5P5sLzWfwnqUkYoBhGRlfaaYZbsXVWOTTXcgEeyepvCeLNT
vB1oDvYbnmXzBQx1Xr4W4kSwf8sMLVRwDSWUPDfbY4zEH5AeP6BWXcd5jExu7veB6uc5OLzwymJa
1/hPeEIATxawIyw+Ryfvk03FG0HiEhKlnUuCtGfpWzluubVNstWLBhPwKRV74KaqTpavcpQVmRH8
sLCAqcYtIGUEU4bnIPcIEx95Oj9lrsnHzLzluSJLvv5SNBEecS65pO0038HxEsObPYwZjHYEdYNx
Wq6uzPlDs7YARwgRziOQpGPMQa7NbN//n77CWTITNKhScLVMQtHZBmwiogoosF6RuDbDUmBv9Iht
dqON5m1P4kqTlWZL+br/oI51PNHH7/1G6jQtzrepOTXnIqIdysQyADtHr2dFRioyWpTZ5JBVPpUP
EQP3oq8wCp+blPm5jUZZF8KdjyY02cG5u/3VPHcAJ3/OdvcXec08CGdOa5GFyYHOtDNbqFqo/xyE
QjpyCv2G9QvKQ4vDR1zMOrECdJ6Zh+LprPujVnvm+LGKVl+EDuVu1LTCT1o4J4dDEEOxL32jcmU/
amVcEiL9Xg8WfSiEYnERlzbQ+eeEIZeFU3zxMqkfImOq3OZiQJzAipqOLGuPjVQvx9CRwO7k4uwf
N9tYyk1BMRIZunFai7MHfCEYyzMFsnw0ADXPQx0OaECDhei3nukLFby1AozpgiaO+hyknzn7Pz8c
0uzpmp8Cm7r3/NQ08vJ69eOWdYzH2USFIXfqkrG3QtPuLPmr8Lk4W+t/a9FzNSz1D7xMFZvFieym
9dSrLipStkUo+BJUKmlL054xmyQVQ3eZpmoSi2LpmnXIskFeoUK0nZmnjz6S07Hs7tPugKo659m/
EqF374C6K40U0JoEtE+AZuubMy4bsnhLYG0IQ0jsxWGralQonUbi2PrdzrgSlEd3NIAf2tghnDAt
c4Ml4X3HIo9ZVUYcsFw85wrtXQW6w4zf11h82/CSlSOuyErH/Jkomb/k7TDwC5RUBAu1Hcl9XsQi
w3V4USkKTsySPMsaXlA6Gy7WEuQPcMhHqG7Cvoc5xOAMwrbXirHa6raEsrfTnq4SAOEPzo6G8TI1
LAOkEDsjzU1Q7FlLszCAm0HcjItyibP8brkFIYpJsKGN0YCKav52VHKB7Pz6raCyZ9vSPgjSwhdj
2YOnMTfoqrq5Xvg4h7GeJpzpfAVebGX5Rpq1stN0bXxviZP3aEsGjG4EM2c6yP8fZ83OjuSpsIDN
0ZrRJ7VhqlTWMkb3+XuQhP1Xh+GyH9DXZxDRgGtkpQkQMqQNE226859uCFyEm4oS0IMiyfOwjTzm
HMH8Qu3RF048o7NMsDZXrMZKCYajHfAs3oFg4D6JvbBmzigzgMFYb+HLfC19Ep5hIxIk+UbZLlIV
RcWWlOzxivVaKp9wr4n4pTHqRV0+ji7W3OABylcKo46RMOakY9tON4QlUUgPQKXh64Ty8z6aQvr4
WVuiZ1u68Fc4JWsLhWF6J79FJwslrOFFsWkKuCyP2Mj8KB5GB8Sc0mv76WoM40m9OpwGBfjs9+mA
23SLSSyL12h0W0ZGE/qwVELfKNxjGeqMUZDdEfhWB9J1HQITHSW5Ygz25NKwXkQ9B/Pc790z1ihN
SC/fHMwgiz/p8/xixeWOYzsTgxV0Vx8rmmmKLFQ4WtMiAGszqgzrXTfQPlkeQpSxFgCYaixwa58C
ZUcur0ezkoFo7vWkwVv5M5aLknyw7CN420FQ0QjzF/3AuEwbZSDBdrW0qfuiWTBMOQlvpMVjmcrf
qRuICyzg9bGwN65CTGrOLHeGdeQJMwZHwdS+Z+KfS4Jb3Ahqwye0f9snIOpHvbGvLpLBrH920F0L
BlZJvAEF9VPg40rHpHoYKxhz2lekp3ZT6IHeQ6jMSZflvAfcb+cFrJ/ICiQKLviJ+SA5BKwoFlld
0OTLQ2qFwU8t/FCC3yvK7QBMwRi/cOYhTa3zp8QvNgL9Le0j9+cRm5KnBfBaaJTBDBdUF28zrgnw
uQSVV+RqLKUclYFFzcnWVzUd05tHofw2FMBNpGtHbxAvUUDjSSm5jTgD0JNuete/IIejX9bVetmh
J4i0HITpWigSmLf4+eZcfBdpWGcELXm6X0sl801om4cpTCa8i857DSZaBEMuEO2rzvIGcIey4NRl
IohfETxIb+RQY5SjDboIl5xo7QbDMQYvAa7fWzrIf06R4XNHMq8DQvPct/8E6izRXSVwwIAGWrg0
Zf2ELOSKYzzbL1OqB7t+mDmX4m7Vxj6JazjfhXGRK87/oZMDaUynUSwB8NWsWj9kShkQkvtSxSFc
UZ++w9iV1sUsr2BQfHhP8a9CpEL6g2xn6JaXmmDXdrG2465U74154+Wz74EiDI1zBYaQ8nc0TgtZ
fUnfahn4hSlhmARd5PPnOQierRHhr3kSLMClz7TcPS2K0Eh/uJU+TBuXFVbp860csevPPMC+bjqE
18T3Z6F1mqtYxbDMjcP+2aSsjmVSA4lWueHCnWKlc6a7+A/bvgAyDCGq0hq6ItUpe6jtUrxsTHsk
NbfXdfwx5pW7lAAiQVOnGjykDj+CLNmammO3kP+8ySdKKoAn1bQNCF39+JTNDF3bSanRa5hdCFKy
B5b7b3qmea9sqAI2MiZt6Fh5wOo84AptID+9oor6lIQ3Xu5hxT1pJUgHLuna/txvwEHMkrIMAseI
9skmeoK0rkzGvSapC2Y9t43ax5xnISlnVISwqmdVGemToFKVf8Pcj1hQbYuchcEqRVBzMuAJ3vjk
qDSQWqbGdUIqbc/JjBMyyBtTsERhNPG2uxk5lVeWuxxHsaLxXUY5O5MWKgQ/fbym9sLasC0HJSiN
RW2GLX+KZOC1kjJcDLBbzF2JD9hzW1pAXn55nRgvx9u4eT81gZs1bmLXWARZsXbbx/kakB/ijm6f
QB7sMDzYJcpnywAQEgOrHGqbkjYHQ2OS3Hh/mEeufkddGJ8iQmB2QAZjWKN+3NiKcYZbJWlFTKN/
bHYYxdqoZzRaVoSF1KbkFy4RxBBl+/rbURmeQT4ORZ9JbD6Fh6aFQn1I5vxFyGNsnCkiE43WU1cY
6tKBfMelfd3YRDA47GfAPMqCqOeQgeFlpg31sgRaOheT4RC0fGkOVFUw4JQtAA6II3pI+HwNkbdX
GzxytXnWV4KRZgSuUwrj8IV+O6MQrOiIcmDtnK4P47ko8ZLZai8FgROV+0+t7vwFTlLg8ZOoVqBt
kOdxs/mygdXVx7YgO+gHLhPRyPqbbDcQZFbBHg10KPm9oQMC1FXTUBKto4exqMu12UMREXx0PqOd
rIjbw8eLsQlWviVoDIXfnmOw4Ock6Wsl1hNMFvvVz3OhX/vK66CeWDWW/iRrIUhkWGaXU2rsKo84
UlOEazlIhN0lhKZK76jrtdDE0FXNpnV/kV/7MdEAK7WgVv8NuoaB6pHqOUQOEpOW7UVnFvMaii5v
zvogzx2f2ddfPATt6XdkRuChB1vyiTqh6/AbaXqx2QWPuypvXpwxcPV+LjZ8BtjJburNKUWrnk0T
RzNIKUpfp8gAB5EELAH+B/2QVgCZrTKhFmDjHticj1mjode0KPzG8wl/0dTJzHjqwmY+adoeYBgn
8dRsVsmA57e8iAUbdn+RWxtmmiJ5pqtsFxiMRF0K07ywkHu1rd0cSrH0xejGlRmESUTuG/J8QyeE
iui3IUV8xFMM7itdrtwYiEihbuYHGPYOA/X/TE1oI7CqCSETmZMGTLDXNOado1yGCArXWvxnLzfb
DUiAgVJWbzvnH9/+D6x1KQ3/rR1G2lfpSLoI9WMW80gXFSMzHQ0NWQDseGI9bDkyLGBshfhYeYqH
0bJga4ZujIBi8eVUEnyZw1ECf8rObN32CSouAQ+Hz85BT3QiNdCgYAOxjdIEagIR8vOTQsi+ZBuC
57Q8qjoFjpMn9XGi+KufGhll9Z9FOWA/HTcZY2PdoGI5bFTXEeEZFR5lXgWo+QI+odo7PfhOZLl3
wgnic/DRhF9qOscouK5uaJMWzMQBCOVeuXN1by9ptQglaewIT5jJtNiwY/1lQbRYNf35JCClQ/8B
3UKeYhJ5VH/ot4QC938oUMPgb243eYogLVkRdtfljkQl2zyzoTNP1Lr1XWT7zOuKWlGqyA8TCe68
l9JbOjPHTq3n3nQhIXkzGpGBBdr8SmQzJ+7QfslHdD6aXogC3ZpVRTQU2U0GUSNmjrZW9GA6PdQq
5ZfJo7Jxd3VfBwxJPKcH8gybWtjaXff2sGfDt8uexAprSYEmWWgwn+ZYqm5F50P86+bS0zIrHo2U
3TZffh+p8posYBIIoczBniC8WioCtiu28kXTeM10wzzjHhajHEAV649Ho1tncPXzucO/Phqqnb4V
1hIqwITivZPIgrhUXZ6bmWQ/xgfSlnFdJ+wtnM7CwL+3P2J18khfPTTGMmdwT9ZrfoK4LdFDbbIJ
/giw+NbzDCDE/dSy6qOjmFEsL9+ISVzf+6T/hn0R1b0+QImuMa8qvWVlc+D6APjzB334qRwf7KGb
Zxo2EFTuIOsyaqvqYCHjPbOH4oBIuJyw1y9MIQzKSdr90mlkDWfiFycTaf/rYejPDnw7KYpuWKtX
2Kp6LkFyC56NaUySXJ9cAILdkHXysz3UZ6O6Cg+7q/xT0NppPbioA1k1azBgsjFrm1vKIBTgUZaX
btykkqku8W44OxgB3WCAr/ZHlHchUT3R4ApWxL1nJZvpKkAamGqeRlbAUt6gdE7lBY9Q5Jwpjq7e
2u2BISyIrx0tdLhix0t7ZfKwgjS1RHASxTbdNIb+VckgRljD8R/ydcmsLyjbJMGmtEnf/rigqcOF
1cfnIE7XSQdJl+2GBLBiMb1HsoNH02w1twgaaygmwM2+cEOppEcABoeepDbn3yfSryHtgxtdlgjS
CiGpTtRX8J8PmWIyYQ1C3bFQL33m3527fIUFYkNahC8G5q/hln0US+fxo1824DIrAxx+pr07ih0b
WtffkdVjlaNEfPVhUtyewyIi69W5qhC2TeFihEUF0ySzP+fRNVsPc1tlKtlq06xEgV28UEObpsdg
FrAXRWUDoKVM2rBEZ7sLeDxgY6WrpMnIUec78GhtZJgnBWfwmrgVx1cw6cNd9izBzuXK5mg7rcQI
qc4Hh1CSfSKdCrggCYTbgJvYpcwQJhiv52WuMLo7xgao4WtZstiv5NPa5UiIcFu+XrjKhbBAMoBx
/vqKIINzpETMRRBUDadmWiCbkc4mplldi0nYyzkCwak/X9d5Ixc+Y2diRm5nHgbM3acZ4MRuph12
3h15vhrIbW7X/2I6gt8UzCAOv17Opq5T+YKqunb3scW2vKgiIsWodyCHhd/ricK0+2iuftgYBEWH
WwX1MB0kKrz2RfNxUeOywOgK/9d6g5OWHNtAdMbJkV9TkF33vPrszq6OoxXe8IdSZ1rqPpaet4ZD
CpBWQm/sKCeMAoB3kkjjc5ADg7cmOAqZQ70OnWIoRk6gF8OujNxPb143PREbjeJlWbvppwCGpXHU
QT6xfLe/YlKjxDEMeGFdtiEtI2AK72hHKm9mYHKcjbVQf41q+u0zOSn9nQnmu9i9JsYPW1fRJ3bm
uCjzhrnwfxiDLyVWZNSpM7am11RueAgKU2Vd5+Cdj9qGiCeN6WUX08dJSzvmQAZfIeNm2e9GYhR1
ggzCNQkIa+/x668/lZgpMcJdkKJ3j7JutEkYIMuH6O7LtcE3zhzzRL9CMPvLWjguwWBy62BevhP8
M0coYifhJcrjMuqgEorjcY0cEAhYEuAI4YiepOmWYE1otgM6McSnYJrGdwOpkTIWCmIfFKgMBAlO
6ob1kEIcNmYB3C1uXIBw2HSF689J60pkwE68HufOcfgZIulglI1ESuNz5z0pcUba7yN936R83bpn
0zlJDxz3g4RrPpLoXtkEj3lO7Ti8RlclA5eltBGA+zfRvQlonQCEZ/9J+1NDemNeW9aoqXtw96+M
3Gg7+ywJyaHu9jS+fQGN56DrQdi2S3zAk2WK+gpAAiBymt7RLnVquSgkxYsmVE4SerYUGvvosmeb
JNkFPP0pfc8rHWPwFn3cbhObAlHY9pvtUnnbq25ojyrg0WYACvkWt2djslFkfgMZXEMAi9O3CSYK
Jtm2opWspqqXHyAb0H9P+8+5OaTSGDWVqaNYTiNdmelLiPShSLHEDOxebR2BGPtiRhsg/UiPHRJ8
XfUJ+NShk6B/egU1Zi1cxYJbS9bsQvJlfcQWjdwqQMO2pa/5JpL3k5GFNzAPA+ecNnuSBaLGm6ZW
8CrZ6jfcB1HmIBPsQAbTNDjIUlWPlRBusdXLdIr1Fw4m9RZdpUXGnz5t49CnrjN438UrZo+CoG0A
RYhbqe7RtKLREPtg0dW9M9SfwXB0Zgi5NZ8Zbfb+q4DjKEa4HOtFvvupBuyZvSbgswEgT30wOBnK
3BYgtesqqNVPEBcF+0fBptmRBQUemoV8D5fR6Cpv2BtlZY6LVXKgrj3vvgMPyLaa1R9KGlgGQ1D9
H+U6iICAY5QzG0g9IMLmQvb7zMJtd8XgsvRwu4aoFn4CXXnHVserxa+wWXaS260LF+yXPUhPeF73
M6XcegCYLznnDq1kbDiooim2lSlHaQRBSgatIksDzHWUroGph66EYrgARpD63m4h6WklcgWq1rZY
nlOeqWddTpolA2rTgUwUq3oJEhAr6ODD6UIar4ZFfEvaCd5wtdT7hOFJTA7m8l/7RssJFh1S3fMD
CzNa9zYDqulUqMA+iGBiJkSSnoQBnaJoxFQ6VEAH7V+lOPUPb6LMvychD/wF3y8hl/dIBFsaPU28
gWwaJfx0i5W1DAjjZYc8+w7cp7GwFTVr398scDtcb8n0qdv68Bo3U9Ves1urktk28EX4t93lZAkV
pRDpVGiMY3eIH+OE/jTYMK8TeQL6Qra8O7GR+9Q4WkK77iuKWuMK2ZLFVm2BNZom8t2Nd02UTlac
oRdOVCOmS3/NSg1LOtgq3KifUC8RsnxRLXWuTrFv2/CChbvxCvROrcJU1LlIX/yqrc8rug8QO/1X
61adZbdvPj5+GGyXi+XqGR8tgWtOWO8aU2zDSGDquYfQQ9fMVpv14T8rlU7FSMSCzq7S6oDeRJNL
DEnNdmszxdH/UekioKkJhskR0WWlO6jYrCOm4t7v40KdffIgsGC/LBraFZYtAxbTQHpor8HvWt2R
kXx61GRvJQliKs73z5zp0HMGRwNXbuflSQ14WNksyAG+cUua18OpsKl3Wh9TWjbpwA5IKkw2oapl
I1NeAqjpKzNVHf1djx1z9Em0NHdQ18lObie/ObRg98T2rj5Wmveaj2RuOISJ1hXY3DjBI/FdR/+A
5gAc50M1na76PFJvrBboR+ieyzBZ/ZTVPQrePc4pJa4sM13X6if1qD6+FoDl073RD7mW/uPt/Zra
n5GOzWoGMCWJrDWGvt7Xw4zElNcx3EJRSF3QYKNqcETkx1QapCjCoPC0lz7vcMAByK5M8hmQEmiq
pbSGDIw4uitIuvy8kvE8co0+UNSkewFd6vP/pZ2B5JHunyxv7D91tDKdva6x0R3eeeiWaviBIQej
5D2NrMtKvtocrkRcT8umY6GHyDbaEfLSn5tjjSVPkGg00X0RuWbF8vKIIQ50r11KSgt7KfEQPPwH
8iVomh3CvzBqDLRB2RxW9XpCsL3P/XigD5C9ROOeX9oFK3EN0yqaxrQwcg2IxkLi4pVf0lXNJ5JO
lK9Bg0L2jKAYvcxUFtCyBFJ6kyyoySzRwrbvAuah3AOwgxbspmIvo1TL/2EYWFrRLiQtLzPBkgp6
LRY5tVcKhmrAjDcqrTJlLXMUYfPUTDUDLgI4Y3e2VBylFnbcxa3PXeyvjNINANp/4TQ52TG9rfHo
8vCye5bdgI7f9qqLciiVEHI0ciErjjrN5P8FL8AkztgKz6Nja6ha9TxhKMCHYgtldDKvvguZet0q
4Kqti+yAycagiDa9TzdZ5a1Pkpvthhvb2FyMXRRYI8YIYBo6TMPrYTFDEQCIyF3+uaF7yp/nkTKO
i4dxfqoDPYKxi7Tlif1V11sTO1fW7d1/2kkrdjzlSTd3UwVgbG8d5yQGWh8wV8eZuCM8kyBtcrqW
nSTlmABIlpbXJVf4ebmi0rgIRJfQKLpkBg1kiGfigBK+BfyazyaX6YVws2ADjhDEHCnyY13hX7oq
HzpR+gmeHPBpTZVB2Ewfv12b7KpWzowWHPkD0w0fIgyuHa4vUFpg3B040IZ+LEJPsUyW1ykzz4D3
I10pcmnetjGTHdnNhWTtoeh6Cno2OOS4Hw75WyXGJnkx+3GbWv1T736aBYuAwKPe4mLwDV1F5jzX
WlaIvv1FnhIefkp6Gea2yebLgGTd2OJtFlDb3t28H8rZo6m3eoHG7JyUWg5bGAh50hfspNxWvrqK
IZLmfxkSkgFPsii2mSi970d/cmzFFnFeW40zuiXbcPK8DeNjy8SzluseRxebjG8UDu7tnF/cixnx
MeD/yTnGds0g1AbiFOsLO1bcPKyhH77h6J+g7EAJoO839Hout2qsx6YUZ2dL3LJysmP9QrmRlOMh
7eDmghFj/oBdQENcrLCCj185NXvK4vxHPXnA8oqGO/IFSAE8x6f08mg5wFtAsJbWWEwSl0fFaioo
vNvXjLgG49+/qmJCwYKhDhsYYGQY7Zxfp8X49L1AqYDgDLaRo02i1SL0KNj2iem2dXvklq5vHux1
jyPSUL3aAc3vKtma2J+EjgLEOPLlh+0ba4UrhrCwOP3YvrHBccYQAze7QNyQyRhPpbgKGq8v7WJM
oF3JR9zeJEOmn53/RRUbbPniTI9FvqBSk92VUlRk6zioYxVDx0bAJjM3OuBSBbYaqE7718H1Dpvt
GuUxZ2GQL267QB30hq6TzZVn2PNoE9vhWRC4eEoCcewlxcdvHu0CaCytvNKpeD82hIT48u2cspn5
L2/fuKaEnRGOk3I4KI3ZxIITiqipBNekfg/3TBtlwcH+G3IG/vc2F8BDwPUjDKc8fQHf+wEmRvjl
/ebOU4ulfLEKlv4PXCww/tjtv3RZQbEvvSe0a4ml9FzbevSKilU7c/oGtzgvT7AjI6bI2xF3vw/H
LELBPaTuZLs772etRUZ8Gzsiqg+XOAfreBqswayC3EzKM3CWB/nZkrJ2jhyegk1kuoQHXx9m8BUF
KBGcp1QBxE2Xud8NdvD8/fBVz5W2VPELRLOT0Q3hjiGtf5xLCKN8KlvbuxN/N3iheBzLtyFK7WiL
plYrWi0tkcrJBEp77Vk97LUUWdywIsKLp4e/Q1rCaqZkaJXyvcZ9cGKqKGVEPHF1t8V99Obnkuz/
kKLh2aYxLNk+nVn2JN/eMAZ+FvlL+f239tMt1fAVG9n6DfxDX1abvFAE9ElSaR9y8ENw3owVYqGm
ovpzV3jAe2ipyKJiB6c/xyxRRsc+nE0ZVP8b0UzhfwypIQunQzDmSIHAWx8r/Quqr6UF1ft7/QRs
w3lMYiNZ50iiKtNE+lHv+LhgGVZno98CpgV0y0OblLXPyJE8m/qPot9/WSyS2FhbqpE1gX8e3URc
mp+p/ZuPzP1nkD4EYmp1NyCl0zsrqHj5/2fVQLu0hJosZMp1f92ldu4xkV9e4VqaRvxP47Hjf90p
8yFIHvy3PMZ2Bjsn2SEZowqNASpdMVDN+5OUSNc/Czv9jTTpRSt6vWJfLxIhRkT5O5iT6TiBR0f8
OrVBPCDSOLe7M/9B81SR7BvICxE2RwenQ3b/qkwh6/KNxsVpFW9g1mbIXZyx5lAhfX306U/rK5Yu
QdQRr124JJuzKBM3r7An/TXr3usHn9xxVj4GaVT4K2bh0Ynjlp2Pttr2GE60ORrfjI3CeU6l47jL
WB7UlPMXaiq0JEAiH9otMEGUaThPlURiDmHoEv7J7LrK/pifgbAg24XZUYynWIgxGrPzeTfltO/u
/eLcmQ73MzOD7l/5mUlmYv+i5pz9MGokuKVo7zj9KFYwBQtCEzd0Dd4yt98N+X7n6awMnfDMVLIu
IepOi7XJmP1P0eZWYxghSI+IrLX9LG647kBX41VX8pZ9wHn5hP6ab1lIAixciZFZ1gk5kf+zNylO
OKMjZaW79hfWBxoADfPVzrZt/Tg/1cCu19xGQy6U8K6aULBW5lCE7YD+kjtWq7y2lm4/7w+XzLFX
FHIl4SLwgdxIDTQX/cmjm/exMBQRsB4Xsjfy3h801RVcZUh85B38/h161sSWJCf7nNyMFkNNTxzC
XQoWMB3QBqSDQ6miid0kPWfRbyqzKTA7rKRxTMpr8YHDNVKGbux4XEc4BpdT8Oi84QNdDMRC67VV
g8Ti7SCRdi3SdZIg45ZWhlHA9WPP8K4eDZ7sXW9LS4ulS/scSdflQIxVuS861dm6N+jSJ2kJn3wb
pbl6Ls2ohimKiS/t+Cvg18ckU4Hv+UVWSu8FPmwm7ZkBTGLxT/pZNb82GGXbQ+3i6xr0Teee/Igu
zxk46rgIEAoUX2Yk7KPmqpNGKAPhCJ0J205aTOCb8y4L1hg2aJIafhiB6iCKU8Br+NinMFCqZ7rW
Gw2vk2AF035OURi5Lypfc9UtM0eKdsxPJkaJQUsLemL/9+msmF4vhVc0zofmvvkHxG9WWamgZ+p3
VSuicjUIFghlMjxucyx3WFD0EImgmXtV+t0LFXVUbZAWNweEQYnx8VgLsp1eT+Emtpk+8ZxyCHJO
pefrQzrl7ftHZOatKKYtPq5wBdHPibbx+W+Nj0JFvPyFcF3xpW0vHAwDOaefURoilscWVSfJeWLP
1RIabkWRqLvNJXL6oIKdchNGyoiB+nGoo7ziI9adoSrAlkWoJyhsf8yF3j0MLPv9I+qtdBzNfvTE
MmSGjeA9Uyv6xUb4ZRPXEBiUoiRoT3WjatPSw2qpHliSfYdukGqMtpI5BndPl9WNZL8/XH+QaibV
cKlgFv41dnONBBe1lr0O6QBMmrNxRXrP7YVBxGvla4YEVUzFpP7vn4Ny8Vr4c3lfQ01NR2OIW7r9
LvYA/h30qJj0Pdwayo9z62nb/JMI9GbH5m/V/oPwXhuOUSDDyxcuXOaV9GLBGeTBJpz0+jLX9otN
GjOnUnDWFOunqKaHocFDB+/vqEdSnpiYDN0sebXfpd5sIeJxLloZFIqRFNGuPmjcIiAPIwTng1ye
mezvK/TduZSFlrqNSC6NtCl1XGdD58MpF7NrRYr0OxnRbglRS1keGKprcjgGOojoRGfEnrZWDXzZ
NsvJfuig85r06BDUhHU2rHJvVfQZ27rWDl4pPXqd0roC2tLZWxmlkxZLhApgTDrVuY4mBKO0FQzY
wvJhQOZTuiJrsCgj0wTXHLUajuldG/LYccetTuYTwOqfkzyMQEismgyiPC0qtwR/xOeFDlwPY9FV
W5HJRRbFoJSxVaAiqOMBdqG9BCDRhxBkTr7ZU4gyGpTaK7TqAhidPoC0Y5xG/bTZu/VIxvUUqW5R
tzj/wwBVM75ytKMdL9n16jKy6MSfYpYZSv5LxAtsHV3fZEEDg0XFI+D4KPqqdeU41UK6VZez17GZ
HKIc3Q/T1bhExmi8AW4xue2MCZgPVZlXVESb/AO6QPOZyTbw+KMXwaSUZRd2FtGAWGbUbL4g8jMX
9LUT2z5rvnO1Jz74eh2JuHo4apKnBM9WdE/tOF4YPFAgkzWML1lfILZGU35PAX52l1cDFnb15yFN
YgMUi7lM72ZcsmR6Njx0OgylcpYFhnGr1s25pMd1BDCSK9pvIUinv420HXs3HQhLr/znZWKSSGDr
a/8XABpzpEUeRKgCVHq+Wr6MMnARd5I3iYJQaqE4doM8FFdAu+GjbxejAI0/EIt+iXZT+5gfEB5/
NSqlXOxiQQgSesms/DIXbNxTqTybCfmNJSWkMqmL5N6WieEEmL1YfVp91oT8XV97JmJMYczhRDK/
Vrd9v8ihQr2A0K/TCQDPvCtEhnuoms+3v4AzYue6LJSw8a+UuOZDeFNg+cGaG2b+1NBLJM+wBL7Z
FHY7aLZ3fNaDKqNF+yLAiLcl8tdVqBD3mS+IWXbGgf5xG1EnfqOGxZ+YJilp4aCsJdgI0l0T9ieJ
W0K6eCm16OYp++pjKdVC4aVwLsgn1uWwakBkbKuZ6RZpm36PmNNsHjM+LCehjSjf5VlyqPtZ8Dqd
IAM5VXVJdsE3Ha/Mgkq8Oi74y82XqOTtOggBbxLW/tX3WTUrEgRNPDRZsFytRUyJmcXYMqr2imym
6+lMOHVTSLI7t0LQUX010XR1x44gln9mEiZ2VopqmCVSZtaZ+VfEdwtzSBoxCm3I4QscjIE+dvQu
1ChzbSMQYTbOgzYrRyiNR2XNwIOtJ0nWupVHryDxqgejzMm48cj2LLvE3nI4yQgtoLffqYHPk3WF
GFG2WUh5qwt4j8Hgj1mXS+ftNQigQQGPK/QgEeES8Bi9XHLYa0LN9aWgTNhpBPMvSAiwvxDrIeWo
uvobR3YihBOu0mIViapIxGSxideLHafcOEjCyecZhvYH7HlNkqmajV+v1a8OKh2fDHbxLhwce83z
47m9X/FMgHVhkPlmtVZUnmPIv5GZv36/zBbB6yQ82OLfxI4o1G4egG3Mf3RQ2txWuWQuso0HSVjr
h7fgNwkrsS+TKjnFxPL0A0MsgYROwLErQeCgV7oQtAdp95DmTEP3Gu1BNiCWjF30eSLU2Z/kP6hi
rndml4+MBelfppvON3T8FfILsmSjBugY2hUUcTgapmRM1cpr5zXqMPdKTK4OaCgrcybiE4wuWOIV
FFK8DIee98W6rK3sYYD7MebHZS59oJmJyMbR8G/7AGZE3gnfUOzAm7E5ylYmt1pdnOr9AujRW6Hg
lJ66ui6rrVbDvGEwVW70fNR9zyfIg2rdYqXRSmuom9tHMPCY/FjflNpep98AivynjlYPCYyJ9W2r
NVlnBjJ7SSbVwaPC9OrjDGnia9tuYtit+92qpDu5w+ymqELGxzuDgqUy4AjJjiryYb6qYSk8bxLp
fjjsSN0Vtc34P1Gj6e4MhgQF9xF0TPWiQ+c1GCUVIxz+xcZqN6s6H47WoNVbiTRdwq86RjWfybKY
fIkqDO0iq772DXjfv6cePreUFqv5Nv8WCcURw+Klv6hIu7aTT4fKOyNiqIXeC+xpgoHCSQTw6hTn
qUh4yJyvlR5ySEYDaIFBmT7FsvKJz+sU27UeWECBuiCGs14BUER9yttTV6YHlEf+4VTUcb+ackh3
2sSdtQgsX47B7gEPhBiULwUy3f43QOuhksgA00dTjXjqChnD4Fezyn+e0uDNBxdGOttV+DE7jg9X
XbaAF8rZyoKktv2OXSdCo70unxU+Cio4D2UKp8GTezurBhboBQvWGiMpmwVYFoO5NMuQWQGNiLmq
rxEOPBULbsN+l5VvWWKtF7JPKoXfRaN1h7+4C1ie+Eu+yZKWuktkpMpv0TCeJPUqaIXXxhtrOjx4
MguCavVXEpXujDCyU32yt3+pS8RP82yHOHsCvgFGlW5wOWRtrSWVicbrw4jreU76cRVqRUpgX0l3
efVKvbsm2QGGyqsXwTIzNNrLNqGPGKEGnQPfxj0wnugk11PTM8HhAFygQynxSVGktGa7luprHXBP
TClHE71lc8JZ+y4bk6sqCt2PgThLi5S9c9M3czdKI82wmXOljgmoNluqqEQTX7TkxaELFEuZyv9F
a4f9JB1gZY84PpifaaLvtJpQF1N7kSnJYO/AlVBlsX/g0X/sQf6P92HG54K/lkG82LCEpdITU0Wn
ySRsT/mDPmTdTg0ZeKRWRXFgXGGiKBPBbikaHhqVrFVITHEKiGTPiaT6aPT6U+A59dBOqMlmqJ89
7KSOM0Z1tjL90nWgqTaHg1hIsfr8dR5DkrxtmD+sDvwv6TAlMzBcHvi3FqRkrflORe2IdMRXjiii
ztDl45T2+HYwqhZ2HqTnq6T/1zp66S9m9gb2GS3lhdL1M9kJ5KNSIr1pgn9lFFFQXuk9AULmxYXI
QdoQHgUF/P2ZS1ILa7u0kA9z7npmIWmiGIvoIqP4b8WNJG/Bvj0q5PwdjUyeTfZlB5anc6BbRM68
+bXO1RYaRbzaJ9GlR2mDejnfn79w9q29gj0dB1Z+pkMTe0LlXJ4a2S9xMErZv91XQH5blegKkEgZ
CdYkj0ctPXm5YqaD5tScpfkPNoMvpnvipOODQcz9qCJU7fUY28oouTsUZ5G/YQKhz4vgYQuxu5HZ
zw1aPuTRu0IjmWPiOo5rls6+SrRSAQfLiCy56S17aL2K0PDBlW9Ra0O3qx102nlGi7KMScRcmstg
y25p2L8l9s4TDyBB9QZKCuhGH0EhFR+myfstJaZetkvWMRunimu3gpnYKFol9PrL2vEfZD6bB2uJ
NACIL9kvW7hwt7wN4ZppNDcpdyAycrAxvXr84oPW6F4M0s59sZtCgE2WC50Dwd6tD61grMWqBdrL
NBsONXoJ3Qm9k1TPaRLaqncAoUnr/PDbbdDAWXFQZIY2FDq8y3qtq3Z/U4y6tShTHdfupfYsCOGa
rDVZAkyBfVzj9dkNxgc7Ha51pdkVbhYt4ZrGr/HUCEJhhmxg4fNY1eiuT2Ry+yglPBhtYzmCYWcc
oqGSPqoMtGk3liR14E3DcUUud7tII8X2bhZC2JA/nqR4tUpbwo2zMett2+G0jCBoC2tYh779fS2u
NZ9vHK8EY6Yu0IL/OPpXKUr4Gf6mrx4cgcAsh1IyPfsOLLXHpVRvFM0oFOuljAbKPkrrcPFXwdSS
9eiFH43XQKlcJAtftWNUO+Lodxh7zaSrNbz0j07oF2wrwe7680G9Pq6rcTdX2peh6D96MhOQUas0
ZAXBQ3qy4206WZagNGMtPGTavMXegcfgahgNsmuQZfJHiWeNTVQOjFZ9S/WV+K6iN/pQ7fLKO2Fs
btNrE9P/hrHvlWDaKnPu6mrZolZi/IiYlohHdF80NOG7P6/sqUOojTyskYgOQ4K8un+Fh9oySNpE
3WYteZFdQtsw3p3dCQtmKU27BTMGOF8f3CRcLbstXC9rxL5wtagpnbvhbCQmV/jTayWtNL1e4zfj
T3ezp+jFf9QHprT1CPY61xosoUTyzmDEwArcNCykQsZ8IVJvpsbCf0IKHOsgLITr6hp5UJnBJsF8
vJYBiDNjBFOAy3Z+job4E33up30mdmLH5ux9vsd79BDJidifmdMee/jRpeekdtUyBPmLcm40cduo
SQ5AFJx3c0DViYmwkhQ+Pw8tQTcOvj3L9Tch/pvfSBVxjoAiU3v4jybb9QxzQc7jYkVt53pMYrvS
22C9/Barp0TMlU3lm7zowRUQLvdw6iKRsmn/D04OPbavju3a772edwh0T6HW4G5AfgtNv/pMa4N6
yjTI9lv8FAPYUgpXTZ42S/QedfQtokoDmLjnSlbda4yY86bd/emqS1yFPJmc91FJN5hDDB6U+d/B
n+ri9CzbpLZHAOcMFaInECwXC8kav+mxi8wtnU2wWKA6KUBJOzwtXzn7b8f0w4dLcxjMGJ/x4LVz
KzAnp21BFagyULnHDX+JDK9BvuJ9ZSnfzBUMC+pCQhjmsE1zBwBi6I5TqwIvm3i1UiGLhzqyb9qd
l2yokIyLmMUIm6fOMmQOwIZpr6D1beXoPYFV0Bbv0+WFUe9/QWAaaezdATKptKchENkvI4KgjTvj
hRurptKmTLCGISpHNgfD2n1h0R/YoEo8Z/9D5Q5X4i3014/gFZ8N6uOCGFYeE9emaUFLQ5Utzcth
JSkP49ULdjinkOK0/6lNMqb9TTg3hWDtcnPBmE2AFCszqJxaQhGCfdXHnabEJUNU/2WGrH/ZMcd6
vq8hZ4MYuJXaSQuJ6EXn9IQXAvr8Z6rNY3HSXXO8T34wbjURCdXBk+gWkyDIa7oXjTp4MU3Bjgfc
yx24G8n+jhG023A4N/0YLfZjYTHtTXVUQo9yxPujJjqf2xj3HUV7sVdVJ+RbNx2YG+mWWrRLDIxN
70OSVv3oW7LAOznNK3Prgp+whYulwHj8hb37hX5IBM+HhDg1qU0A88MxqcnFz/EV7Waw9hW1pBCd
aNXskzGpztMYmo7FZbvO9QWnqM4a/1UYLODr0izJ3/UMEbp43ACl6z/DxFWJLYakWEpJgN3e+Mac
wZIC8AqrR5TCXRECN1wIlSMukNhTUN/2RcTN09IZPTis1IARG/Ygj0ftfxa3C/Pedf/M8u50VrSW
4aq4n4h1wu8yoqjWGQusLRo3j4NlNm5DWLuw0HE9qBfPsU3RhPqi2eHtxobtN4kKarRk7PdSrWrX
90j0qfcIlUoEVEZoF/oYdz3JeEH0YWN4Kf1Xz7fUxruv5kdX+/YmbwmAGMPhvfWjvUVzVb1zZjfP
pY1tf6SOApycj8F+Oraw7ssnCwRIJQOti5JRul7W70bxIdr4UJ7NzI4hzPljXrMRSgs2B/U4vfO4
vpmXKMK8zvvCrGage58oeI2kUmHbAAed8eKNM5U6RU2NK07eFi9Oy7v6KN2k22R9CGd9LGDgsc1t
vEzif5S8eh4bXEmlhwWgTlew5WkACaK4miPNfV8i3DqjeEFA5Qbrkfu6m5gZZA3cs6EgKTn5BaID
VAXd/Ot5sNnxj45gpnhnJvkCfSBB4gncyZb7RL0wj5sZi3Lf62OcE5fM4/yRy7NbYsH4n5BLW/HZ
IgfJOhI2jArO0w9YpbCzlLWhVPg1aSnQZ7Bb3cjPa9hjRIJIN4Er/Iyzh1vYqfgqI5tHXkW72psQ
0W+Gm7aUteYN4wRt/Ea9DBMfC91IzVBZSd71tMy7HMDQsf5gcueiNkTtTPRc1+qyTAOcd7tNbkkR
QfpbGae3rdE9UumTmjpjHOAKGkZDLXE7EYn6k3kZsXIu2XVcBFzgoa0yHVjwIe0oZhl1c34pohpJ
hifJMXliB4XkeFKN8icSX8dVIJCcrXh+iNPwdBj7AkYImQ+++2n16egSar0eDOtH4olc8mXKEeEE
Kpb4eR2KbBRxOU6mJSXVUL4pYehguHluGxbHEDJ6hXak4PWiaQBYLeZ+hkdm8qphKbbyYU+PNJqC
hYOYjqoUYx9AzRh2DiLhiNZ2kPgBhkKxtv2rmjcjeIYHvNvHre3LbU5wpMjcIGGrCakkuXwMuxzx
cHvDrepiTDQQWOAQ6GfjZ+IjzEeRtcb8vDLc4x4bvi1TNPT4o/Ik1LG74Mae23+S7+WtH97Eq8sz
TtqbWrkvUELrcicXSNnYOHEO0scgupK/tBHJG+aS4SDnI7Q4OX6tCNn56BFdxDU8oPlvN4YPSAmJ
yk1VlIhau3UU9Ug5yDY+fHLjbDa7O3efuIumkL5qrl3kLipOM462NjC29Zmfp8Qygn1+DuVrl7va
y1b2EzAzQ9dDAfJDrPIQaXSjT5QwqaaYiawoqOkXgNJWGtbiB4drRSHHZNc6cBClBC1Ou8rVa2w/
dn3g3BXOBbHbJT9bShPtkuD4fr8U2Z2Z39hWuZPm+z88mIl6IxS+L/gWNfCurs9TytBywCBVW/Nh
hvSZWLPl+BZ6jShTXRyWh3wcn8/iv7dd+dV77W1NSHVPWbunsYzEDxzvBoGLoVhrlqNQmWr8ltCx
JnH4Y7/UREdR5zgOc5eWGcdi5uJr3Z4SLBd8BLWyNG9umngzploZq8zhqlW0oYUYI/2a0q4oyzvg
VvbCbP+5l4kBhX1p4WsFwt31EstRzUngYSOtbvL3es4vWm6zxvHmssYNqHxfjcY1wXyy4IdZ/vwR
yPDE5l12m0ZCDuoOCEUB9z7qFrm5oUNDy29ywWpnKh3m0aknhvSCJV8IjKVutqla8IO2WMJoJRmv
0f0ywrQ73vrGJRc+OQKUmRv/mWzmCXEmzFg4teZun+a3n49ocPtTjAF1KcG5+D3KHnbLVwOe0kiP
1hyFVIOIeBIq8yyclHpcDquw5OT/WvgMa5YGOMWmQArun6cExTK6a5kyEETBM26MeZtm9Vh1Cpba
P/A7Es/HT6IwSK7uonD+FQMS7HNJPBaSGFvHvr5S1Gxn1T0RCZ6hDmICxOvL1oG3aURwVb4ovw1r
2XAJ43oy7azTjpuiPppDIf+Z8CFnCE8JCyuU+eM8CYBI8onhpM2vDyYsq0YzAoQ40aBSt7B38M57
TAVRjG9BB2kdKUBU7rP53dfZLPpSn3QyooSQafzoVrf/9qGJ+v5OgGD7r3xniX+bMP+NbLpmNgW1
pndxPRVGpkw29hkvv85/7INLhGZ2o5IlQdLdgFsfQHOfAzXprAtgtpRdjOKCv8tTfUTEKNzJ3C0e
4gu1F/d88PXmOtT4sBqgW7/Un4N7b6fjDA9Nu9sYfu8Us0rYqa+9aGIM9m5WVtLq3Kvu3jCOnGJX
smCtgJqvFpu+JCR+R1WCi+IHNyu30r5GcVZ10DxpWe0eHAyIRmvN9QS9xalB2ZeQcXsae8v1zGP2
iUj/bzSRbL5KFWo4DlFn1tsjLiyMHWE6PHt45Z3OOtoM0w1NzmooDXUMHipBF23Juj2IMD4l5WOL
Xq1g/dTa4wZ6OCIBIVskydqWygSmTV9AZFe6OtEugF/1syI5VvfnlyRKa/eZDaQ7CBpuEOoiMaCk
afzI3TUi2gcJVmYEfJiDXR36w8oDkprXYuPxz1tH9xrFTkeAWA/35DvXkpoK/M3EVG6oHpsCJHEM
pHhws/6EDU2+s0MBu/WjA+M3YYBVj7WpjzpYaKRaCUn60PcJ1YHr8W4/xfSn+T4aiSxpwse7FPeK
IDb6eqq4WefLRMef3zs401r4Qeq87IcAbWagJ3adMGFcUcbEKcZuBb+SUUAcJZfniLo7GnAcDv1a
rMiGfyam54iSOovfi75PNUrdS19gTHgFXIb/Gug8Wb2LJGDBYXHe9zAq1F1uIwF0qbti9tJnUBT3
DmYMLtdk9X/Mvl8M5f38IlQ2+HJvpTZVUhFiDmdRxvyARQ1OFPj9G0Mnqs7TfeSfLLtMgbjULnrd
FGLmMundxdy/ByEhaaPDRpRqw3b8eD+IuYgxx0Y4G51cToxpMrnRQb8XA4OaNMKOtf+acKYC6si8
KIm/K1+AK0WLc6KEKDT7Uw/7Fx9079bzlECLIGwAAgX74seyf+rXUhwkcwlrgAKs4thXZKPz9azU
9PjBXZAEIh1c58ts5N+C5c8UesvRqJPkAuhoNe+V/z4tvNhcPFWeeLQzXCiv+HDkXq728xLODibV
CT7P8C9boIRMGscxHlkLiAmF48vZ4s1MO30RTFS/bP+D/MERhm0uoTLFecTYWKVArbxEO+K0vzIc
tf6oHVHxFbmVDu2l86eIg/YZWLvSUKUY/jwozNI9yfX8/BOcT1QqLA5qYKIm+Eu950PFSaWbmw2T
dNYBCOzCAxJNoOnS/NC0G9NJyVj3Vsr0j/Sjzu03iGpBKNYHLXJTACcW1shPeGe1kq/NtjQ2gyrx
pYbv4d+kWJUv1q2Y82xuPv0NNUuROsFw3DABM7DUDP+HeWhJH+nF6c+THNOlw4zPYg+FTfxcE2Ou
RlkrteG/dsu1NIgw0T/S8Lsi73FdNrP0MW6pGZioTzK3MjNV7bOfkwxXVFbkpYdH0+fWRyVem6ZH
tLyTb+Q+27JJO2RGn0gVg1nLLOMib2AbAjC/PUbz3vXOtJw9OcrXK4Qg9lJnSFG3VykYWv/85fAo
YrkKf74a1FUp/Hhh/EVNim4YFZa1H8sGORpowLu0Fyy5A15aE0mvMLS2xbILrW+36mPUc6+O4ITF
7txUSNaYeIr9WWw1g+Dgd+luFBNnuPc+IyvxGMr+D8nTQuaEIHuoec8iXHmZaSu1rl8bi/Dld92/
AhTKytyXZHYRQ3p/bbYoJ89SsTheCytmwK+T2NF8eU3ycUb//92y9zm7iqQq7dCRsAyp+rwL2VUC
Tb09MaSeBQTlzR7mN61jyZ8lhfJE2yYWI2g+WupLsR4YkthUC6lcjvbCWF7IedSz/2bz/GGMPfn8
boK9aPs5UM3d9YfkFz9GWTOGin2KeSs4jp2rETEVIpFbjLKK23ceGX9wzFZ8lWOnxHWPFt4mTian
OifQYtvV6ozQ/bPsbWbeUxdyQmn8MLksu8otTTysud3aZlB8r2tE0zKeF/CbbpOTdzLxevEzjxkc
CFYzDnKRE3glaMhTzSsuuEzxR7QMoOkcAco/+JtnM6j15K0ecahS6qQ8ZQhBHyvvknqbrGy968qC
WaQVeRNPuFB/k5M1iTCtdKAGxNIsOe10bSsaM2yZrYeur9p1QfuPsIZMxAUfmr7B3YNp3QMjlHmH
b00MLo6OnOGRUJuSTtKV1n8e9YAgEskt47pE8CK3wfH9AsNg1zJVuyChaK0QfOVa8zSLnzUgVKfN
0NhvFVdb5Qbap+55WMgH+KmSnMrPydZUg46iL7u+O0hvyQCEr9HCnWOZ0+JROUaDXbWZAp4mCuhX
qNKpNhzeVwC00PUugcDPyl+uAUM5ZN7nXY2lJ4HrhD+m9ZlHWgCuf2dOKeeQcveeQzsl28v6XmsR
EIJEOoTnaVfN+Fi9DKSWeTo2M4qkZRZhnKs6AEfp/i6WQ1MTmKE/f/e+qAIZIYomT35mKXJTyilk
FY9sSnf4bIAbry9f6QlxGZlq2f/QxMxaAX3vZdQPV3D4FB2YGzDVhV6egL7BAeuv2iJzemT5XrX0
8GE87nv4XKh22+ZEq0WcoUpX9/7z3+SwzQCmtdBF88+zsRwvuV3RbQuY2ccBsHO4AbmbaPx+xo+q
BeUPNddWkx7WPBq6CE7uwc0lYreIYGeXGUt/4foQwsN3OyptaDgcdkcbqe6VhzESZcvb+/jFWeP2
roZdxenFBa6c/4MvHwMB8/MfIm4DoxBmtEBAGtbTnwwtWc1C9JFjLwdd/rlG6yCwJWVpyY8t2Qa9
dU0Q6WwnMYUR/py2SsjxfvQ9b+15Esl0onn4UBKwfwuBIhCFmO38if9a6TTvJhMRa7xWB/Zs7KvZ
26DL3z7kqxFUeIhciAlMPZdxGvqxQus7QFM7nySAQQZXYbDn6x6zS+P0okxej/xqPxIaNIQybPh2
XiUe8gnUioJ4B/Lypa1avyV6zTvN5y3ZQpHhqJkDQbUsdB7V0K8T3EVRr003XvaJ986LArVzcYOp
P3UGMapdlPXkVGwWYQLHm5qGakr0nxKs+gke1dGGXAsxQNclEizqppNNgoWqnWgdT0dYA7d1B+HU
z+7KdIQFEYG2yTSC+nBFzResLFIKrzFLL4J7Zeqn1Yivkyuqymfg4B7mw8cwV6c3gewevl/bFsb7
OclgaUiLKok/gvP1wJFzOzHcC9f8DQpGS7yBhPpe1gn+3FL6TAS3hGUSc0s3tWY+HeQWtCtfpeg5
FK2N6FRNaJlvoHnDPI7DeOImARuWdNQhsGKHz085j4nQBGp/9RRUDs1wQiYIShpOtZqYl60Y4zNF
qlmU8+O6k26YuUqsj/vP+w6t7ba7cumOwCKG3akdp1vDWirG2NfC6HNrLpmOs1b8U4u9JF0udA3c
whIMy2hh2IqvYBs7di3QIxB3kdnGp8T9GF/aBAyqbTBLWhd0qtpBDXPWdBiEQ7eCQBc3MwU1OUpq
aJqyr0qiu7REYEIeFuSIJrq2lqki6soudixNODLbyhu8LhFAAjLS112F9skz0xFfUqdQj7hyxR6F
szwkGd1E47zQ2jS2m0itBFn8f1yNRqb3bak60M36Xe/9V4onqDj5xvNiFVFDhDIuAgq8b64NaNrB
dSj1oyqJtPWskD1am6s9Q7VmoFw5LUxOJbFw7llw5yTU+lwda6CFTdYBvp4pchV1KdBu4OKLAF9+
ljhG3JO1VELHL6XMzpIKryIBlbsbXMH53LJMTor2NsFlna2cg1CCWJLDg10W43vDOetYUIGwkFNX
DO9USwrNRdWSP1CH06C1dtjUN92Ys3wx/Hzmkyo2kbXNgyOSUikWZGnu/jKqoT3HKn/gxGbEcE9T
q0W153NX5gQbyJE5AJ7ePt0rWUheAc9TF3o9qlnjMoclqzpf+++K60FD0iqEQ2V8tbPyVoyJqidD
m9agw2HRSaqdcT5ddM9vZrZ6k8dPr8L+W3HCbHk2oCmZ7N9kDzR1pv3/KnpYAC/L1L4H1KZFIqjg
s7zQQAKvbJ1gqZtfaUBDDrfSaIH1Jur/qcsULWPEvPSGWQKBkG9v9/W8s2C2gw7QiQB9PoqmTpTT
+ZKCXyAdTDl2KH6d0O9V3g8Q/UB+gqrfkWRh/JKXeXMiM4I63rQbp4hATIjGEqIPCUTjSlTHAm86
INV9w5ytzC+NXILtai3NYwqe5ei7jzO3NRS4pUIxN8Z9U01h9YYZ+s2wsuz3UIN4ULeKG4K8wkLO
qcBePiilwWI6OEuU/OIKm8jv4NRiDvELbNTIgm1Fx7ZFfGit9ItNcZ2Y60X6E5nSz4bc8vDzE/JH
pVags5rrRHMQrphjVX5bPJy0bboF8Q1c0MwVfRe62ryu/Gbxh76r5rl2emYFX40ElzirbICUy03g
2KHcqBP/6skdJXBtYcvJDJJOUsIJ/jl85SyT/syc7OdHl0BwvBDfGV5puwmDJilkD7kMUw6dJ/ua
TfXF7w3zJ0BL2h8XumesQ/HIy9e9HWBylbO9p/y0OZLlG6sUC04wfJPSvdl8wqCyDrTkARhgY1+n
TORCFJ4e7Ti3T7qqVSjJ7UwUlDZ+MoS0FW0gf/M1P3BgvHgaN+whY9EAh0dL2N4R8btazrgTbndM
EOFoMnV/6pAeRpO+INjCc/bsxmtcGNPAMVPQYkhoNn+WngLUGe1HuVImNl+3sNo9dgYfou+IAJD4
mlTX0BrQE5cFY3bD4hxBB9NNhRzeFFwRQ+/UQzIndUovC9QgMzPYkomXwUkvWdERXFIU4Pr3ZpcY
k/UGj8/3Sz/gRJhsAiR0QUJWOpGNJxbZicyc2oASyWvNtWDTMOld6yMG1ZQ5XCTy6cwyquH7Ob9C
gN6AuFmyYDWgrG1efYXMvgn7Rsy1PvsPWIFSMOOqtWZCPm79hLulsPqUs+OEX1O/tikw9LE4EQ2C
0dXtHIgFmMhQ53Vwz2CoI8BHxhiopijWaznjU20vJ3VYKDNy0c+FNvM0k8RTJWriyJ7X0XK9NI7u
pfaj5sOp4+XLWnbjK4ciNkUEspEkwXabMDrJkbcvBzCtfHJuaEnQUWjzkv++XcK43AggQB3v06RI
Or+gu0cdPXahc2CSuFRwNuts3JfTPayMKI8Bo7Aya2w/GogQtS1F5gKudPgMAPlyBxEIRpLIRYZK
TE+nc55SwVib0Sb5YlTVobOHu3lwpVIBInKC6vsfykeONGjBr4tODfV2hhgf+l4gyyZ8XeHIbYhu
FBhy0cZwEcNhOQ0Yo6KiJV3qtTQD6xMYNPHHWJ7MZdaGWF1+mN/b9YIW1ol0CPkoU9t28w7kkJ3v
m5k5qhQxT+SRcJbh4EChUvyJvSCdzdWIQL5WFDVk0izl7VfBqot2E4SejjFZb4Kby6y51iDHDF7J
vEoLkunmynyNQWdW0NiSw/gCyIcdX8Yb45jCqaLuJzVhzsbwk94xTwMRCVJcBoWlTqoyPcRfQYkF
GQ4NBOfR077uexg+vLCZ7ZqoH0hpLfY5mak9w8sVeA1ZQgVmffv9E9vPpqBHV3HYZ7VeLd/XJYiu
WU9LzvxhZ0CsE949iqoigHhcPjbTtQlkHbq5UHQY/YsFgo320wUaA0lNNZ5G9W2ptdzwlLGmBzWv
VPJTRY2jrWQF9PD74vN1HGRFk70H0/bXM1q9xP9h3IHe6OtldVLpkNae++STxhNJE/EWUDCA8kvu
WDJR4fR5D6SgZTWgs84hbRk2LMciYZcsMo3AO0XXuA0qvkbg47qtm/j3XgSnNT147gYusEo6SYmW
SXP+0p9cjWc21k7y8R7vZJFglXWnrOgzVa6hrFhaFcsbsEK5jo/zZqDOlcMoCBw5nZOBv3ej30Vt
tdXaJjcuKODv9X43WFjQs+hs46RzF0DYWe8GxgLO79sVRDfhT9lkMucCg/Q2BuUxf6TfRka4ZhwE
R1gzLyAGmdFKuvwDgYxTbNxVldi+TKWHXT3c4BxBa71xo7JGkuUGqfJdQYw4Sxjfwh7+6DhRX4he
X+558aBcWsTDth4QIUzRDSDJXHzBG59dzqb2WjXz6KjCAgtzg5YNekklJDPsCfwEo/cUUEoKCQPM
FidYJEDRnU6tFL6VKTukhBqqbi0Br/s023p4tVzsdGyc0rpBIOzQKwOl01sYJlq6A7dS1sD9Tz1J
IYKVgD8AKxF5omLkOpudtVlvqDWSn9BYFFUAyvPoCbNGr2Fqb13z4zYsyHe8DEwLiyRlGYDduTOP
kiiDpNcc6PFNCkEtFTqTt+p3MsF2nGIFizN4/LZWwIMkH2t/FhMXqVPuq20scekdXOsR3QG6sjuZ
Bk3+fzZV1L7ztikGxYGGHTaugk6gs0CKtg7MbOre3h5RvPVZrPC+izfBorlI29AH8y/8Y1XsfDWv
8Yy1CTcwYgWj3TzFNv58kcojKXsnAD31odxgUP1u4IWyPfd/3rcrhCjTFiJGKTwi0KlMqtA2Gg/v
TsMeoXao2RNDpcTUWm5YEC9RaDxU8usfpB/e4FQXcYN37fX7MmywRU8lMHWjGH2dZ0QVxDNuwOsQ
VRogp26sCMwBV+pNrkvJA64oWvk9CsHjwPUY8WENMlFG0ydignutQKg/R3NbSs0r6EUhjpFIMbC8
bLt4ax/4d9C9vzxrBehyyc+S4xFMknNUUUKYfcpmqD8olyP7LG9Cv5to2fJSkhag9DowPJKzWgnE
ED5eSjoUydRKHKgz3jJCcoPteX8iLZe9S66WG/ETqeUXeM0ye84smUKvomCoYiTHh/MZll+XIJOe
KDIJTVRujgrfAF0oo/QRwLrjJp8gDurNEZEipkoI/xjX+Es5zpdQAM2spz2myQnLnliRBFspKV0e
VtL0BWcPjfOXEX19xJS4DYZ3sIA1H8UiHeUIrH/3PTKFAf+Kxs5RVJSMe1ytOcaYARjMdDEDuH7I
Q3/uPxXM1uHUpoQfWiIawDUpXTT/ss1tjocrkyP4wTyTb2OCGiyDnTzcLRYZDwUg2B/k1TZGLGPQ
LQjrISmmQoaHpT0BtURQQXw6cdlGD/6DdOZe8mhjcukrfM/ey07OfF7m654wgxAQeRNjuw22K5PM
jbGHuy6ZzDtzq+pA6Nn59vAxTXQVA95YbJKoFn27+zgF6OlvDJw/o8AVOlR2TqfvKLFTAbuVP+Ii
fO2TcconkTaKbIvBLhrjQsL29L0XGajOfvR+PLctWxoSkuA39p3P62uP81FfqqndHNSllg2+V60z
OY4DBL5Ic+8hwPsW5BoFL5GBos8tAIG8ImaQ0O4Imjbaa7yQRAQJUTOoXYFMEDkM3LizzeeswKr3
mGhqb+sJyzYYGaAlE9BQWT+h2O0hICvSew7b5y+8rluWezk4tC8ov7XsNiFJROFKV4Ajv0bAEorN
2FUEiMUOJcICKgkL3cCKQI/YMyDHETC0mnurnR6WAUBQvhO6MtEi44mthPEvWqDRsdNSIQuKUVHR
X2f94tISVnLTJ9NzDhs6IafbS5iVGj3st8JHhH33mAV/4ENhy+Wj1SsJcxf2ONDfpZsk2PLRHN77
roixOzS4JA1/sBlXzDKe2HgoNgqLlcHh/TwQHga5TKIyqMZ3TnobfFI3mERL/6X5DeZd5neM88z/
1kYVtHl4AP7pTbWTbbUAtwvxwnBHXJZgjslUn4YdVhbA7xjpu0alv5Xa/Bep4SDgwc+FTpRIsWH9
TVU9tEKGl6ODWObW2KGGSXfB3Dc/gH5ftkc3Ilzk852+uQKA1X66H6BJVzIkTCW/rEATut3qDpfY
j7ZWELNUxoc3foBwH8bxTwX+OM/DbOk13IxN6wWwb+6RR0KRt4ihkrHHdfH3YpDwprs3yzNkgucz
4MJaihpaQ68Hcpy0eBDjeOG9SBdq/t9oGWj70adaDZm8LLa0bbF98khnqq6p1MxP85EhAzLsYtBy
T7lArhAXO+inC7lj9ag1WPdACqaDx1a8iF3CT9QA/dN146msSAnvtSpcJhLbWVOf7Ll6WmvfaM1J
reZVppZdbFjCfstKenpSbEsEjRozV8PtspPYcWGK5yDxjccvaaqooz1rQ0jB4ngmSh9k5px7+v8b
yqi//Ov5On7SMbV8C4ZKfHixTe6aZB8kp5zteajyT966LNNA6v96KTBed3aAa88am8xEv3a35BNO
aT1b8i1eSzGGjORaBMU/h/Tg71N/MIdsTA5FBPt3Vx17Yi6YKplLiKkBngxrDCI1BB6r549BPwzr
8fBFVZYHvrlJc3zQ1UPL0SP41h311+t3+xOGz4H64gxc6nfy7X/OtQXsOCg5TLH/SC/Om8HslyiK
g4RS1WwZ/uG5NO0VTbvCUg0VCCgc5QeanTgDCGWJZmHvR2fI10pi+I1gtvSnXrRTS23pQpQYNHeQ
/6RBMgsXIUx7IzUEmbS3RUFCmYZTdq0UASKrIDo5sOUk+0VhsGcThnGyFm8/Aio+IEXRjVe6r3Bf
9vRhUKQLqkvEMXT9R9OIU/bX1mgN2JAeEWZJGRWDgWKn9ecrKTP+e9nHF+VB35SJyJUfGtcnVyRI
Xb6TQjiTFdH34R0hK5cQA7edp0RhB5DTbNEar+9HkGAEdG0XvlPO53wAK17uGHOdZg2lSGtQXXf2
+87EanWm8OEIs14VCCrmbJG6ltSYgRyHaQ1SDMbZawdF5bebzjhP8iywy34MwU6zOYCFdvItSwT5
P16q5vAw9TDy2hNaWCsGeZNljlZqoeNuT5TflMMM/bnXb0P71KSw2IX1MhPKVDe4tr3GEficXfy/
dkUM+lqXX/9B3J2tz66+9/iRDGosOm5RrovqrNr3yNGXI63BRdZnTI/+3fyzhGn/skWUhh40CpIR
X4XtYBSDAWWU34dUkiig8TOYzYd9xHqIHpV/I3F2RalQLXm+NtDY733MnBposAqxrk1DjxjrrKE8
vVpCBveowtKViCj39hoAM7HbexyzsJ3Ih6C3I/Kc97x7EFKLQYdzD9HQ394gTk67a5+S4M+ZH6Hl
LYoRAKu+ugZvWcdmYI+WnbICa8Vomzh0bGKRcAwGZinXpiPXDqgJQZcUpVmXEOTBAeSD/9RJrTfD
H2l4cl5ZDyvMtV7iLsSpnBnBEqlweOc76rVmxMSdKo595gzik+XfD3HyPmSwQMwGR0dbMV2k6LTs
xCSJU3fo5yqrEg2HPAquRH6oAMgG/7eYDyIr/wxLmGRhCEE4bsrI/8t9f0IuIzH2v6LRhuKta4QM
7dypoLiD/K+bzUi+/UgbgQmxWC8JXEJ3yPSp2T4RCR20fHcL9uYCx1mYpH2awCNKf+PZonG/ZVZT
z9BoLhOfZnH5YQK3TUonah+8k412NYlVL7na7xCtE/9dBErVgVUD9I6jcjQpMjcJs/efxNhujlys
YOO9VcnjiDLlXChR5fFSCJMqFQJms50C314X5L0ySMKiwLiWLUfnIjcl3WXrUTYoNm4DfKXbHc25
cfwNsjXzwDTxnvpE3DXXj69ILeKdyvRCqHwxm/IAN3TgqmQ6+M/0DZ7BqoKbnK3amzus4igqxfMw
azNw2EGCFsqsR66lGKTcA5/szcmVBuwDEWG2UtxmPyDPEFOSfuk5bNqD6TnPzt00azC632ZT8VfB
U/yIECpVqtnW3eK13dxwYzm0OWs1Y6bNHbNOSmvQLh/XBnlk/CanS7SD1Uy7VAdwbZxDHB67qnFM
vQH53gzo3wHGLHFZ9bi76DUiVpQs9WJeU3gkZpvRjS61Y5yePDDYf1beyr5MttwHHGdoCxcBxoaR
RTe+6o7mn4+tA9Yvha6rFHAHFbjU31n8jADXRZlDes97jsarSOqC/WcHe7/DLT6zUFKDDRstnfo8
/k+j3vaf0kTszcSaldF9R3takwX4Jm7IUG/u2nJZzZhFhjpEQWbwpiNwr2McFfx+OfgTJ3Sf+O5f
jg62lRQYjk5c10KPZtFLrvII5J9k7hdcximzSgLdL6GMZ3GdywrDklVchh5t1epA5FBi/ouGwmlJ
Sc2jKOINNCtEQ7XUNJnV4pxjuYJXLEqakdGNXFBCTnbNyJLgumXoo4xhTbpGHnYKae/vVqMfFX5A
Fgrg4gcoZzf2M+01Y5+M3ZcqORKWGUg2McbLnZw5WeZISw7HQzzu27f518EhdvWtCmy5EZIbuCfG
Gwu5mjol+9rkzX4gj+XfBk5B8GUHZbjTvIfUZ7RO1e4pno5JAMSLKAfBuEa0JQWkp8F8bybQi67k
iFzUhfwnRzJDUtW0EBIYBZwaIyu1EXzGuzZGxSgPMWPXZx7pP+hoBMIxBVcluIpnyRNnT/krYbEN
jqZIaPMTOh+gGwGrX99rw5H6oSvBoOgBqRc8J107CS9F1UW68+Fe3q39E6n5JTz+yDCjlhbPWyaQ
JLEpwf5fYon68UCVZt5D3Y5nhDbnlSsbETLe7z5cMP9/KAMVS9IudjUOR93iPIfqnssaI+9zhc3N
JLdpnPQKGjR5stoLrBQcq4nl+Vkr0+Xc+vlcMk2WJbamN0s/ZTOpo675m/t+TcGOkjIi04MX7ZoP
ZXXzwo6VJnB8qfj3iD7R/66GtZH1pTK4OguaCZIZMqSegO4YCKmdbL9SE92dmzWMJghWD2oBvIhF
G7RbdzJFCjQWOQhF83iI4W9+4W4j8Wo83ylyjHzHzLLZVXWNEvGrAjo2eQea0ai6Fxa8PpqIEA2B
owCpK/ZxVUdos8UkLFNrVUqVuYYGZ5v9D4xUmo88OkPz3UvZTM6UFH/xYA+0XF3Jwp84+KNm2uDd
2PBOzZx5byi9eDQ4VZLejNP85ap0a1NBLjxfSePEulctyfa77TapQ8HuozgAlCNSQ3A1gF1pIxAx
ftiH3KlwReKIoiAwpv7goC2xb8Xj6R3vGslp/w1IQ54PNTEdbVzRjIpOEvEHV/yZcFEH/JmCMS9g
thBsEWFOTWyhheQ+52WOIhyoSxP5uRFEkr4KL92J5pOLCfRuLUqEQZVJRm8pgJR4X6z5M+VZtEWW
frbzg734JybOtQkAwC6c2S+bTACfuRMthuwkfjaOWN9LbTYCHVj22pKQ1HJP0MH4mHrrnI8CRRIO
vQ/o8rLG8cHWDXCYD/3FEDVpmJkcGyfxGOyVsZH4Msnyuan2wkzJWZ+NWDtFMpFDjUFyQqQyYX46
CDd1CxQdgnIIZI2GDnjWQoqEHkFUF6QtKmUxYz82HapeaF4l1GZKlBR+hqj+1DpBa1UeMO2uvtd3
899z9SFaCOw2HQO9Fda06KFNGygnxU0SUr5yb5TK00C6+1WYe7fdpyQUyFCPFxno9ur0Flev9LdA
SGzhye8GL4sgJg0hVYcbeMQqzj+AH2Y+a07RgK9MiPIiNfpvcVTlLLubHMtqTQbSBYCRsbAsjehJ
erWqtOS1kkMQ6x/LrxvVI8njxsQkPtNbLjgr+lNG6MfPWyOx9GUsLmkU3W12/vT32Qav9toe3lG1
v7WE/93GP/9WUGv1iAc4C7FZiRM/X8qd1/lWFoFYocEprLy2xk2F94broq0wc6DdzBBCvN7a/LTV
KrJygWAkmBOwObLhadGCvEephL67Qyfs+DxtmIFwEWBXjGuy/EsKE++ZV5yEg/6RxLjKp3A/VaDQ
l9jTvYAjGkY1YqgZ47OOmesYExA9G6f/JGyaTKCENGTtiZ/BzBldbQLlZGOXrLmcueZsrnOfamEH
Cwl4lTZIWVomuJ251swYuq3cFm35mlNgLbrXAimYvSyGduCIy5bo5MwecpFUY1JhEA+zLHXdkVj/
qbHvyANJI0xMU9yP4MSpRQtY5GNXdJKMNJxW2ht9atfMa8vMJkZbh/3kegioY/JEB7mYgsIpliK5
1K7rjL4VIHophM3YjSvxE0nXmhtUnp9TGKrMmqKeJBVuONN+bNksIj3c6XlGKTgbqvlYajXgBvM3
qD1wK5au+8curs9DCz1QEX5jAsCdrqX9doTVuCTbzbwYlPt4R9ghWh4SbcHtJ3yUEoHx5UM6yyAR
astXIY44tWrGcifXrxQLJrEj2g3lmaAMeTsWF7DvTxo6gzHkwC8kW3uvfZA1SU9hLfUBKn4jpe5w
v27G7eY3ucnI89SsKevYAyiEAugs2LlJX0PImmI2gk+Vqm6E5hpp5x1nwGPEce9ZEzIb8WzfvyDl
YwZPK7RJsTZef9Ml3jBZe0DvttzW1d87J9i7jB0WLNlChM2N+huS211urwUwCZhMdSgfnLJRqYMB
+dKah0XGswtjIxhZn3/r8aCfigWCndLDGocSktGCQU2UWC63DTBWfRH5XnccIv+gPn/ha/Xp22BZ
fIxgwTU4mmC7Y4Arcmo60X/T4zp/MybXkXkGnxH1uiewU1V/YigyCqGfB+MATighcGDtjSnTJAIN
4FELnZVQ380OMtE9YeBolzBpaJC4oSdzlPgyIH+Uus7IT/JQgBwHsHmUFHfMFsoEZftzdoNRQvaP
dCjXoT995iDO47cnVi/nZ8+C/FoHliyhW5dAPLtSIlieFjzbNDJC1lumc94je/MOPLgnYDYllrWK
k8QxOEZLFwlfIpcHPIjFVMDsAmo4cgpt2xGeY4mE/Fxtat8L/QWIIti5YZ2Sr9zrTih1dDu/0fYn
Kzp1Sw4nKXqHf1scNznJ2Y7qHAMYUDeoDZmOs24/mwAULGKxcbXWri+PVj95G7qGCfEpHFuCJJrd
CtYr+pbrDzJsUhmzOWlJbOfAPBzCPOubTTr0L/SLC20BwpDMhzzvaF9f37GCusyStN5BUC/aCRtl
MqRo8inWgNdAwcEtPGkxYhputspBdJck8bWN6MONeg4j3s9IbCotgggUAG8VPgaBq7gMdr4irr38
tQj5kU8TQLvQ7q9XYLSMF9lEl+Mr/IwpVXiwqOcWlR6RshnO3dqnBiJJ07L3Bv7wcuo+ObSEnYYc
q0Eoc6YTzuavIXboSMarRcWhqU9jS9lY7FYpHcmBIOZbw+8pqkenwSJpW5+lJ6uHlT15kXfC6BSA
t+yra0/WPrHg2vm+3B+O96nfJ5ZWRf7kvZGsV2f5cEp2TUtYj5AmtHsbWYyZMVgg1G5wtthIxzZP
066yaatf0eHhgIYVb2KBUnCBvscWwN36WgNKFTGTqWLQ9tVXQfs/nB6avXikHruSa0IsI7peQC7a
c7kuvuZw7z+EXPzE9SS61Per0/e2q/4p60ePcOZjP+1eM81Lt3IYnoV9BQgB0h3t677RRtuFPHlY
XRhk29iBixhQDn8uurpOsrgf37r5r/daAjH1B3vqt5GbZy3Vymy3hob5IjiODmnQWhGJzt0ZVioi
Hmf/Scx1XuIR/hdQF54G0DulDBLzN9tTDLkI4m9ra+SmcFtIxgRtoGmyz666JNbTHcXce54f38Xt
thTEuCa1OSJa60FO1hnJ8Ylm8j7peJrC/cMCVJ4vs5q96tZkAoxubXoDZlSe97HYAAzl0X/VpHdD
vXDzMmv1DaM/IOI2g7GyGDUaDAK90Ppt3+4zLTsqX2DUbmNGF0GPmkPEC+20Awukh/SrSK/loS9X
abE8K0K7UcwisuKNuXEsayxqF2ZrVzQ4TNdK/Hu7lbWp8arpFpdeKYzt68oxJdqXYCVJ+PgqPYUN
uUKhac9eSUmBPIbFCjVXH3IcS0JPCnkB2Y9lpB6MiuxVpfRfCeJTXyUNaVhl8OsBFhwqrpvrbgo3
vvMy5Ouy42/jiCEFiMol51lCCLLmU0SOJY6/yXclAWbEujMRYD2vePgFN1YjGvINd760dJibYH4v
kz4mx1VR86W4Te7Fyq0vB/7ytkNIzHLQuJ7jjRfdM6Q2BHFLiKER7yartQ+5mGBKz64JTLGqstxu
EFyGcsz2x3eDiA05JQOJjy0ZpyfpBPHRe6dKHINOHrr44flpFO7xqQGiS8hrZ+y53ApM0L/Mkoy5
78Cz2CHYwtrUfof6CtHWKFsJiria1GUu9C7PJRZyEYNwlukznv4w9YSxm9uO/j/MID60Z6hCg3tu
4LBM5yScYxKPTJF6QiMl+hnJXpeTOnkbet1+yEV4VBSxzOfTSbVLmh5GT0ef0E3aZE5vdsnydiue
QR229fip+r4Y/uDyAF1Klm5XfujDNM8w6DleffCugtKaN8BGLDrEeHwOErXbRGLxKnBtysHMCFZ9
JbbzkbtHh5Bblu/gvsZsEHymgAxU727lcGJ3PqebIBTNStp0Z/HxG4B1K1LMm3kcSiuX4om+LNLY
K5yviUnuAKbLMrvy0oDottr2vUVG8ZW7eEzzBpMgECmB1cr6VKjyl/HOUPrm2xP5BpPVsbur39Mv
FTTLi14zPkeH1U0mghnwHAvM1YhYCc7zbnv8w3r95JglGu5UCim4ru3Zv+VAXMT4OygKjKs4iMzo
ybdJqd+Kz/F2f/XxgOyMBJc7noNO2F56ya6U9AdJAd1pEWRsqiyovf3hGpx9GcQH0ZXZPy8TV8kF
P7qr2bePQj+VXwK+mpasrUwKr4pwV/4E31ZfQAZMjUTZOkbmeXHO5bcxVtQDhTVxCapL7jwLCdPO
sQiiBpjK3tivosq8WpfNnYWhHLzFLDZ58dSdQZE/l5y+CMKGz3ciAOOrIc/QWeWix7uQMfNQ2nVH
nukneTsRL7aYCWnF0SyrRTOONRQl9PqSOKWVBx7mln1HJMjoqE6fa6SwLh1aRTej7Z1QJNxNfVAT
lsfZfGttKOgv1srxaQ/GP/frg/XNB6N7qoUCQK3k5EIcByetOCJIiPZTpj6DW7u+TatD5C749aWx
dFS9mJ5aGFOR7IEoT5UlyQMr5cr4YdrXD6tivqbEIsaYtd1UuAXmf7uA2jy4tw1XnvPPd6zlDj8S
tPnHoFrVghQSg3f4PrMrfsKgYnz5BnIkxYLU1JTQ7+IbMLQRYQLJkRHoSspbXvWCOujroj1n8vzt
pS/+0CBOB6eqNTI7RxbQ4yklpx1Yx5MPhhy6U5jyQSiACxMYsC+ub910F6kNU/YOcYtSPsUiK4Jn
JU/LIFHS0oKf8wa18zh5VKPI7ECFA2SdAOPBAzOFnrn//5YYlUZJOcoonp1rZI7xK89A5Jsh3fPi
ZUXHIEYi3TSj2tsIbq8KHSo5ddxZNTWHaAZToV6x47xY2TFdKPZy4lx2ATh1XgqPm3/vF6naX2aG
XScuedOOZ+iuePDmcM/rIde0jESyvbBlQtx/DXsrtjHVdwy201DjfvZJp9jWcjViJjP57fqO5NEN
/9hgvwskyh4SLUvy+cCeKNEPpPoYH9fnuAZ1QpxAUWq/FFlAT4vh3aktCt5LQfZ2q9WBF880hjWK
6zX1i2mHCGD2Xl0ZHunTczyrsSbDcFPxPTVqj1CQhNJ4D0G6WESA391VCUUKl3K7tJvGDfbHvBWU
XrQk4AgFYGO7vH4htuc7gzXLQolgmYxP4S08T6/NME2vz2eh7xrLJ7WRyx8xV10of2FnqvEO2zMK
JSTVWn51epLTwx/1rpF0pPTFnfHxv4DQCgxppYj+u1L2APSv3+g5YUD4NsJMQDH+Wpf0lb1vIvNX
WxvuzLP4FITJtF37O4ZQOH2/gmNYTFRlwch7lcEPwvwD/djWLtUYHhb7XhE4JQ6EqwX9E4OV01Pz
VtmMomfYilBlTKZYyIa6ZmW0s6I3Qcn8teNyg6JVnCABwIL4PfShIfLDoKO96yp8WGNf83MPQCZu
aE+8WCHOawTdaUOZEw+yxJ+7oq1knNT3V7atStiBSwiGbLAe9AkQWVaieIuJfQ8ShJwMN/eet2I/
JLsd65uqQFW4+PrtOwWFe3epfzDIm27gpi7lDYXUK2seV6kwGGuSAuC0d5IMFeO8V4NkMO7vyYY2
WCDkbj1gqmBIkmlv+VAad94sFxWIIcypWEe9wmNr4p/KphJ5/PaHZQS2xa6yn6NIV6NppFwD7vKJ
+7l1MOhj0Mm244vhcSg+36KTUFyiGhk3CBWCKe+PvJYnsjXP/9h4+v7JsdW/HGCtK68UmQgijRkM
RcDGs/vNVyS9kSYZ0KNbtljNf8kXJBSpYsGD/mbfZOIw/YRSIcnDo88lFPHGROyBwNGDzbNGeAon
jBFS2Kv4hMtGpi003AZlXyr5GXus/DasiBsu9tUf+tdONH7z4aqUuljqVerGWNAZZ9z9O0W5MrbU
x6ULOGQnehI0Ae68D7c7+qrclFN557om2EmPE5XlkY8bqbm6nuozovGPS0lOvzpG5zXsG/6opbQf
wrQY3yDxFvameYfDNbqAAOZdUgCL70faWR1bU4PyzwS1tnvics6mRdc9nVRpb0wH/1LpWDtPt1pc
xBzgqGEwiz+wqpdYf1JUiREY+EcEPC+aROmQZnjrdiIFjKCte9bQ5ZAerHQJQ2OzRao0FJOYuLRQ
2pOSzZ4jv1dbnfvV675fKXBjA9V0kMYqnARYgEdL4p+82ZYoV0X9M6e3uvfdrUFA6gaEvuyjCEum
FpkfBRa0po3+s2DmIVAikAlK7UoFaBdng+hzJBqRjuafBAeZOl+3DQJrx/CCoGkT/5RW2PY3QZqk
Em9p8jcl3tqjhM1aUWqeiB75KENE26QNN161ZddSIFpZswDj/jO+DG//88K33ckQKVF0SWjR4YC5
27Gbrnx4dzTgGDeOFaYyhKhb1OcNVSaz4pk6QcDDfiaxWsbdqZ75iEUeE5h2ULHsGGYp4GMyfYdP
EKBr0ChVSbX2AVY36g7uVUVKQ2TvVymmbAdUBYPIk65O4IFpYRxVGNlDT82sFhJnXMm94Sw49k8E
KzItCW9XPPJKn8Jcj/zcQJuV419DyzdB1YnUA6dka0nHU0/sh4UinZAO4izQKmD96+0WHFn6v02G
7gSniPi880FjO5J7N4fIE68RxTM0vQ8vIx1Oq0n/V6vMJE6fq+hJZ1H23zwCdZQ3kKvNkc2rKILO
4tqF8tHXnaDhT9vN0ELuepfA4A9hVVRzvfZxViLsfHGyKo7soRAF59QRovnxYH99ojBR7ZM8zd4W
zJ5qQHsN0drnkP6wYVtjBXnHMjKEdBmDocHyOztZnN7pJOHUIQyUUe+KiiZzCdAC3KQm5THc3ROK
kSLv1ZFb7w+mmoU0n+H84IYsFHsF/FH8zOCHKqLYt0zWqp1hud8VJaZL3/T/P+W8MVYE+8+hEMJC
cXlqj90C+/5Ca4yfmP392aBhgY/gGILKu2H4cTbGwnnv9SJCJ743SJQng9XXm3lci6yynIGqr1fI
Gd6BazsrXMT/YavVooiCmDyQnK7EGc8xrvD00CCWyRAlWNS4sUN41RmHhKKPbEMQuyi781HOc73N
PY5RMDVsNpKORCq2SRZHfI5TWS9by34ijKU1e+x7K2qHaACDr49mQi9L1g3CZm4LHVG82iTx6/Ja
W1dnIL44WLOo7C9r2q6581EQ4s9wqvtZer4lecEvYr+ao8wvHP6F6N3dEb8NdsZ54BV0UbDtvO5E
f94EWdCvHHjkX6J3XScCtfopiW6972j55CvL6+zGdkKW2vo8lXYZT7m4JVSlsPd49JiAE8lS282/
TD7jRKZEkT84KUSPVaVmedOYMsW5QZ0JWKLB8eYPV5Pt3hsctDDcjOhvWpcTlqUHxsshXBpM17mx
9/U+qhqUb+/9AKIJh41Ykhj1SDJRqoewOajUZFEBZ+x619TPNGg8cqwIfq0SsbLF8L8t8DaVUPHm
3olrxvJBt7w+srNkN9tP1P2brxvBmz0AoeX5y+3nWIEhj7dAXXFQF5rfTjk/VTlYwnPOQTeD1SwM
aHSsP+ROeCwwa7kWnpwqKCNQgQqi1rFYSiBt7p9GZof9HQhRIR+3c1+rgrqu3rSd8dNOCMTet9YK
nNWqWwQbXAUx6Ok0boBeDeOl1WG/5HMjF8dUuy6gx9AShHwAq+aovUqOEbotfx86UgJo4QBnS+qq
cPdEPf7alPr9mRGPbzh9pVMDQfUOx6qiXDKreIkVII90jezPt+23GCSowTtFpsiMEtUgkf/gK5Id
S8REx6s9to5+lvnskv8hYoMoWGrrn5AVFppiOb1TAzKN+faBcUNzzooc6XW5QJHk4tZyGaRprrHN
elgJnPYIejV7Sf3PekZ3I7RSMnSLwIoXJJjzbxY6GC+tkieJX095CtU+PWwHkD2SsaJAcq7sQs5k
s5GYUUWdWvv1WlKP8kCvrwvcA3jTk8Li7SaunD/WpAynqEAoeYZdhiClA6rpkAapxCdLMA3ca5jV
OvHE4EI+alIUKwsAYxytYehcJP80TwpTLe7nslcfw2FU6kffBjQX3dLkEU3bHsOtlKRAt7Zj4uoz
6E3tRDsY3MXrOlYN2JesUa4CPc4C4plvqh3hUZHIT5GyocQBhIls+tlL5gnJ3UbuDFHMj6X/PR9H
juhqMtJT9DPoTRZzvb4i4QlRJXX/GHMD72Cjw1xUgy5hDSe2hUuyY1Q9peXGM20M4kQ+IjGUcPh8
xzAFscnh75X0MxV3o8HA/tX3onORfBy2FVSRe4rGxzCNCLRA16MOedmxnS/b8Qs7EoGAUkSUDTdj
y+in6Xj8oSK1/ic1WrSzoRshkNqqFSCffO21wKGZYMfwWolvA66TrZciVFHUvr6nAkZI7Mkfr7Hf
cz4PrwlMf+kOdfANDtaGrxqOlbkwtNj3HLuaEYOBiTH59njBV2QktXB6QVkhj7ChrPE6+VhzOZbK
KedAkVQluo57ZUKZG8J975bw+cvDEY0MpbroqBwR/dtdGD3uJuKWt/FZV5a/jfQ9XjdZrNw/bZL5
o9YOstZp8zHgx0siGNbzVyBPJ3hUpXgXvLPqe9GxCn3TLIV/zgJdyTPgmJbZbKvdGpj14121azRP
kkARO8MCDAEfF3c7xRFDM9rQD/hUd8WfvP7DdX3YA275ffd/OaqB+wayl766WL6FFVTMRlffoBbF
aSfgR8ce+fEgpXljSY/fVmmDY9joA2JCjnmUb1ZSlkqpxm9QzN3mmG3FSS8nNce7c9qF/avdFA7T
bytumGMbVo4Y5E+ZZkqbcZQBBglNZCq6cUFeYLm4wUo+B3zSO6+PmUlliIEZNz5WJlwBwVYePmwo
WufiBHQxCatMi3jik4h8ljE08DiHz2GtGURPtkJmTxD+8zzNL793yUKRn1LDVpmnTEqqbnzYV50b
rFZoUnyvp0V79/eJ+Hv+lMCwTk5TVomoeDAQEtT/i7pURcUHaAYf+ebrtbnW5qzzTL1ftp69BmWN
FRqOWfWBx9zOdp82uQYnWA0Wl+UQOO+PwhK2Lkm16LU+O0bcKztYLIuPFrcRzvfmIL5DBejeDl3z
SESqZ3coaEpMdZkNlLruG1Njl6phhJ0iOMd1Dmt9jKw5m/JJOGSwVPsnXjro2FJ/0JXYkdEpnECI
bow1mDd2eTWULsArFWtr+YdnbjZ1atx2Ea2LsLXDqwTYzp/mkb40nS7RG4pNzGbL17aud1pxxuLq
vdxioVfZhFf8WLiaQ3J9vhF3MJ9Qkeglzx2ucgl5Zo6ewKZT98i6ImvhYWeQbR2IxdOATZYc90C6
PPFTArXHCGcbdkKE4dk9bqSXJxxkzjsI8OeZ6ls9XAOH2cElZ7AgkCNYp6EWu/AmDreSWCiftIYD
1keXIl4IWJSSjk9/pYtB3ozVLH7g9KWD4wQJFDyH1DyHOELBEs2nnlDNU3fEwV0HZ6sxtpdOMkNk
p5qNE7DemTvxMvi/nTDqodj4GZo0x0U3IXvFRoPzHgpkPAJfblXQYGCzusl2+75DwvQmTYzyz1+9
cih5BkwGj6F4pbKsCGa1hUMCtDyS1foQaJO8s+O+AdCDzZBOHeEdd+hhfE0bOcu3uLnhUO1lh/uz
SofNOjwB6WqKzf1rjQJm6iuaYZKKVfIRcFEB3Qafh5n/YkvKzgHAH9CLfqH5vRijxCiirMg3Hwov
7TYRLx9iKM3BRyhncCwCKvpBRmPIrpDP5ixku7MVM315KldWj7txghdOcXKrndUkLkcxmcG7V6B6
Y2FKnFZbenZwtokJJOb6jqFs+PIMsEWg1l+qXjqk499lhoZxd9QR5OVtzh+mPQgZeyZLiIbQdk5M
TrGp7WdZYq7gFumi5TilUzcU+NQBrNlSKukBrboSLilV+guWYsOOk6wRYtk/vR9Zs6IZyQKhFtv5
tVGzYjUNUMJMtUjFDOmBI8uAPeuydgWyCEguyWMjnX/piLQODZC6elu/E33Q4YZ6AN+9cUzJRwvB
S22vnGDPy0StjygHDVPP5n73vDwAXBxJw8AHJV1zaG+IbrdUpBaglUD0P86HTkoi8I4iClLK5Y64
hrtPw9imHZb1HaO2p/rsfWSYuDeegcl8Heq7AQLnmz8U/lluk8Ltn3eB3M07coTwmI01C8UEtjUr
14ScBo/i7OoVPnx6q97FFysZdiKDnOnrhdqC4ire+M69WXWWXV/o/8RW/pxvS2L++uhZ1TrxHj8c
lIoT3epBeIgHkWSLllwMGAfBAmuwN89iR9iMx6iCJOpByngJom5LR4Aixjr+gq9+jqzDieJa2sZX
2IsDvXBUljR3LIF76yJMDd8NDTyi/1hSc6g/GnURX14RTvik0OEsbEljpBbAVvAvrTYmacEIvHGm
sEDQC9mUFIEGhnb/IVPSdZZv3uhuKl0so8bOmfjkMpaI0bNN3w6xNAmRXUOpfSbsRbLzBM281nf3
DjQ+aM+foJJs/oyWgcIiAanlQw2AyQN8wQgpUHKh/ZjcrjZ89IiHNkP+l4BEBXlVBa8dVznim7T3
Tb5vxawEdxp7aJyMZMVpyu+5JNcsaFnqlxxfF7CzfE7iEFa750nv1G+BPvNfgOEBMppo2gPIQwMn
4pil0CWOv4fXK0g2CYuMoYDr5/3tmCrHOhV6hZtqUxsYcb8Nu2j6PhFcAizAS5s6jQxQBeCOHlhi
F9o4drcfRZKtLxhFFkzfk6NH/+ifJy167H17icQpqOh88rPBEAnbMQgrpeUuPAiYrBNb47tl25Bw
oNaLISqMSUdHsf/oAKuvKP5quejvyiLZzQL7K6xatdt4Gv3VM6wYe4opDF6EdYgCFHXIyaA0kSOL
k6sdjUR0c5ac+8bH5rDxklB98WXlT+x93JUye222yDX3ranTPl1G9QavehCQndeEtbOjmiJTdQZs
ZkFYSdUylUSpkPl4YDYMy2/i3iYYqnkIUAsLImx04IFwRssI5PAPXnZSgKhbvWDmZ97HdjE1n/ZO
yjagfH0Y0xIhdcNZnMk1+d8QjU1ICqsoa68+mwEbeviT/8l3Q5++FGgVyD9jk9KfPlnzqrjRKker
WfRDH+c94Skg3q6I5hcXKnkzm9XH48r0gEtzGlljY0CMoO8ON/2OKvM87iaf7bYs1A+5ZB33GTnL
CKas6F4atNp6JJEQYA+BHNNzmwNANk12UOyJbw9DnJVGxDhputw4Je/rv6l/o2f1BaFp0WK9FYE9
1z85qx++28+WdoMb7mnz6cIqv1wkoQKX5KJ1RhN5ZRz8M8dT83+THS18/ALdRD3YbGmbA06BkTcx
hxBHMOEmxDMk+JTQ7Xh36c/DBHw6KwUqygurHP5Ki8tEuQWCiwbTAj/bvXvJaCNveC++uhZsoNsl
z4557x8DMizhsv1WTSFB8LqWUhPTCgG8WxLpKrkx9UIPYWWbMdViHxvvZ0LMuj9Q5tYLD5ezINkI
+Uf7/yk9oM8/LVTNi7wG3aAHEGR/LguLAweTtsxiqgH9t+vq0avGhpCHsNdTrVvT/RYx9yxyTYDi
VlytKyQ253UYTlR0/EXvrjcUubCVSlkHNHo9hu4Oq+PNfs/cV2a3xldVKy3cP8P3ANDgVpLmdfTR
qQQNjhMzIW0Q22qMTn6jM4GCcKdPL4OdhV1j//QNdkwOaoHVDh8/CyyO1iitKQFAC6yrA3iFt/2i
sKM/gHgmiBFtkQAxFuo2AA2jUweXOPhvNG5xgVqe3JWiAksowgHUPAIbjUvtYV8csuHGJLcf0MTD
O67Lb+WvwCO8+VmH/rouRPrDZZZemUe2Wundv+CD4n9yoeVyJS/BE0uCNxA2ghryhpoBphHdQUKy
7q+HwSnsh9LPhsdM6eTv8rtRx7qmNXm7QbvfKNvDzqiwMWJfwbP/ocqdf6hQ7cICQmvcdCtCeKNG
vxnJP8huFg0jnXQuA/ueX+zIyPwNSgSe8shbW5/fcPctWwxHBs4h4jMWAkqFc3RyCstckHqxjTET
LQHtFHy0t7+72S1ri43TVjv96vkIsmohs8D3ZszLLDoDT1sr7ixnJ+gbed5QToVhDd3/Hp+5pkDB
n5uliazQl1MYdQOqgnFC/j91MGt2GbZ10yQh5qVc3cGc0wOIiUw7B/gQfCzterqs8JwlTNgyBY8v
7VodAO4kYd8yBRuIg8B1EqsaZYc10r8x4UiDRtZztoBUeGmzwCAyDFzTvT+to6NHEdUgg2wovcD6
ihEBrzl7vgNSUW2oSrSgqBZvdY5ZuGPaJOU7jXwUKdQdMxAt5hxP1U2uNlMS3GioKtBl8KJyC8AW
483l1NmMQwMndRrHwA7pMiUOT4o+fX5Q7ky6mqSerpWCsMTC5BI6sDj29lxDGwQv48NJTcoIVS9K
/72n4Ue6TY2HzgYrQQv+0LLkXbNk0xl0zFDKqAo9Vjq0Fsa+LHn03y4iRuKZKYlHsH/ig6mC2/ni
H/u8yJEQQFQ1HOtfkzsUlVwfybVX4UoZ/SmSwjI3EtaDprUgEeUrljPCaey5Y9rwLH5m5kS+imMe
iiwcICCAG1gGFvpELm1NCxu4osMv21IIB8+HqtQGWyvq2e3OJ0zbr0GMTOycrrNtSXTKmpKV50Rv
ULqPcK57PTXWL0p8yX52ZGHlynNclLXi9dt+uD9ZSjKyB4RLkNEarhnxGThcw62cr7mDmsvtQo3Y
j+uZuQayzsAqONxi1qNd24x8kgIgjVahbWGYEA7YQGpEYlvAcjVusAZceJmu1FokueLnWfBzJPer
2bij2B4R7aOF/hrF8fjpgiYf/xP93NEsdjiIhn+Ptfl2iGvp12RpdVkWIiGaRuWQX926IQncGejT
7jGCUdsOvDSf78TY7M7au9yuMFfoZhDjRRQVw0tUfvpnmzR3weSeEneKld8SNBMFe/Nx67n/EGGN
mrEMgJjWOxiPD4XO8Bq1LWi14+VwDeb0MSkgGARCPvW+Fq5reN/KycUSGH78OO6gH87y5xf9BT82
bs1BredbMaOkDZKDMaCz+/dfLGetgKGIyzv5p0gOdksGCbqCqzzvfxGmoqMgki+p9GgM8Ufo4ZQf
5fS1szKza+9hUDBqXl+A0lSshtwZ+idWKbrR4pV1Ae7efY7Nwy2BM3R4KNeYTSznSsjo820UG4wF
rNesAJUBybhCaSzTqujb6cU6t4jzAHbDrm0WA/Dp4q37JQ3gOaDkMioFfyY2Qv0JjECXy1kSt9ex
7N+g06YBn+W7dA7clkepKb5LsH1IqBNVvBqT7K+qB3HIJUxpqm6JXKNX3ugQqi2ECV9v6aT0jmzj
vgnDtb3Qa4KMZOLnVJPeqAm5jpaCgzwpKLsu6qjO71UTcqaTGn8l1hn4Lx0AEyQ3PSWvvVmyyhxj
PwgSCNYez/B2aSo7zaXr25lGoF8XMO14wCViUAIN5o5M6db+0tM2y0gHZ/3NOu9rk8VHSdZ+S8Lw
4Fm0rJfCG0mG9ah3t23PPDYW3/pzkGPEGXh6hLcHoNGuWVjMwCfWmYd85DjYblqO2ewLcfXrqG9V
1vXg/oykhGy80bGtw5kRqry4AbKI24D5mJ8rF8JZbsAD/+cxcgQkh3Jap+LhqTBsMdSIpGWCHbEW
OQKYbeRgIsFBh3WiXD+dQTgC7UKfObHK8Npr2RsFUbqr4lb3fQ3zhWhLA6iBgBsd4PWAYngjtfqW
J61XghXnJGGfqu84YkLQknt7iVaPXrLeLGyOjEzryOvL2O/lsdp3mnH0MZGCogm8JCqckjnOEIVG
xeWoJWYrPy7ux0M8GDf9BPxQZfIxZ3XreACYxh9dp+DeK3dSb+a7xuVOgsA7f6EVBnjte/KGhDUy
StUTMfhWZlqCm6IpZLvak77XomjiNBU+idDPHyCZNgeVfMaXonC/s5JShrlOWKy8Y0WxXjSqoT7j
s8JpF92OZ2aACNBi9B+f72FkhixZ2voXv6sF4jbxIYPqg5lzT/98bdpROA2jIKxgJt77d4YQym1c
oKxzzt7GlUgZQGFN/P4j8GQskrd0CyJ5l4qzBP4kwqA2s8NrZrtajnuptcLxuoh5OeXhiIX6lM44
N5xX2wlb73MHogBr14patgz53KqciCGeeCauS9aYl95LUQ0s6se0Y6tKBs1JN/a7mKhZnrS6914f
qvk9IbYtxXQNo5CJyV5tAGt0z7P6duPSoBHJeZ7bYMcinuLH838R+xGYOjy2pBPY0gnC7gMUu4aM
/MO/5d3CyBAp0Ve/KUT+XdR5GraoKSM01FFL5M/TZWy0WaOYLwjrI9jJREGqaDXo9Kgw+Yb+4PTC
SJYgBm8ZyRuX+lrd1d74qqaQyhjgJuAfwzS1tdxvdjq8Lx5F6qMjuuVKDzUPuG5g2C0HcJ1c6OLC
h7v4PCUeTnOA/lHcvif42mGr/bmwUC2UcaFnxRzGIPGycaiE6gQMMWpAX5+LDqKQTBSp0bSH9ieS
8qTK9iqzKGMPVSTy32RoCghc6pCkmgGzy4NSglP8dlKKVEHPoBbXySm8cXFJJmLs4sV4cv9SDYXN
uvd1QC3oL5DOVu0GMCrhnMSvRKJ4xYRIpWjTBPVCmtdk7j9VqxpPu3/OCFffWiYW8hMKhTqU0mfc
6PniIC2fYrKh8AiSwMjIL6tnk9HdIqkroXV/U7p5owyF4LBHtCy41Y+rvZvd7TCf1Q+gNW7RILvb
uZKmpwDI7U+0ZH6QbSfE5aoxNCIsTNm7Yly25HVrkSCtXZxmsa7OnAKUeqEK5bpl9CQFizRtRNjJ
d68jK9W0mKYheIv9UiZmAFnvNRm6kawLkFtFF0VeG8KAP+VpE2QN4K2kh8ZrcQB9cZla8zcdm18B
d98kvhXinqVEHsSiNgSEn+7KRpwzt0Ng+65rPltsWNq6Fkn4dXnX2Y6kLlomb2joo4BpIJtJYtS+
QFJ0dREayfCt4VADvqARGVIeUtY5DEbNFS3mq7kV00j6RmCnl0Tw9HD0GbBpw5KRHvWwbML3ZaHo
fn20Wqm2BrImlYgKt7lsiv5K/9Jz50EGN8UnRKzJ6y5mAgHTkp4YH1rCqBpre3r6qQyQuDbaEfe3
0VrhjoMBRhik4MS1W6IOa/Mxl98oW7H5mV92w/gVRo43YgbjHJntDL10w4BmpwVHqGt8e5VbFaTv
TeTgXyC57kvd5KvEqgcQFAU7z9FN0C6I7e2hwmXuQv4wsBrbl4wFHX/fPSzM6WPX188/8DXOIP77
UVarZlGr6gxF/p4KUFQON2PjUhi0xWmwLXxllz/hk+QmCsY1Vy4KMPlQJKaIWulOY/f80Uky/ogV
Qq6Q0DibaBXy9o21lUqkBpUF7zgr5aKotTCmOVTPlAdumbUpqp5clCynQSYyjo04BD29nfmGoPAU
+AzAePq6HTyW4GuvAPhr5L0p7FBuXnf5fX2J2AOgbteSt4VHJDivzwsbPphUMB450lcx5v5ELJ+h
oFGhoOwjqlUseai520KSjNDwnwN0PD4q8AvBPBhAeOdOIXVoV+H1jYskBKAk87u7p4zr8MmU1SKU
7DCk2gmL34yhlZ4q470zEg90KrsiAjymuyOr5MYuskP2V2RzYCkajtkIlALRk7K+kRazWLkygp+Q
DZqN9rTt7sgo7NvUjWmp6B1BDdgeeLvl3npcjIEZUlXlxgnBf2WfCgF2fAdyFCu1czyY/2WStV03
wmANIDjc4FAL6t4hSAzubUDEHK7VKCC8AlEIysRhzd4AeQneKRxRJ1aZRaHHucGlXkCM9QuNP66F
sCFPEbQ9qXqWhEkEUCCA1+bxLpNEZOAWgDOGN1749s5VyWkxYExpL5JX6CKaCh7N0GcDOkr32Faz
iv/9/REEIpJ9rjKbLTjGqoSUpXvnw0tNutkT4hmxSfOmTevBr3VFjd1iCEsu3uL106DVJ9V4VHcx
rghZk+T1T/vUwXcz86df6pbk2UBxFPD0fs3SHXHJSSxzZPsSWKyP2SUurSdsqpXJ2XLvcXFCChCQ
15Lw4pYLOWizqrDKAFyUuk0wg7WEIe0AxCvK8RaxM4opkspHhXOxxU/p855GJlFbrJRLbsljHTDb
38QOyLIJkthLsn2aP16XTq4udQLhwUb6M00q2xsgjODurAzvokBC+yEVvhQD25FLtAWeXB0iWvoG
YogJVEHcfAt1KO3Aw522hn4TAzCoz9wibqzk4bIsORmqr3nZfsDJiWcveoDmhern2RXtxSXAnnzA
aBcX/1lyWfKc3q3jpgtVoUZtmwoGpOiWrxZ34gWxieoCUvlt0F/BC1N1cjxcd76UneREDNhUmZ4B
6AViJMNOj1ZDrhzmghsRKCd5CqNYRbIMo8F+oKjBUpwqmSf9nI4W7rhMHbBvOdmDEgkp526iU6KZ
TfladmZyKIbrox54LOajajvGEUAuEPx8cADSL4FN4Shg8dhEjtMoZBptvfo1ozY/I3/RXUZO8wsv
UvihlvPU1DEiU3psZNsHJkiVMR37gsvbH7NQPSCqEvfEvkWtjo1EkqkhgutFIFeMjeFqAHt43btQ
aijzO7fgsuiklwnyiHTuPn8xC5dsTgc9e+wNj6IkS3MrIZb0X3XLzxP53QyJqVW7l57/sWmD6HQu
z7o0lIRhSc6eHTnMkpgMb4Npm6gjZmUut04SxumwU4txRUH7V6YALTB4KlAVtVrbTyEePnLTTWTK
oymIpXAs8+JTOkCAJjWLubOYUwn5F6RsO4DM0VmJeMzCLP3stfoPHtV8wSTM+ezErYUHkPpUnXtI
xaPWVP/w581FRGpqkyQ2NVteo4vx/dhfFCkagiEeMRQdVbYqftblnv3TmyX63ErNZLuB5F+zPrA/
VvbduwcgfGvZtk67AXhWAyXHCEqPp/p0u9XStbeZfmLt7LWgws30C1WUxmLEOsAXz6e/tblD+zFQ
nGSVD8z6WRIhyK7r9XBDZKhacT9cFqTsbtBGw9CJstCz9BKyUoeZ0/bjxo8NMnXLyxTzMUg8Gqim
jKay1gC1687k3oiA5skLH9GgQrkcv9iWFrKpc53z6Xr2b7xBJrUXYQ3YAs96HP8Ay0CT3IiFT7Mz
sS2s6vW7uc1J7Iht8fmu5ozPNe/qBCq47q5x6CnyRU+q9lZmG40d99jOCk+DQtjPl/K5HvjG7GBH
BoGYScowwczlatRcZAa7iy9BjoVHTTDbfdaKuY9UUmhNJjMc6i8XyKYB5Xx4ukxXgcUnrU7Xg+Xn
TY4WOwssKQCTEXXJSnpJxxsufGYe1SBc3ettNtVepcVrIfG8ofGcQcKWD9AuneooF1s7nRuu/Fw4
/mdebz2lTrwN5K0QM9BnE5/xun11JTmbxmzilDpn8j2NuA8Qi96w72DVvKQLShSUhQtLIgHk+OKo
SD26G+bliYSVUbqynIUQlXaS9drYKzPglPoCdW95vJFP1rtQ7bN+8hwWeIOYBBQoQ4S3Qwq2uim6
VBz/JGeMm9k3qfCmbYcipNSnFKUHmOqU4QfHNjY9uI8dQUJg5IqdZa1C0LgjQlNqRqrn4DX/t1SC
1dtdYqdUG/8AiOFtmLLVHdhbGv9zvrrb0PUU1Ubo7ul8OOIOd330CGOw0tRCPkH0CQ+YzqzNH5jy
c3MOGaSLt6Saz3RQZuFnAnKHoynllXAp3g7+fDYyGBd3A1AVFnIBjq2zl8CpmfcUhdMYfc4psfaD
Mkuq9/SgR74uIv89Pk6zktNAVCKEBkOzLPJEGeMyGd/z502ZbIy08jKRRLSrhBgmHcwNWHHKtZYT
TuW5mIhUAosMCR2Z0J23O5vB4gAjRzUMbYK8RP+ZiQemJzZUktK8fB+ZYSAoSOCRlx7z3p9LWNTU
vyYYfTr6/lAC26zCeE0MBlL5ZGkovNKpZMCaxPquxBTiLrumEOYIYwX2fe4T7vYipUm42MeSG0V0
gbTbD3al4HVRv51RTzVW2RKGgsi+FjDNceAdHMdMR+P6CktMrB37O7DAvhhQRIcUyY2r7rqj0UC4
tPSl3fXo+RvaMBNE7Q==
`protect end_protected

