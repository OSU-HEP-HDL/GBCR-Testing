

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oYYUZ0MeKqJUJoI7DJiuvSB+q5Ix+Iwj9N3EwG3d9aznfrZuw1+Fc2PVy4cVNiksbh9EhD023m7N
/1rZI7UBsA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BmgMGlUziZwp4Aeom40PM0gFb+Lk4HIg7NJ8Ke6/iR/nzJgqwxvBOYZHlsOO/Hp8XOgAeNb9Zd4o
mPFcvStSgKrLqxBJrTC4jOtTOOUVOGECik9X7RElVDiKeZuCTuuYfKks1rnTANMNKsXOPeJj6Svr
YyXA9D2NRP6YkUNuPRY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1jtnTjcMZBAylJ3gewlkrSdkM4rrC/SF7w+2Gpl8C9SK/D8Tzq+D0qrZVMnmX2MWMKbqqYu6bkIj
sy7Xox+kttnLUyhBRsrBNs6gr3T0xsxsJ7Gnyco/P3Bde80gstdJ+PNfjg9uJOXa0R4ym9WtfNGf
swawtPDRNO3XB4oPqX/YBORxc12Z2+Xzlc5kJQDf1WM1UoKUm0j7+JBzjmig2WrmokL853BM29jT
4Ht91JL1B2bOy9A+fEpZnVLxL5NzuQ9svrSJluHfL94vaMxePXlPq6InH4B+XQp0TAFlIitjElNz
4mBAF7U6zb9GPz8ite7f9+Ofg2sCbTc7qhRaHA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gQeqr96ZiBT2MmGHCpbhB9Ma/ONapmaS0FJH16GFlg7E/VRDUjqbqiiC9oovpVsOBnNDQZNmXNgv
dI/YoLxA/mPd3NXizDTj33SvvwJdHC+sPFJrC6pT5rNUHqY3WkLW4EktYj3xtwACazlM0R3H+N1W
ZL2jtTv4hCIZZw83DISHIwGMevxP0unAXWFpAlJTyOmzC5wsjnlwvjA6I18++KC1ECVIFCC+grSL
XEAA1xdZCU131f12m2UaGi1yGaQH3scoEe37TXsoGUkWCMAn3jD7PddNt1X5zhoSRxPsOfUDmtSO
kCNVtrnPznMY8kVS/SdMToJlnwH2sKbHJZ6YoQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aYbz66wynlNa4RYsWnE11uoqAUkMOGD1rK3oC0qHnHAmOdMhPdz4cV/CAQENwbN3ryQY7/k4qEBR
2l3bOqYxA0+CBRl+jt8CXXxWU8WE2qwf32lPVes4/pVAbKANmE02/Ysj4IR7MGLvUvtr934XOsBK
cCc/KqvEbWgnnzkEdl16nzyz9Je6iY7Ni836+/z9BA/OYPszoNI5lKgO/06ni9esrcL9aCuvKXjM
Vplsu70i86fjOGURYjM2YFmCk8Xng1M6ROF+0KD+TufNMvK1W5if6MPJr/BsB83OF/hzcDKyULpB
p2+Eliq8StuhC0n7jUXEo6ZGATEY2a8DWEYVhQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B8e2xR5DNyjb6SEEOPCOnfB9/yUC8O8izWpzVz5s4/hfcHkvr1SHS13gqMQDj1DN3uSpaoGxcSIv
a3uLHDL4nIDztAAEPOvl5rp/eCLKhGUauWJKGzgIaInIPCBXw0hsptiyzlIicQEO3rsxoS+LR4e9
ltN4asLfvR5i5+Aru5E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o08P3wLx4KXr1Q02DiaLH2vPxf0H1jXIwF3rbwsiMxYgYGWIJGF4/mxUFC7J/WeIjcsQFoTUns3o
ZlNZWWRR36HJ1r2GmZoMunV8HAWjNjCUrk6RBWvB/4dYllizQVzRhb+3YUjmiSEMr4rkGsWsR9/t
W+i6luLQskwMDbMnn7puINFUehSDaOzDytgvFigNs9cj7haJi7XjPeMPUBa/JbbTJGFnxz8xzl03
55+BSHF5m9JHUn2eN7uDkExSgYolpcYI1EQnoCH8U6Zfcweg7A+n5SfklkTKUeWInYHoz9tHbIHA
y9aJwNoT7f6uxEt4GVf7oKjEfFlxUe/yajXHuw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132672)
`protect data_block
ooDQOnVmP1FtSEjJMBtrfhRlRL1MIXfeZ8qojblwwgfZUEndvH0EAk8QQH9+gc1CXq3N2H/OgoFs
hQKTuMle9WxO7HibFyU9sVIhrhEhe3w8lVavg/lFgNL+NSJeuFeo0TU6mDGLh+F4a0MNQz/jksFy
zXEphyI2ERz2At09PDLFdFgbdXG2xv8FDISH9mrwtR8EuUr9OwrmF8VI0OhIx2TAObiZ2hRUaNri
aVTcb5zH7yVNr/JOqpSo/SAA2Cnk9Xm1MolIjbRAHX5aeDZxNATd6GiGnFzn+UrUVz8QozaMrdP/
Es3NW39s0q3iir5JH+zSJJ6MMZPsyYENcxIhFcNT06iZbhlWL90t9/FC3rlH86GrBfbpxVTm03C+
oFS4r3swk3enGT/6Hu3e0oYkKUWgEr6XCi0Fp4rCcVU65odCDpy/FZiw3ndIuK716Iidjy6Kvy56
yKhIcQqMxG3Qr3ARgLQIvj5gByojEoB2xbhvxlOWBIwish1UjLfnn9CYmOy6q0Nb5/CqOchUO+iy
JfvJcd1nPURMz+SwUad7GAmMp1Gueckx/nopDm7vxmxfQLsVB6BrvlV8whzkBBJDP0Mn+oMMIwtp
b7PKx+DVYqrcOI+p3/3L53dKilb1P55Ydp47WE54ELfAK9JNC7Z5Js+Jawo9ZTGd2fh66BlAL1sj
pRTUSQHA3BMaC67XAILjyxd/SzPvZlWy9Eka1VDmJ0oF12/7awM1yBtKaypwClerjv1rHABo7XGg
saSflqQIA/EnA5zsun1UVECKkXm6AGMHvQOVLK/3pkia4yYNSKqv/xaX3egEDlJcSr94qfwk3Wz1
cQu9CqJbPaKX2MB14fs6xZK61lkkZVIQc+Q8nr2fBWkhE7fSOk5vtgWZlAKV2PLk5iA5jPgfQvwc
idHZr9BH9iAn14+OMykSL8QVqYLYcicTNnUwJvF375fcGXd/EgnZYVAN0HP0vGVPrealUijZp65S
cT9wqNjtNJtZ4OpoZUNqoQux6IHg75Mh1VD8BIUCmLe7T9pyEu0pcLFMR0i9g2h4PTyIRBlOydtn
O5UNpUm0tQeI9mXa09aoWdjCg90FjiL++GHgy4XGoU+V0t2/ePC03e/dHj+RLJmpjHIuZtkdQ3hE
6nWKwWVdduDaao5PXUM3uRIjkxfRDMZQIhiwisAKelDjrreiwejeLpoImRWvuE0ccyXSPA25+p3/
P+CufxCadZfa0CWxUgx6mWlfwdSNQWKFdW9gTrSoy62CHzHrifhDkeYLYGy9qYtAvIg2nvgaQpZC
p7KWkIYtPlCcMDm/MolRUK3hRsgmYLdkUdXhrbPeDsYC1BbcZ1sNEwELAH3J/wcGRbBn1pSVzwTS
CWeJwz2HXsI/+6rKLNNmj5vJjxyDFyCFIkUa5gLneFxnJ+RL4VH8UV6mtDnuhVeun/8186BZ0Hec
MtlacCYV8g3xG2OLFbFQpdHsqrnbIEF35a7P+qPP3IpiL+38hIAA6C/4uMbF5W9Pr6pfnA3yCjMs
h8v1E87jl8r1BMjdsLqeBfK/cQdwyhUdFIjhkLwySD087f/fUrcAnQ5ICZ+fyF5/l0RFephJxLXh
fpY6IDdkKF7QNW2WdJrbxknx5WGarj9HZ23d7/6StSN5TETlKMt9cOY7WSmI+BHkZZ60IQvjPOGH
ty35hTtJJuU5wFlSMB9AoqbH2cWWTFEUv0fRgKi7R2sXuXJ03InlwmuqSZqiEWJfTRf32SPB743X
S3sj3Yk4BGTgwpShg1l8KbqVpS4Z1ev7HUo7RMz+wx0Zsp0MT2GXgPJ/73MD5bAbpOrarkVp7gN+
kT55/6yNjFv5amiVR6nFbPgeZcOYGnFAf0a13x7ob/4UkD3+uQLtAOrjsprw4LKdovJ2aJUAbuU4
Jy+dzGppi2dDPKV4L1Qhj0vmz+fwpvjYwNVMBh5+KGPwE2VV2F8fYpfhQVyVMob3qSc/iEJKFbIE
qYfJADLnj86gI49so6wL3ftHJtQ2+q2P0gq8/VFceluENPiXwoYZz+LCvGZZfUgommR+onE18ttI
c6z4Ld5xxAZj5oDtIvWD+6YkjiwK+JmzBOrgXTVS4Jl0+Oy9afRQfxZeEwYaUE5vXZfIFgd8uvcl
HEL4SS4vILubVWlZ3Wj8w64ggRDWOjsS9g6PS0vULnvI+SI92J9Yi7k0kKRfA+ODSLS4N+s98Ct6
Tpxviz+AQ2SJ8+iTFXCEChzmVl5jcVqVaAsHWXGRaDkt+qAX3ygjtPNBI5p/h/cmjLUBnYn5285B
lf51PHR4xy98B3s5bpUvuHUGcWm5wVpYKuuyeq7CruqtSbeouqERkbDamT7ytPWtU91bC2ttr0hR
KLAyoh5VRetxRy5sYoZr9ne+L/IuaXKTDJv62Z8nEI8JOvWUo/OQTCW7H/v+gpeEhIACxcZbFepB
MU/ejnoV0c56G17Mvfr4cNOofcVHEzOYoH3J/Eai+ktLCSZIDkWDr4f7MnmwKmydcFeetoM2nhah
JrDzw9QYfIjVmzg3eWcoeukxueb3P8rOW2L2/XCzLWKH72DIDyZVd4xjPCJbiyAFKOUwT8mPieOk
CvKCmozbat+iXP2DXojXUWTZt6LZN9fSJAtlj4dzd7Rpwo3PLree63wNPvHZ2arKXRJ/QeThh9gO
oflPcdM/29Yqq8soVu1ji8vp3J6BKTk+3skZgwbl2Q5hKZPJ5A15qNQVvVXMxgtc/w9f4URaquTD
7bnTKifxZBP+2oQeLEF7wuYepnIjh7sbo7c2zD5nadqmZimKz05Q5EDlznqMvOTwGmIQsXJcxSmS
xlrEogzPsZoMDSdO0fknMQAqhUarXzS33i/yznKR6EMHGFqlWWUxGrBmEcDfQNW+iD5y4Vh+B4dU
CQ8DkSL+uPoy2rTcGY29Lm6DredY612BTXiWO9zSedk3foh3bJD0U7LHuLSs5OMCJNh8Be3J106f
RNPyA4qEn/cyVoWCQmJ86uGWvoHBah3NSiLtAUYJKHlGc++NPV7HoefVMn13uApDDMBPMZjP2D2/
VydTLwKPyoptWO88Q+8U9FEfH7FElP5oeIz+O/7a3s0zCdjOmByG1lj69r0cyotmX47zvRh39Tjo
N25/gFgEVQdBpSVCl1b86slof5idmYslVxRqs0s38rlG7zUT1zQy0Eig0brEHojH0/YWt7lWbF1j
cX8RxktrJgW5X3lDy4p8L6HiI+tCHfblHOj3SXDNSqQVPJqmFq7k5AfwYXCBOgykpZil26eqJpih
8bqqCw+AI++HeSFFcjTZMR2UXhR9XSN8HeMsXSYkuL9Vr23va86gaHmamJ3HD9hM91WT2KG/4ZXl
JpXNscBrKlEP0+9JULRLJecDJb0BMU3LagHkCE24YSj+QyQcH4HkMuQ5d8GPCKE2pbqVm7l1j5RX
+NNtq3fKCOLHowdxtN5EuAiiO5of+dWVIxPC69QwyN2JK+Hr+ZPotRLyEbPh7V0ShCgEeqefoBgC
k+GTZ7lgxeuN0hk9bVYXzZnv3ha1A/Uu6GJVR5Bgi1gLQFuUiV6LpleDN4WI3iFsDSlEwFPGDWBf
7GEoA5iFLR3ukhi+e2cg5pGrqaVpKdwm2qyg2WhxYlzS8eQcPCLzXopb88r59I9mTIKfeTQlIZJ4
84W37W7Fvm5VgMR766R/cFJ80F1TA2VeCavcj1ysZfH83lECy+XlY37Ya36QlxwP61lwaIWqqtPM
ea3Xc3Jciqh5EQfhp9RLMWUkRkEUCKRgvILiUavimKzKMokwusfCLKEj8bErnmCO2djGu4+kOGC2
tx55baNVhcY0XlbXR9a87JIz1GUNBexDSpBS+MUO/r8OqLzUoaZnNfDe2bffxAH6TZgb70m2ULeu
lHxlv1RmDJnZfTrDhkH0ETi2C0M+hjQ74nA2xujPE1gApV7cr/neRIlHBfKLTKzVfsDSPi7Nv5V3
NHgtDVSUIVDzIk8KqN1DhONo3munj++z2kO30JWIEvabGaaEJzp3kjp8Ht+UmpZay8ncb8vyviSc
2Y6hvbl8x7hrFRZNLBARAadUuPOKLyzQkPbNBlqhZgpfVYsItWmG4cyeS8Z+sxhkrAZmpbOsgI89
18SVNaglM83LMgjyzOu+lPyP1fQ04gar18SbyGwXUKNlOYWjdB7lMXZ8HXKj3f6owjxdx+8CtyoN
5hYELq0FkfFuewSuOWZPz5ZMpDIPR3ZFvVidT59fy+9zkQE7rO1HsO/MojhjBIXaFYL7SKzkW7b5
i8+MzcSZIkxQXBDaHJJ/nK+0r5roneuGmHCzIize7+8IVMv+0k4NVOlyACcGbxFAs/oyvbxGS3NX
INqoEuuHaSGNu4Qv1AJxJK2oWSekKuM2R09FTdboR51aq/m2Ocu7SRwtPc7MJ3+rvRXkZnH9c/kt
PfpjMwqD/OGfPkjwR48XiksTA3wt5c1nxKUvWVP5QJkIEXMzr58DJt1AjphNv/igRm2ydSMPYi3M
x0NV3h4oy41JsPLgQf7p5dcgJ5b5aoyXHqMyeQ+MJu37oSPT/dBe80O09MURk/GSVBiRBcI11d2G
dSo6yYHR1T1m3Gl2z+AhLpFI8MUUBy3TjbQ7EaTSyugr/WsC1mI4nWPlnta6IjEXn1lh+r/8aUSO
wcuRToFfq7/9PGeNxB1pww8/2yCIQDV2G9qgh6IqX1sgrKIOmCOZl51jjZQPc1BRMQtFfIus3vcV
6WIqvCxUlf/RWMnE/87pJ4tU0QEAFeJE7vUBOYa4NIJp2r7lQB3QOlFMKDBbzN8oYZ/Z6z0qqBZb
PJEKmMXfQKv8tKGgGnG/KMOa+KdQ9zBo0f7zaPRLm6qg+0xiVb9vvtOUDgIrcE6AY0IlgbZygW+6
QVzvLN3eK2F8bc8OAbCqf/9hrasj4ae03NltpIly+lKojIjw5QMzF3OXB8pcFieNgeWuYYuRrfUk
L3sMnf913JKS1W0PKVMEMVFRL2bvfm2591g37cxkZT2RkIEJNOCEe7lR5Uhs3y0QWALYGSfOV2r8
yq8CuWewPYWSmeLJmWwKJB2DYzNPquL1ckLkQfvJSV8uHUOUELpHsWjpkBmIvXnGMPZ27lGrls3W
qN7wNUF+/bEUnFW7bzVo3m5w1xPwbyvwIUr2/CPEgi0t3cYHaa3Uh5JYDf4wCVgxzTtNW2GHIoU+
E/z9wBkn93RE9LkMHKtoBBMI4aY65Jk6IRTESNMIXmLogdj3fzspjBbl7M6iEoGtkK0wfW1tyZze
Syj5UQoqHi//x1Cg+cgWaG3RpI4n/Nf9dr3WrrKQ+I+JnoSDwOsr/yHPnQv2tTkX6+kF3o4D7c/w
HLmFZdE5fDStvpCkpwwxaOM4AGQcSS+eVFgoqrv+DB14oBcM5NYiOny3fdcaXdIpvbLoldNv/SUX
f6baHBT2mRUZB9txNI26XHb7sRUxxxSJOpWpWBsdTMX4wx5veVAj/NhEKAAb9GomJ4Fd3R2WlK/T
V3BwJ7ChxT9s+0V7UvQgNtSn5IN5F8NPYebfoK3LwiztQ8+/FD5x/sJzu3/vut6Sze6+3+7Ym2dA
xSOW7FasB2oB8uu3YPamKugnHYuD5G/rFpwMlPzlnkUrV9qLrNGGH18exO/FnFiuGip0XRpgNX++
274C8RgVpJ9jtEiZVDp4N8eZQ+4wSYlF0H/WB41NS6VIn0Evhj1nV6lEQg94Ynvp1nWAmWqEAbEE
ASC8RG71OVhEamVb/dLpd/+BoykQ18pSJqVUjvOnX91m0DzQlXFN2jR+K2jCfUaL2oRId/H5RiIG
xiWfhmykemKofwaB1t3ysylPJcZr5UR+LQP5ca+t1F2VQ19gtJS7cV7xqbub2fSgWitMgFFaIqTP
0WU0NIjhyWbbiAyIw3zQerobWacT3n5xPjV9v7pnr96j9Lr4j7oo7NLiTuPqgeL+FUZVyu/LRYUg
AlaYvPePBcNhGVYuo5VD0DZCm+ALi6z/Y45/7wwm4el0OJ+5nKyy/fz57r7bGLSqV8LA3e4TU8mz
Z3kTq1KdS63F1D4mW5w0ib4lj/6dlhdrsVE41zkDltIjDRDFGRXQ1DaXGhGSSljgfgL/aGag/XpV
NNOIr9mBqQFHufDujkjKeuFGve8JSksq9vd8dnqNwc6oMzYg0BoNDW951hRj+vcEiLXqzER7tpg+
ubGewS5RAg0E2gT1tOSIvYwWaWjYCHtdfvTQ7uElbUlWEVk+8Xv1zICt1hADqV/tMmri1bapAbHk
fwVrSJ2GNwMURf3/HrmZyTYh3GtVyVxlildMddXleJ0ky8t/+gUIV1N08dmpN44dUJ0qLyrYnjEW
8nWyu4xUwF4R54o0f9TN0di+/i4T83u0jP8cpbEcbyB/Z55ZSr6LUPBbQeeghcq5zqmVoMxv8StD
tsoOX/wxLgazgnpi8H3prblmnFv/vkYl0ppB8oVitd4E+ziPoXKjQB7V4WuBwfd0Sq2HW05MmNJJ
+9UR3QNVS0GN/upzEvLEZ5B9olOYPbGCYSKH+vwMLyJaTXLIXI9tYuO5+e7vctRcyfZP2b4lTtHA
RsX6qIEpPxiPqkLwGxQRHOgyWs0Wnub0M8vW6QP4b5bpVX6ccAZL++LOuVHx9XdYpWtjMAPL0neG
ZucplpieUldu95kj+NhdQNeoKZKqn0BA6GCws9Jw5WByW8SZINCXETKiV7Egh9kuithmlVhv04Wc
BZ4rXWdkmMy2HtsHGsrqXdxXdyBp2OAtcdYkqg+uZP/jbfQuYSqUtevpF3pKkGr6PlvD5wOSv9nG
bxRo79T789cYiA6+qYG6+LTSLmoCE9aZfqrXoSu6VIWT0n1Otzp5+pYsNiGTm5Ah5ym9tL0hAzRg
GbHkO0My2K0++vbg2Ou7MgBdVKlOxY5PA/Q3qh0E7LutoZjk58/vWetjkgohmJjGJxqq5Tsx8Sn+
+znFFPrLFYvLLhAgloaJDxILkByB9aTOeS1uQb8Xaonb7BOKwP73QoFOp4umNb+gZfWfCObAWMOV
CDmvdXNLH+UDDbd7/uuqYwsRNdMp90U583QXJeF/+vwf8uBjuwvg+gISMuESMM6GbYPSKYiQB/Hb
GkzVRMRf2sVx8+ePcqd+AGF2Z8TzxKSPXDg/c4b9pcZQ1xU5B03+wOYl747g5T3+AcHliA7gFBMu
7S4OlvLCp5X+O7TCuHp5OP8N6V3Z3D0ixjsWQYN95yg5S9CWkP5o9xREFYgjtQoIYUNd2s/B+IxO
h0rDmYN/X3hK5sOBCitzk6uiNuKcydGYrOjTRZ2ZXj868jO/+mQmddK1f9BTsmdaAwHVsmI8Eeo7
w0mhQanB2bTwXP2n6l5DZFVghgEvoi1W0bF6gQ7IACFj7FDZ98sD6g9RQDtadkPv3qof3qL1TT1b
Y1ZM3WQa1yshutLAXo2Gra39mxQ6ixp/r97AK9YUYf0+RW4d+NTknw2KfeTjcJKVx/AQDERQfYBn
5+rfrX7VoMLV/CC0sC2hyHsbfUkmoUd7T9Yw4qmgqYzfrAvVZOg/ATI6IDkTqowRmvck2Hv7wMDk
RXEMDC4TTvw9yKoamHUb19Ql851TUmHKw1VhNu0Kj6KuufEQc48xQgoxkq1YHxqr22JzDALpupmA
AQzTInykJe6qc4LHFJj3a7DC/SmQjfQu4pMu3vvN9ELYslySWBiCtsX+AV95rGhgG8jiFwfaWL4z
jSIrXQTGaX4zuAqHf4VnNb2ZEQxPCi76SGKOD8K0xx/WNxNovleV3tX9l2NPm6mUgDeugOljKxpV
/+72eWahNe9rHBcl/RBusmnp4qXd7t40jXCRiOdvsKYrfHQgFhi0f+XU1lIDstiPzFHl5V27RXjJ
OuvTgjagZdWcrcDrO9RI5jXQm9+tHJU4dJCK4HljidpZ0lM45Kz+ro7iqIUR3t2YPi9llRoE8QPI
kNnhqlBIK1LzNPNa+Czd5sfasNEiOKzb7OUIOrUxR+Dlt8cOuRnfCWEmyAgI7jGOmudqauoInxkY
5dEjvap5G2q2XqlNWicP04j/QqV/5TVMaKxSh1BTAvI1Jviy6/HOwVPMTVU45kyLllHwGIUDCa9Q
nSL9EwY5WJvr3rTp7s8GXNVAitAjVzFmqL70kfejr4fN1v7TexaRF8moXyQjUnbI9kJm9a6dz5u9
FbOq2wxlWmRCb9oq7EBViCBaC83Wb7BrqmjPUSI7ypuEqWdiQvn3PyQKUzk4VlHwZIJVzrFx4+4Z
gDgggZguf2feNjOhBpy3wX6U3cmVWrqFHEdsWHg6QZfP0V+d5wi9E0hSFADlYd43zMsmd021OcMG
T5W9R9jBIs7SpnXcWUAP5/J2njjGusG2sL6U+ZHNkfItN+eenZAw48qPRVSgc2Wr8HfRpWXmvUrq
g6Y3J47M2uA5pb2tt95fsGnsyewnez0taJeXYEajcPdOfrUJsZkinbqFJSdHRyddhfe2IlxQ2MGq
oZ9755IpSteoloXHIQKAH5XEOP7KiZpTjuxh+ATK0S4qGTsg6km9ytnwruFm9tDTr0/1lLPzRpph
g10fqVqZLz5WG2JFrKuUirb5q0TFZrlVeH8Db9cg9cZ8EV6mSINpDUPUM5T19GgeT/MagIsvO7Dr
1rF3MWZY5NWVi+nZLsmMGwiZxyiTW9UW+LNYU5azjSaPHpAh+Z7dqVI1pVPXTcTSHmHq3EdWRMAm
AYMhPRnbrqQus2ViTMasE7kURNT9bfazevMCFawy1nmfqi/J07rcn3Kchsf43ZUx8vAG1jBr8fOH
Z1bSKZDKd5Gp8E+4Tm8nCPcdYQD5qLLJlg446NR/ZJ8OtLT/KqtL07JrQGpw7CwO+EzUXyplOD5C
ZCcVKHhETo9EdaKiElMnFxGil3x6DVGWCu/2FSuciWEC5ryhXhY/rqW2rcLdgrytfjRy1zHg/Fka
51afJLMbnVt1e/xkFJw2VsJErKLrphwXTWHnz4hpN3S+WpHbmjCflEQjA+hLDcdwBSBEvM+z6g+S
l4wcBAYEv8OOQg+sXpl9FSvHFp6x+OkZbJVB/guoQOYzezwc9hczkz3syP1xHBhZ2tAooEwxrx7D
MOepsIbmE5MJJtJ4VRav4U+etUt6ZRRenPFZb04Kl1Q3TM7B+GtMr+v8oCHs5VW7xB69OEjet93H
eKAuweaMiwemAB1cxOoMaT2Uc93bwg65FgLLo9DIksOuAlsk4kdy0mfa0ECJf1wm0sm55nMDd/yo
6Rc1yfqJzKszse4R09TfV7o89M9s957yKY6EyNBKQj2Y83fTxmTwK7zUakQk5ypsNlot8NOyZFwa
0FxXljhbce9odhIEN250rs+I/rNmZwFORkbVQBxQE4eMUsmM/CmrmC4ZARS48XZRoLCZR+Os6fpO
JdWU8xC8CH3mXybdrirGr74yau+WtNeswO5LMzU9GahDhnjmPtKXU1LTCpLcST2Ss5o6N+p/0LCg
HUlw25VgVcvVqYaTAk5/yKCs3NRqrcwWOJKySnJSi7OukBoDm2L2A3p6IEIl5h7zNh4HOs7nBIWb
57HPwh+ZxklFBeIUhmcfX42XBiP7dKt5H6OI+iToDBtcpNFt8UKm2qrxkhOG9rBHf+tFij1NQUTu
iswILiSigbwWWAvKuXYJuQ6Cs8f3WEcwKN+2LvBw/1Mf4ItIhYw1vrqILEnu6OLao5Dh6D4suN91
lPs3Ek8jAitEMP2yh4PJOAoS5tmSohdyqv9wzPHOU2J1LonHmbVBJZkAZUdmLmnZVCivvVK3DcYd
SS9vCknVS/56KHJemHQTjdEViMlXoJuIvTxZgPwS28a7j7v9F8rIuD6i2vV6GKtVDlwi/3FUiLl7
xuTQKsHwOCKVGH2SNo1l2fg9jeQ+eHTd/FEfL0Vu9rGaK5mphc22R6CqQdLA0Ts5zztk14D92Eq2
uKA028x2mcKisWfwMmjm3kL8muCh46idBSYzRaZOIj/sNRbeB8Nt87Zqno7wwIlLVOhs76pFzSRi
jYLa97ad0SxAafj84bUKjrAQBceOvzrmfD5pDX+Dq/HJu3bZEaJ4RrH/DZIm4Yv0rJeBOMCwt1xM
pCaHomiUI7FmY4TzfpkR5NIJCLoY5vSe/I6Uhhj8KUfjychBvKOrXjfnYXvP8aJbOKw9NNJHevqB
8cRUa+kNKlm9H3txLaHaRxwEuelWXYX3dnOXKujcc7y4EjeP4ilCMtVoFKNIlugIkrLUlQtwFiGq
lt7o1IxXDOuPeMkOvl3Z64GcHX8GT7QfmMZd7ettrqVw+iSKVqzh8w6Qz2v9SLsigCOfyZVc2BqR
ekGz9iOuVBRpR0S/qudd7DTcFQxAO/gvMyXtSkEgY4sMJj8a6w1PACJuA/CjzwIug6BC1BfCfZtA
zEXbcSXqe+hvbHdpTiKINpl8jsNCR0pSnXquUn0VP63AdOKg2LvlwGxmaY8NQqCnlVDIo1IR1Tmt
wODwCbIGsAZkpXer+hqymPamSutKiFK0hvm7EKwTqyK8YbFCKwO0pItvk/qxLTreCyLlQWWCQA7G
67ILDhk0aVf5gMpZM8KbGgDHBDIsFKGTFNUdtZBE0JAXUnJDSequ9MyA8K+3bMqNCfopdJ37Dyd5
9mOiKAukBVXJ/UA9nKjjWfL5L4bQRiv6xLUrCSsjc+8on/XTv+w3Zg+tYnfQv8n+fcevn1uK5R4L
n7n9to+/VWmrs1HStalaRRwvBjAPcVHu+fSvLdotH91oRqiqKxi5eBE2Q7IODDjUqZuWo3GjK/Qq
1/gYe4STyyNiJUF6ICNcF9kpklEsmwKJLSyIKWKSdsR3PenU3XCkROrCFVFzGHqZrB7xEl2g2SCv
HR3O5haS5yTr1s7xlM2al7Yk1UIl/EYkfseTTb7D5gYO5s6SyYwfifJfTphaZIldD6LUSVCUMX2p
xf+PPXwf9mYGq0gGW4F1y/dOFk7/LOvWn1Z/dmy3OQRw/IdVeN808aR5n4ohxywLSo5rYIJcrx6C
dsU5QWwQMZwGjo8SxC59abRBqzW4qgDOcL6VvfxSTywYzy7qjT5sL55KEE55a71FMpakarM/tVEP
pUGNKdC1K59uyiJKMlKt3QX+CV1+YU3vcOQzVXKCs9Ha9U1tHdze3HrsQr9Vx7fPZEFpQw8zsIMS
boicRI7/qWWQ2PKClva/6JLEHsQilFSwB6t70NdWWk1Q+N3mQChSVT7C1no9BryJNsBUNHbzciew
Ohe/it1Yxvc03BtF6i70XVkYNeOq63fMV68XsUaArsAlV1xkokDhrCbIPrLIzpqZPPNl+++cZG48
dci32+Im3FSjnHD1de76HSpAyFBJKY7siJdAmbt5dXWF3WI9ow8xZSdvZJMCvsA0guqjYIGeyk/9
NaszljneHGa+JAeDtZ85VeqnmfWQI5p4rxJqwXLLecx51h8t50AVwgGPLhT/n/16KPGuX06KxaIB
sp2XOjEsMwTylQFIU0cve4Zsgye1u4lHiabnF2qSY2mNK2/nqbnwbVI6+flajcbTZGDrrT3E352p
MnhyNiAbtjovrgU/NIY+34iz/kWYLKH1SkdepR/4yK7xu6uOFW0iOI+b+IsbeTP14c9BYxIlt7Cg
iHxoI8a2k3D4+ai4sZoS3FvL2T4+WuGZrwGKGF9vl4pKwg1Wi0STk6VUsmLEnBRhXBPkRxjIHD8D
dD4iZ+xJuJ4X1NqbJjI5I8Fq/+bbHAPcO8cx9A27dKvTqX5UedIX17ZKS1cIYhjjpe7pd47jcyy1
ms3w4qUeTUICV5cKFEgv5myGVnFoJydVFm0ba9cn2W44vC1GVjrtqRzFm42yz0rQ0gvjXDPzwIgU
mv0hr6ZMqGoY7DWzGyk7Y2iPNiWAjDq1wRn+cBkp4+YfDRQOouKu25a9VR4fxNwYlGOBQ9clqiNZ
QdR6LzLLfnTPSF38ytaBLeToACTlwuuI0AqyUi1uhF403SPbNyQO4PMCFhpAan1XgJN2unnQeuBX
bpmhcgPAAL1aS2huXpF1Htjw4uCnd1rSiaYvRjf2ZcC4t+YAWvrNo36Vk3ES13FTcxFVB2kHVGzY
2mCMg0P99yEo11OePucvUCobstrnkxTjliucTK+0L4Wacn4x+VVwC5fDHB6Q7Zi3bwVksP44TA6r
2P50r8ZytKVirgrjRi6F3Xt6ZWlCbpOooie9i250nBeZoS7SM3iMBwfebrtpDpfj6p6vNnP9/Avj
S5fFwlX22ooBH7ulqxWmXRzu7xRt5pfSn169iw10bOX2y7DlLH42vciWumI9qqPUPCPiDJthKzTd
uBscCXJcwL7F72WybK4Ix69vGqr6dSmYWmxwEEQ+HHXlIkfCWsMO0uKJL/J7tV7dOOXRxmmiot3z
FZ8iUwepJlBpf9MGlD0vazWEIjEH0NKm9R35HPqftS7HWYoq2iKat3yFF2f3wkemwru0XXSwK3qt
qGttP7zN5Xd+ME0kmXXCqevWfYrcX7K2T6tTEZPDFtvIYq2ZIMfGge0Maz8VFk1KYG3XCLeqsO7P
sGHgeAk2ow31b9pVW+bgz9MHfiAPkuq0PIc3MbH0bquzqB2I2ac7ahrh/bckyJEP1xJo6xFFM7Df
MbY5OkxxE62C+qdW4llYl0odtnUk3j25AYIQBgVcyfju0LFW9D+k7KYkBrcMjrIazEGIxDDSIzPu
4GooPsGA+K39H/ySudXg3KKrr7fHbZBfjGqXe3p9Cjl7BjvXZBpijFwMgywbVC7QBtsbh+8Glm5c
t1aqUetSktFvgOoC7bauNho6M0+GgL50EUr6QyLe+/eMbghHeFpaK2sTshAwjBFiH5DZHDVs/JyL
257meD1L+UkuEfRZfKEMZ16uwb0uUsNMUnCjeRlhxTF+xnjAxNc1t16qr2K+gtgObGLXEmZ2U0qA
b1VDH6EkwUCUJO2PMZhDJ/kT+7tpOM3aKUySD+Zq5s9ybuvaTB901+k8dyD0sPwj5yBpIfEt0uLw
HXWhWCKGJVnIVzNsgoIDjGgMiEvlKi3EmDAyOQ8Xaf6GCwdHVtI/CuA7cyev4AKFJ4TmrWSQpQgA
uBJ9bTMMv86u2UPMHwfz13Mw7hEh8PbNdiwYPX4qtC0o98FDdgt0mHIGASnT8IsVG1fiM27uoCYv
IRyyolyhgm7DAZDaaJVJ5RdT5O4Dx8pT1AqSy7REHQ5dKeQBwx0uwIsob1rOH4ODnCmavMZ+2+2u
qizzuLKZ/W6Iba7KzPO4QOJO5CnJSsgh2OX2cL47653s5gxG5VulM6S2IreyNSsClCZmVds1k3le
sFvmrZyw39mkm9T8w8HJ6+bRiMptllmSGXpnQIzjpLQ8xU3Jt79Ntw/QAwfIbN4OpW2hWiBy2pul
n6h1S5OxH/hpJWwpgyed1QBw3feOzvjUkc01nrxiZUdTKC74gGF/uoQ/A8BoMmBskOEiVZI9fAim
n5GSiQdju1ylqWthYkPGkVGoZgjxvCnLR0Vjt72y+oQG5BGd8CF7TkiAeHR3KIgKQ/Bbi3XXlyGo
rp0HzUTmwqZeugr/uDePydkGXY1I2i03pDz9kt7dn/taipaSkYmOB5OQtVI8sxk03+XjaBUloUrG
r6G00Et1V9O8YcUvnRzD8NXnz993CBDFoPMEl/5Oc46rNoZ2al3EmwabObMGhshCeA3MR/nPvHIZ
nPWVaAN1pQaVqSpLdXaLdWaupXrJdCCRJu7K3tgxdro34xU+k4s1wPHkELYfZgbLFYXZSHAfqvD7
7KXtZzsJCuU1cpspTDj74/DT9+S76znXt3vCn9/dborIFuuYu7H0zinM6FRTC/6YNL9L645ySUKp
GmnXDxv726YBW136wgmoVTwXKscT6wikeE5SZBaEuGRdQDfHs1Il9nbAye5HDSKV1+ME9Y14bDFX
QfHj6YXtxnXQJwFceLVuI6Qp7UvA++qTEUBwyyn8N4eIWYYJBCu6tJ/FrvegdEHAsJbMHeUDREpo
Vz38zVPSGD78LJKFrxbm31PMvsXy86eLoICRX4pSL6GOjHOGw/5EZanXWDs6SD2mTySUS0osA7xl
yUlCtw9VMUd0jX6PXqvpzNQPtzfGClkxltOMHpqtLJ/AXJc0yZ4KLqPB64UB3TcHT9IXmAmv6JuC
dVR9UPv512YfADHjOy3EpOPW4g1LSDYeXZLH5e6VQgsO5hhv0eacNpVjA3WZvO2PLMtgFRwObEdF
B553TMuxLMAdouxrcB1lsNqR724pr2BL4aWe3YNCDmfQhWmmc8sdym38EH3WxhABVduD/B9kVCNW
evkjloyGJTeMuqsZ1LcJIyTqW2xgdF++ex9hOImqPTN779az54huskA1xsWWBOpNAQsIxDJdlKpO
Kq5wMPL+AxYnZpakHeU8q+XzwKK7nrAYt0NvOHAuhdEm4UOspD2fWuUoeb9jwERuLWJk/PO9a+Xr
Xyx1odO9b0BH5HRYUeKK5+EdpQ9ap5Lz8jRDn9uiV6qQTvaFNGuTmiNKDtBwIRGDh7GWPxDHXuai
A6WaV8mwt5Jdm/nCDk8gbIe5lBsfxLWRQ4TiV/cYik3jOYcrqRD7PVpS2LoEd6PtjRe4Q/CsCl7Z
2vEuVrmOVU8NXEXsMOzxliW9Y4urMuwNZGJ6cOsbfWeJmz2T3h2Nl0yGanIII4czC5RhAYGy6c9o
g82/n512t4MSEI8wLpBjXUawtClijWcHME2GwxbSqujAxLY7ZzOsJZvotnG+H/HUQq1nRNgeWBJ0
g2CmhfTOMmkjW5+57hMUag4EXL9WvMvbEqEkUFtrP+JcZCK1LqwlvHB4bhHKSPDkChnjLqewto1c
zDoa/KSKU+o3/hPZJ/exiFujrMvljVjqXBHdaxNWW5RffPcNtiRAvx1DpMnhpaNoctRWEXwOTZUi
VLRnA+e71fyuMP3W40taHCd0bpaO97r6ym2i+/oc9UFYd0FWCDzXC8ulry4zjtXT5C4hzSu3p5gA
y9c1lGkBnlK+GtQdq3GxBThwEGsBFenkKSr0rMQZKlpiZwKO3HM+qgK7lXiqGBG5RUvMRPUqFt9R
8pKxX7vhcMuWVwJOiHYC8hUxUuTMy4YmereTNoU1HzrlfvMhuJUKV5LVNbfB3eom5iyJwkVmKd1W
Rx43fx05uOKDL6d5VDzyZvux9BZVYzy5GdLrsrpm2k5DYOD7a8GKHCKownjzkwataYO2b6IYq+Uq
cIct3MaisxWKkFQs5pK2p9/HqxjHH87iEEZbcnMEMwTZNaj6Pk4fcUgB3jpKvv3Fduzl/zHvhrMz
lXxv0NiQjSy2HpPNFLoRws4fy5IlA+1wuldhemT8E4akr5/cgdDGq7OkiSSHAkxVwKkV/mG29anh
PDn6C7y3b2T11hJcbDp4ADNUXx3uvMMdLWzoz1Hentk/1zHPQiVGypSQ1D2htab/9W3fF08R4i5r
2UwVSgXxLm9MNhQ1sjizhLvymX1Ok5FtRwrA119kGd7ra4oYizViOvfdDtB0kwLm9icHpiWbA37x
3SEdmpzY2aFi4BVWed9YH8KPnz5UMgF+BXkzOyipkJYTrElz2TqofZDajflXfqnl1Ki7OErsNk8D
t4kpd3KQ8zoAi4dZPZdmiReqyXkO9zhlKof2id1UpfwSCd0m+Uj7Rdst8jAdpi1dka8VczUwBkdn
MZ3ZtCKugoRW3DaqrNsB91r+edFvfuzQc3lc4mKIO26Xd3D+L115yjYTvuK+q6a29sYLFTDB2wSU
FkMhlGDSt7ARvAxwC1yVo9dRCjtlVoFsqw90L1bysxhKwlwT6B0ngCViK1Wc4bW2scRAB1Z4CgcG
YSNawfgQyUue56XSmZChLxWEIkF2qRUnMir9GzEoy+BN//ZTFG0lctdNSj8s/UfdeTMk7M6sT33c
XgnmrnTZAw0ji1fEKfztv8ENeVY2/mplrMLSyhPJfHGK4x3DLN2lDogdNF1Q/apGjpSbA42IevQM
1p02iUp6KUb+It528Yt/Bsir8P6H1HsSRXD/zViRWjZmyYTScsnlPqR34fv7dvGJWsp2GTPFe+QE
GVSF0GBhCKSyamHejbgGV3k/k2/vj4alIf3+agC0SN+hw6Hp2CiJ+Jz+JksAvhXi5kFR2nhLMWKn
+Ns13sNvMKu9exB76zYHIk0trcAHh50L4EV/hnN+fT5/tgXB0WE0oFM0xUu/JqOSge4ICvDWtjtI
1JFqLXcaWIRJVG9TCEZ8VhgHmmse2jm0T3xsFqsvqFUPTX6PX6bQPKRBOO0/Mb5WRa4uignVjRU2
9tkk4Ab0IAIAm00O2Fsb6qy3FnCUkIdw0pgXmuR21/cMXyDjCzy2nN/KrXlTAx2EHO8IgoI4f7r5
IBv9BYSSCFwmzTmABKpgEQb4sFe8qBTvZGQbzknslx6LUT22jPJYbJAWY6EbWqwrui+N3LuBZ8rd
dph/0t0xunXmd4uW4TCG98EYMDbyyJExyHIjBdwgF9z5uSlWhIXQZgZlHUcdOfJO0C0lGixr9F2D
L2MAK7xAXulXi10GpgqJs8I01CRvll/9KhNINt93liA3fEi2QPj3VGasLWf5HGkZsryi7yhiD+eR
RxDaEAvsolCS5k2hFJ2P/VHW77FM+JS1LA0L8lCSQ77/U8VFwaxn/Mc/c7QFgiOShJLekYaGSlWh
ukMw07stxJRSibhlq7V48eFGTu9pztts7bdaTfBiXtZDHt+gTPzao0NVCdMP39NRJC7rUvv445Mr
He0TF51+GzTWXhgmXyqPZ/zfvpmcZzaup8YQxjKs2CSBKYxiKrsceRyGbVo7mtlZbfC2xD7IAKf9
Kx/u9ujk7Lwy9YMi1qtSetQApJpoNkqffXGxsd2YIjVtEsEBobMxMllW9dzThjntFoCO6HrSLAB3
4/TbcUQyZOMyPTERm8IKKN/9KIjzOOABgfdDDcvlv7Razg4PpKwPvc2zrZycsxVYx+faUzSwdv3u
A1HYdDIJzg2vaoBqTxdW2HtYPX2nqacgsK4An0kuc/56iunkQytGbVBkLoMfZj6IImbiChsscPEW
ldLjL3UCt7ZZjK3epCDdfk9JH2Z3nzR/LUeCt5+y4D+0z+AmvuCKuCPRTwHfZHfPv/AD6zYbiZw3
otdgahXZZn2WOKQbAj3YbL2VTh7RBIFOPqVfv2Mkrt5Hq07m5xcynV8Vn6w4hL0XBGykbH/gjzJt
yvgzU8WSImLhhELRD8OQN+NxJP18q/WvSqQ4Pry6JFX1c7g6/XZ5MNRSNCmPEp0l6KOZP8F1NMbD
+YxCS6g8S0o7R+ZaTSlObu0YeE+qT9so+m/+Pyg2WWvmhUP1GZnZxeKj3rCaT9h4dfY0xac1lyVG
3sMi5/1huftR7MsWdHM4DvRkQzHZdEPQ5mGrpQCcReNphsEQD4eBWVfjBr0/ZxKPB+EKR73xDBn1
MpP8hkCuXJLrVPGCNQUlCxdfQu4C+4XxoIQoN6EYFsf4YZTX3MDFOTtkBFufXAx8TCCMLbetxiPv
jLimpcNHMAS03ee8S+Ux0PfgzmTuXC4DNFGw1P+sgomW0BWVGUoXu9lDeJ0oRD5JB7yDkmFOBYFp
Y4x/kGGza/B+AcdGZ7Hcj0t3qFhdcPVg5pMI2dlMJkk2R7l0SIuakH2XBQHdIrAzF9xO31r2gV3Q
RkBGT4zUaj6HhKcpyk9sm6Fgh23buq/3LnlYEvrO4MT9ah6sn2Lw7vAM1nED0MQNZXswZCFlvIeU
tUBFutOwEDkOwi9VxQVPFOs3J3ngIpmFHybwXJpwyj9SXN6etvgG/2Z1MCi2utJUPiHjb8WfcyZV
5uGgEIADaJ7aZIQHiYBzQj1gvEC1maigcwi626vpuMl229x3OObghk8fhSy+NnUb1WI5u0r2WBkS
09GzGkkkP6ADNG2q5nTFd1mZMr78s58jJEQDdi3KtSkTpTV98kBeJ9gMWZA75Jbcr4h7ag2YTk0P
d/RJrCYiqGNFaLAzveO0l66FUHFDQnrwaF7y1qO2M//woDTv/W5/fB/tv5inbbajBVFPaDRHvP8D
tt+fqm8Klw3e2x26yJWz3sMNtoBkN7p7Ol9wpgv0V/OTRtbzk1FU9ZnFe1V+WwA8HP/ugHcZaPaC
LF5oMjCdYq+W5njoruzWwRNQ8QE0BFkjNC++QqH1kbamMj+Dj9AguQ0JXchLKYrJ6pQMryxmqsbJ
nj8BLlx8uWCcK+xZPU+cuorAD73rqp/yG/AKtzFsz15TI8F9ToylY/W9YftbWPchfvRRpEt6mrWV
5laMda0vqCm8PlforyhYaeLV5tCT5Xey6ca/HGVi7JbRAmzhNN9vkCqrsoNNJfzBE3fFCH0dg6qB
xgo7eWlx+q4toA5gUEGuhWYR7qUXIDYDbGN2rC1Zr+JBwURFjXheIudWwkq3uEjEgLR5qM7GLm5+
N3iKlOBk61K+MQlE5Q/KvyehpM2Qa76THLx9Y9djMWplCYykvIXIIKf8oY2sMHJtGeIqy/+WL2/b
QnEolnqg4pdpY5OoDF/cT8D+qa1lysxnut63Cs0FILxBSmPVO5oGm97VTaR97IZcXAi/9klRIecY
D4sR9uZMq7i7Wk1BYS8ahSPf8eJX0nSSv2dlo4N6mL4dVWWYLG08Q+2B6fg5I3JFuKVzeq0phfhB
HVs2pj5Dk5AePs//0IIl2xuXurw43zShp94kR0Oxk8i5Sul73vSXUEzlpUB0IzutP7kDTErOO7cB
AKEePpj9cGim2etojNzq19kx0l0qUMhzg3coQ24b3r+zvDl7MjSsEPjMPruiAuHuF5f5xyXs8802
ZoMyEEbr3BS+wCJtWNyAkCw9f64dmGzXgyG8UFco7Qll37FhpuFxs1flcBkF2cjYn1hZZxj6DCN9
+z1DsL0m1OyPOk1Irmjnk6X9QPSe59yfxFuXLtSx6KqAIpbk2aTk2Gxc/I6rS4HH4EJsWYlnAS3X
JR0wXuGzqvC6UD87nTWQgrjSsmMMKJnRo0BfS9QQ0AhCIAYURUqIxzf63EG3OnNreniuY6XXve2G
39aGLJ7jZSbICXoirWUJgSJg1NdulLeZ8ykarzgEpgfEJqz+zCDnl4krubIDYvKd5LUC6Pc3xNkS
19gr9z1ZEbGTDdCcQWYnUWd8D7BpfPHpGaHWoWmnymhk8Tqih3HF40lMv3+uzYh2aLJZg++mFnjv
eILyrk0qqd4vglPAmXmYPjMN2jQ5cWFrGkkUqplPSgEgsgUweAxTsSUuH1F+KG4t4YxEvM+JpCdq
WqE0kU9IuENXrYm/fngew8J8TOw9sWiPHj4K43FfdMN4t6O6UAV8Ne8gLQvD6ZyCvCjG5Xx0AzJ4
6CR3FL2VTnzxQWcdKToX+PkhhJZdnOujxqJ5rrIOfWYhOOzFlpVRBK+difCeaVV4jTbCYHazFiBB
jvNh6NJSJIswPDKrZctxhbyLD0IkZ8npHrOywKJaT85dTG+AqdC1fdT/dLgk/rvXBkqNOGV5k23k
x7XKpqrT2KKJ/vhN5Q+aZPzsOrQ5CFCEWs1RoqVJ+2Z2zDkAIK7d7y9DNLAoJoI/4/zmS39XP/mt
3gTEfiQhhycqUil9KOUWkgjVK6Zt1bk799/GLpIGrt7MTGy53hfrN/BZftG2a3W4WMGqCKe8iBly
61qtXr94Cqt7rRop4mmcH7o8qlruoDtonBJEreNAZpRXV+kHfCQ8gN3Eg2HdnuGL3Cfz96u3346D
IHIgeD5a/5qUqJMmUmcfnFFuwxVd1uxyypwH8glxwUhFlB3ozgiQn2jEfr2Lv2ZwdS5VXGoG3EHp
PZ8hRoYLDkwp4XG/dkPX+885sDsTK6sKI+CAXZzyty/D7JigE7ciynjx2YmkcbAaB5WmWiejWKAw
qUQRyILdmEPjtPRZFcDtdWesARdkB1PwRo3FSIo86on76Gbu99tHCGYipRLK6h3dNG4YwGg1U1QU
zGQYspGu5LWIjvijuv7SocTgY8lyZjud9lgqmOKxafFLOeGEvqXVde80bhfbvHC3R7cGgZcDiECF
US7zhKiltqFN6ZmMLzo3Y64N3KyRsebtL7Ce7LN8sdGE+cfqwcLAGdGl3x0I61uhN7BeHFACuXEg
mgQCLhpECm32uE0kA02ROJ5SdPkSU/xkCgzvVEc1DIFT277mWoS5aNj0KS/Zi/wl5QCF4AJ6hdpO
jy6sg0C0D2Ez60hdJXkPESkk4pIWwCKgmcw6REVGzz5cVdcSNQcklntGU6uzRmjdKILbzjrjHsaK
ja3WhSN4tIsV2lxCvvkuzyZEFCf1f/v1ZRpHPlehbVtn7m+WS2sbSzvz4rWsGK7zVBG0cHxAmDZf
HxgNQk/JEeGWBanBaPQaoFXaTZmDi2TQRWEYmkwkMwsgH9rctdC99zwLLB/Fyi6YmD2UBidFiJTR
/eXh9TumMyVa2ggQkWuzn/03VuEggcSf3ucpKTdH+zk4pimlI3jwduP9EWMVGvZzOs64fZDEG7cA
IPdcZ4CPA/vO2Jup4mNeTRvgMt5icViRMKFejZJaKBr6Q5MouHfNnIxuJto0r1/9VcasD5TGYhCk
wb/EnilEIef4U9AaTCtS1ozSTeQcikw8S2HdVTtr4Dy08b0OkkLscG+zpgICys2uJZqL7gczupRf
JNe4O9R8sb70Mwd3fYgRYNfJJf5q4iGyEFqQezOBW7CB4b3CL0yVVRWMkfTdWpScFP1ijkeHUoBM
nGEezlH4RU4lZk6BS36hosoCwsqMb+Y1YK8xbi+zmiAT14Tb9Xvl0v4hKaNL/ta4it8zZlM9h1it
sL7DlkjlYy6hkFZeCjwR1e542yD07NQIMxlMi834KcGhgltUQmNIpe6qbhthBIlidwLxKZ3Xzw0f
arLZujK1XucGQJe7I6ANYHNjuGl6F4qYqWc1a946Al9q042V76rpwU3UJxz1ZHhDKjdgeptwRJyO
KEtcX5QM6dh8WQQ9nIyYswbhLURXy27uTxVWdSv4n7hcJIdAKjxd7UTllhLXBzFOiv5dF4HHH00O
6idKJV5QieYCBp6lmNcI94gKhEaDC6iVRlk6n/xn2DuefRhawG2tb0pWguoDpSclUG7gnpscvyR+
sOHSzdBX21QH78iTUhJj75R2IspZtBsk19LeRAdsC2sUU2pyVt2HsGK8MqpU6nl+5fZOy/H+aU0H
w7KcT471o3I1gDYO8fOKQTX5a3kIrMOdtkaDWwDMlHgebxkkYk2WiDKvup9k2JY0qg6XlUfOZo7O
mSAqyqENTMUcED8cvygi8jmzFbe6MLayKr1zSnAHCbUQbp3rKe0q7y0jgiY69C10Iob9f08J3Tsf
veyfx6NYNVcdNAofN6M2ifrkEJ2j5sitFooq+/aV/1Zt6Ggh+eEo81VrnjtqX/hO1cGK8S/R+fYB
rKBGM6U1IkhVhH8MgOm+8hTx7h6nZKuPDw3RrIWuRldK/ABkeC2obgJIAn+MBVqus/jipUwq69AK
dwFnTpqiG4aQSgBG2yB6QrikeMoKIZEC06TLOA6bNASNGx1HjxvT+zLBdbPiOzznOqRPkCbUp4nn
bEdw2tTS/x8xd3/sn5nlDt+62k1H6lCi3Y0WonF9+hqJcrAZRdFtzPPuP32RWJVS6tz+BFtRxmSx
nodRu/4sCC1d5UBttHUmDG9OXqm07D1iWeeX//xPkiS1bvPrlOHdQNIRZJrEa3ifBOuzx5pBfL8p
cjDjwfAqQgiyJr5aPSPpU5MO5NnB6TjU7s5QzRQC7HB1TPl0zhQ3UkwicMYQ9w4yytL5ehfLMlFl
O8Xb0aIzjvpx6JUpVWsyORmnzScXDpdrY7YRWuzwXJo6Q0NoOgNWq4ADURBGQaocXh9hG2z4qGAy
Tb9JmH2/CiYR+yopIfsWdNOUehyWc8tNmPPOVLPh9sTwRIDAmRCCIc8TJrW2S1fGqV19Isi2SX1z
vCuTb3FUZbloNwqIVJ8wTal5ks0OCiRF+YkJU/6mX8KnsJJMg4GzZpTmSPMcVGof+IJ9qGm96hew
uh4hpURnLH0fLH1Oy7NX8o+ZVnOy9t6iP1101j9UgFo3aDRT+DW9FOtArjPKvpolzRtwFEDmsziY
J0n+GUCFM5/DTIt13pA2vFkfRjSC071zLe8NoVZJGj3owP0yMDKcFU5bZJKRRQSwPqHl4c45bWaa
lr6TPoAFyzn+KTgUAxidKVnkymci2nrphEpPRJg244mcmWLhnRCcDP3bH4uPO4H7dVmrO3A4yfyI
t6TEvrHCB3k5PjatSBKEDzXdCLMFQZMulCjFI75uA8Ouc3V5xjR4b0hruW/eIqBE+GgHs1+igXAw
olYs13F74/WNdwDsq1Cjnpb26JDcJrMW2TKlevaNKcRPwXV4PjLjhnRu9NCHRO1wzq4BulZtM/wz
5U2FqLCCUAB/BTRWJ13bCPIgoM8pKRnA15zlBd/rmVtNgcTUiKUM3KH+4bQxmFeKnV9CPzbB3O1N
h/msizYRCr/KR+ltVTqr28F/AvWagp1xith8e+oClfTYuEAqQxPFsZQ3mW8LR+0NUZGUqwsuHa4j
eq95BgN3ISY54Swmi59L86eHt9i6bNc81nJqGv2aoCHAKdeYrBdZeDgroCoCBgZ1+Ov0JH9G1Hni
QQJMKG1Tu39fFZp0Gu5s2loCVwGkaXnx3Qj/uALOxBq909LdtrmjHMSDzNcwG7gW/Nt8qDa3Cu/t
uyGlNt0QfpSr1KVdnd8Y+ZAn2zBUyNyEpDobXWkAi38H5czKAZOB6QIBE2/+/s/oawES7vobiifR
jMskQD1sBfV1rOBASH7Djf4Ohc6l10TCglRCI+vAw/gzxkowB18JKmAh+q6xOiECJy6VizuMqyfo
g8G/ZOs46rS2Y5ZcnjBhDWpOWFKiGf7jt3qijHti7HRKzWy6p3DnqoqEafc3gxFD43A079gF+VMS
S/vFjlxpuLj5DL3tE5ur+ZSHwL9pskTmEv6PA4nVEUJ3M0bHf/crmIPIT8YRqCP6r3Aag9zzbbWS
DitgW4fUYQAioU3B/Jdd7BmCztpuO0NU/fKwVH7UCmP1pL+iWT5K6A7aFcZ2WPwMIX6jz9oQGZYA
NINCv+Luu3aiur/ISipMHpfkt7HownO0l3TbpcEsIVaTCrj2a404A5jq0IVn/Ox1GfhzlXwQJbOJ
S3VsLfUlSQ9TbBfio9Vy8qBt2weEM6AecT1z5TBHHbSxSCA5DBRfRclValZw9UOWkdWLmpKrRtWo
3VNhssWVoOoIawVoKPygPcL+STPQUhhFWvot0Px0mfr4QRDIVs7ZTmwv7oMbRWpqyiwVZvwFCt8U
G792nWRtw4Cx2tp9orV78A4Eve+UrD7X2PbZ9v+u50uiHdKB+vD8rqnkSCVkEJDESpIWU5j+H1uW
oQCH7n+DcGAOc7CX1XRnn265NA/n0NJxq3JC+B1z4dCiza67C2ycghLhuMqu113C9FMPXApPPq0s
pCHYQAkjptm+GWJ2CUHfLNwHnupi2GAfIHXuV2Jdnyo3RAasDqjf/aNtTMY9UIkQaMzSKqrrgCpG
ZKCr1kqWkY6ucw4zTVGv6wMFs4L43X6E7zPQ399kSoH4wAE9FRxRYSyW/3P0BcXi6c1O3ohber/A
BksfYeie16QjfjI/9UfxTO4mZJMgDqMvfyMqUq5Gf68mR9YhREfzAb+oOTs/eIBFmeWVEcECNkPy
mCdQOycd1slv0SZaE1gch5ttIMlEWHDXCHhiAQekCR/iZYZEtWoYk4qWCYtXfvHu6AqAZTsKHrrN
NqI7aqGdBP0ZMlhiUq+n8d9IoqB0zvgaQDw3WmfYl4yg1HGUfJnO1AEcMklQdBOf2j1lCq8mkjdw
bVixRR21Y0gSnryGz4lKtaW87e1jEW9Tx7ZeJB1YJfbVoETwnBdRiiMmxp8J+VOEOThvT0GT6LOy
B9SXBXr7AS1hDheSq1rJ+v+bnJbCkgwg4cR2R3oGPFiZlccXW2WPPgePhxBUkFQwlm0Y0GTU5f30
X/lC4zGCsz+SeaWU74nXVu/MMsRfmCnMdWLY6zMwLr35jo/6lQ8T7zbXDzxPMAu+RF+r2t81wUou
SOvoYfwFHhkkmXxHJU9X5SiMroI2V/yCxZ8byHpf8RgQGfoFC3gEydnhghbxDs19q0XtVhkWezuc
GjDgCic4e6Tzhozs3RuTC8vKqwFx4YsAEwpEdR9F76CncMX377oPjo1wDsSrXWmM2mDiZvSxv0W3
KPlGzbwY2PDyk+APDza0qOYK1CORo7BvYdqK8HiDCmhHbyVu2s0Z00pHNeQMXJomiIZo+/hM9VmH
MYR9HCzGKyd4XdiAPC5SQCyJsIZYh3ndYS0gYINupN3wPrFte/z43yyNlKNMrAFRtM5/LcKIEJPw
B6/vREhgJBx44Dg/nFKSdnRuQODR9yhgg4qDrFRWTrUh0RhPYgkYfJjGQeBCQHSn4dw1C2HLH1Gy
IO0jYhQMkTt3zKgFaB5L/jg5WXrFtWTYzVoLIKS/d238ISaU0a5JznmBul0w519iImgvK58fzpz/
wkI7/JU1caC3BB2wlzFb0NkVxjrEO8XzDX0n0ihpZiOaXB1WWtUzpsS/CtUoeV5DP51QWJu2ruJM
RtUouEPNePZiUPWl7bruj/SWPmq1GXd69A92mHn9e/nsWHkmf2Q45hqKzYRnkoO68aE9MzIWy8hk
DOtxgk8HB0U9SX15JF4wl2YVpp0DlERYl1CTo+6+2MgSVoSYK18GlA3wGyWns0AihbPMyGZWAniy
tvfJ54MoHAu/EipRw7GPb7lamfi/vXY9tOqQKZgtNzqSNuk4smb+/tbu1yzW5VWDpmTRUF51W3Ke
/mC6kdr1PJxWV8k2RyKtoE+KSUS5jgr3LMiQnDRBsqwpI9F9ggSO6CsECI9/5CYUk16x4TUSFWwG
RYnADum9xyH0r1bBwrIsUylNSlgy+2DFKidRU+TA4TbBQhUD0hBMEU5nd98Q8hevnEWCujLNhl0J
3HqHV6I1PHwVxBhypdr4DR/dxfVM9FdyUaJz6r8K3APVHC/5yGXwg8srYhs0ofFIRKVOXWQgAf0O
AcvOW6UGS4vdia9sqoABBIr/2Ga+b49CI8Qoiu0pZjttm1A09j3CSbFh6tEPwOF1TX3qOAVobUFX
pjdTtYkrnfJ8sI9Vtib1fiDOsHJ1WCe+ju3LY7OAdq5JiBjxqWqAq0hWM58Qg3fFoxcgI4NtSiMD
lHOTzdWeW+CtUm47+hIps5JSHkwjwyLXY/RHu974EBDhB+V/rRfAdbC1WtEkatUNT0l+4s23LOPe
2AxvxuYtg0MVK5/ObkSRtzKgtR5ib0eLEHr2sPFLxGD5ByWchMwAKB0U83Dv6KLHlomno0EWfypR
nYpRpCKkczM9mlf65pwfWLDn/IHHpnjVvzXwDaqoUong9R6Zlat2n0WaFzNmZ77bdIlcHnmZ5dmr
V5IghbSny5s0YskFm9Rqi67Bmxydy5ZB/nQgMCHxiqFRpcrvt/jn8Q6ERfepPp+xC0wVyocuLX+T
RDactkzeTsd0p+yH6nptTy6de6At2/cfaHnK70Nvvj/e5zrqJrfHjaUpCVOA25KLjOqN2vkveewT
KbifZteUDY18KupHu0q6ldEUdf5epzcy7MZ9rH3L2L2VSWR6LhC41d9YTM1ajlA1S/RS7mnWM11w
d1EaDiHh4Ntj+y6lZ4vcDbmnL5/cwWJtMQDvSmBAWJIfxd0IJFTsEvFUdSorw5//h8wfqwIJKftz
t64Bmpbukd64zv2jlnVPYP2Arnz+ceXCYtJCbTzlr9MDJwO1BnRKpm1I4rc3Noz949xFtMGIZjQz
LDU9dYED2fJ1PZ8mwRwpy3VwCry+2cx7w6egcPomJ4wRIhLliDfNk2WcDJv6iHy2n15hWbmiu2p/
iqeEgipDsxK4089t/Pu0HEEfRH45IXJZg4xfyS+bhdjz/uNCivNFlBL/tOGq3icRs68omC3/kOAM
Ft8bNfHoNlHf0EqnZeU4ndmKrxEyLpYQ6pGCEzw7umtJCloAO0QYi9SDynuT09ML6/8X0kZWTiO1
JvlpwmnEMf0EfQo54lmgTQDZ8AwA12/uHEF9Ld88RfPcaVVZbu7UCTDVUng9uoccBksf+Hof7oH7
Cw4d/Muc8WgYctiY9zAqsTWGQAAav3ePqrYpT1YIkgbtf3zcEfhIS0FSMwVPhebFJqVXjEpEPJbY
HxAxouHeTxF0AwjHGPb4BQhu6/kh0BEPaTAvnCzQ7FMuOkI1i2vQ7naR8S7S1kTQpLDQodSJ568C
krboeEBZRQtpOo+F/mIPUpaYXaeBbkKJYLrgfILOi9+1kn/8fYn+/UVb9WzzgK1U4+5kQLoNqlHu
9/6VpG5X9AhIZFWGTA5qBcGvaUluMZOn8tt0nx5anppqufoS+3Q8m3N8/JNbmbt4Kf9P9KQhY05W
tuOwX0XFpRigCqLrm0kh7t8JtZByncizslL2BMGzmOJVm8zUlatHh9rY6IaCKIHSmPBFAXvqlZA1
DBCmaNz+Mnc23FlX5vjkDniFN/Hb9NANlSAnc++X6Rg+Jq0qlLGlWfWA0bt+nK/+uvsn3vCwu54n
yWJFwbAJ1nYJ9jzZM/ObEbGpQvRROZKTH3GOTpYdcTgTAkNP0Og9kRllWpcmlnyF3xtayCiJ4j9K
2qIhQa/jzmzH34TdUTxV6LR9rdzAc/0yRzlqgfP2sYyl893IkG/KUfchKbLx8zyxexY3JLhWpqaf
szosVyrooulfEirI/jBJGbmc6ZvlKDf2js14kDqp7EWgdpHN+TI8Klc3eVYnqXszbCEmH4a4ugBr
DA961ijzoTw26Idsak5uxdeuMhPiwvyQLDxvzocRQDHt1Yw38v8R2GtkuRxQIZyvFuIHoiae4G6f
eMkLOiTCmx/TV7Fg0P1sjyBV5ZAKzZASRQ0+BiWGoP4f0IKqGuvMy8jx+mbsQYX8q2EgqfpvTMUV
dWdDxECtMPXxyXhX0MVbhpy81nJlGV1XF/fcYKcqESgsZ5y0KLgSacevd+SH1cI9QLwHpEpZJyj3
tavYN/Vih/lUYdUnRvOe8K0n/ZqIewiYLRJXRFSwEKZPcAjK5F06K8RkbdV2VGycfZ6h3FKGCudl
/1CtQ1i+Tr8ncmwdEdl7/JMizLrYO2OIIMS841v6NhYepBn0dsi1TqjF9HDAmJ+mxlqdBX3agT69
r+1ijNl3iENkEZUDG1lU9GEiquQnwP3DuUSgj0S0a0oPP+za2F73IqfV27sEo9LTrUpbfCNPG2KY
SW6ttR1aEIKENx2hN5lNNZumZoFd6yCHtwYvCqzzk3QVknMRuRFpFs5ga0n6IRR9QM+TvcTeF10N
s0rPAIifnEi2CaS2UpOFbfvdTtwK0UpNeqYH1/sXGMS7h1Evl4837JiIRS75H6Qyy5bGpgarP9Y3
3Ihau/6rAj/RveY0Q0BP/jHDNfz6m4BZZb6gN2/iFxrF0tmAbVjrQRgar3gL/RS82v6yT2cuifbe
zMbZRyhwL3PsM+FNdPrOsSYrTd9UPV+UtizMRHuqAeeaxBlXsYHetkejRd06uGm7oeBKJ5TNdatk
L3jTOSH1Owz/AbaqwW8DV8D8iWiPasIg5nmiR7706oH1ATtQTNH51DbolQjYbjJIuJZ0cRhnL+4M
1EUxVLQ08AsRwlIMS58vbqjji+Cy7+YmHBmho+HvUKGVUcy7pmcZusrZXs+DrmkcrRF5WAkPqQV5
5GH0cqCAJcZE0BP46ORxtSWjySmwlN1kmJKi9l6Z9v+juVknrI7rThBs02GYht/QLrrxu2222fsc
bGD29N5YHf/omm4u0p+jIvbiNA1jds6q3SDvlzO1S4OeHAeKmu8mmbunAKfVUkBR/xMXboeKOU9k
h/qR5Avo0MPfQGrZlssV8QaC/nyVC69oSfejhDTwwEX/1Qizmuak5ewIoiGvlseJ0JpHWfQ0+jyy
AJy15nXSVIu3Kjn7nZM9WTmyAgUDxNtlIvyt+GrFFd/hOMpNflGwDzV4Io0NKCODheXBU/fMsatR
d9WkuCduMNb8jY64uqfGjVjbrkg3l3Vr0HOof7cUpDoIqg8iWSTsZ2hg3ZoIGs8clqrkeHEa9jk8
yhER7lNvuIgTDceZmS43yC12yD8HafI1OM9RmIbutSDjv9fdVv0eGkHOGuzAuRX4NM2uUOk+hn1Q
OPRpwSlXEFUAfLX2fkasA0YTODuCgoGbpNCb7uNF5JEavJQGTZn8ZsvcUvCiMK055UKdN03DiBFD
JHgJWjXoPYrDzaKDhxkwp+hoLGgUN50nTw1MwSea2UooMyUsbnQ0Joxwy4+rS6HRWGAVHCpQhy0G
Xs7MX5ehifD0UoFon5JutCCa8KOWxdEyCc2OY2RjGk/9VKQzwhH7h47dHA7nRN5wDqm8wW6YeaUz
9QHBL32m/V0iEJiRq88fYNuCU4mtxz1TYGkSqxs//EnqUWcWlsr8sXroPYHPfQKJ5j1rHtd9ieV+
vDE/K7PiUcEkzP+vxI75EgyCPCo5QJKsZ7ap/KMbusLOiTcEd4L4pqsqt6QUe+WcQ7uj9qCSkjL3
V4d04ynp/1q8nkjwFl6pdWXNjt2XkC5oR9cZ7dTvn96+KmCsasgOmQec1ssUTqv6R3p0ooBE6RpF
qHITLFff4wWezWOYcWWEpxgwtqDglIuios9tpjhgNu4LdBFhiNx4J22OSXIhnAHRUcjtpjojOGBs
0ccTQtqth1TZz75U01QdR78P5QfUxxDCzbmbDqsob7C5rt21xmyCXcoimqh90MCcwcbglqqhzZEE
itRt0+YeXkBb6jtpviVJ7qhi9p8K8pv6U1T/y08kjWjLabtxx4qWV59tQ3GJ8jFlIvI4NYy5O20w
Tmsa8tPm9Oa+QulcqNoROHrJGdyg17QTauxUAbS+qYuX+YqayooqwzcESlay4AUsqDnzkgqKKQQV
S05pN4YRpP4l6v3HbMFiAY/aNdJhEza2HWGoHICD4ygR9U/TS8zPt26EE+8qWCntvsLqRikHpk9H
EspxPjCq7EcvFRoP+vot18+D7IBRUL0aM8CLGTZUZmM/Vt1svlVCfdKW+XTNun/SOKXi8nTZ0ONb
eyfdq4oHF11Jz4FvUu5BkzDUhaRs0VtDO/wy7JLBRVJRLoEVDsaIkPizdyFK6XwmQV8s9OI320vn
xSrNcUGaTPnHguYFgha19e4xxdoAT9Hqkii/Ma0fdmCt5iwLCiLTmbsRPeqzGI5PPM3NCEC60WR0
rR7pIozVvvYMToqTGMyv7tvSLkJhZD3Ue4Cvk4C2NEVCj7FZkk1asgjSVVuJSirmHlW1NB5sQwpu
/4J6VOsBtLpCySzU0r1VkfoHgb7td6YhlgWEcS7BTZeQzyqM58PPKuClcbISqL7JfSrQJRuQ3QAv
5TcyJny+p99xhuEHV9ogdMUpAfFIwppDiNlqvET21lFaNWGNp5LAVALLQcrP+6ryMlbTHmAhw1ZG
qjlQ8spAi5YNDod7HUO/kwEoX/ukWC4HHZxUvdWrEVeWxwJnEFxK/BVfajAb7gTC4krqMJVNHRrh
0t7HNKuRYQh4GKv5KCCCTYAfVrW544qxzouJQkkau3WB2AEsuFm8ZfI04r1mSZYhykodgGTHjFh8
r9/Smf6E7/unytQ5lCzuv7hosrwiebJX69wosgNhljDNDTa9kXUtIb1Xyj+fNayrefMQhWDes/XC
v7ataAkthV0R4R5UNofiu+qsSdi0qeR5PmJhqoD3U7a3UvjftyTBc3zhpendVKnEj98KsRn7OHrD
wAkhLrBLlptuq8ViS558RQybneR2GXXJHBt5+fhyPAJRGA3t9lK02XIKTTRCZse4Lke+10AAMtEb
S2zJPR07MHBoE+8Lykz3oZPsuzzv02EoJkhSXTFOzfvpPx1nb6xGvlPJZLCTKmhjCMCdTUdmE6uf
kjRpK8DDst3rHWBMZPZPjvAwebNXu+VRc6KvOB22fNeF52/eLSvi2lySw7lKjScLl/8CDJ7L1t3M
vEgJ4yXDKAd87dL7+fqS4gh4sU6k2Ifs0NgmV2H9gcyiydxgDX6HB6RvsJbqRWLUQj6Twp1E69A0
UlGtqAZARQeut0imw5VA0ugYTFcfvLHFEl1HYd3+l2SdpgjIDAy/CrcEK0+mUV0KjiJaFi8DIlgg
5iEY05uhJ0gcpZC9xHkbqACCo+BM9hEEc/ks+FIC4K1ukANROsoIdQ8tAgOhNTTWRCkdUT6NnLR2
5/QHyb35K5JjzYBKN9HOuYmwTDLKEJg49PnK7Esq0m6r7pyeEgR2aJovE/Pyi6UoBTxGRtTQC/Xv
T0E8ywpLnPIGVLdEw/kxFtx91g0q+eH0fZ10uxSsuiF6DJjbMmnbVlhGZto4APOBFyHa5mvSXmw6
mn19e4z2tOzRaeYhbVFOSzZ2ZwgABikaPHduAbvD/c8wnQxdrYUZAZrCNYpXYyX21qrNbpZaD5ay
ojeQ+8aJNum4GzhnF3Qw5v16JWgfdTt6wxRbjR0JSigjzZZWU2062xn5nzNrvvQMacqyhbOyysAE
Uty7lmmRyhOSlwEq1I89a1jgd1j2j2OO6zbB/8rB5gs4dAPubHLnnuGlFamVFmURV/81z8DNumdC
LEyp9hZqImcFcvT5xQLPS+lXxCtDn2k1V0y3MYJ29PMzte2kldG/oA/0Y07TYQbAkC5R2c9jRa3A
AoK9omQmVeE/BiCapJvP+bSpTV4Zj1c51eo5h1EsjAoMm3GndTlTqAn3468HZ7vV0ROYZ/GNaXGS
OuygqCA9I0fjOJR/pR1Eg6TMW59DHKbLUdI1gFXtj45uaHDLZ/YQIIk36BL5ngzHwpIwqPxApfgL
1g6UBqZ/LHCW1gHXXyHJGZHzG4DbFCkLa29QTuxq9A6WQIcbqy6I3VLigSZfw+jgy7WrO4+gqjcF
rtwwb1ACkxBPT1erwTYwL9QLK++NLV0gMqUk3rKTBTBXewnPJy0MhMMVaj4JKDP1OH0NSxHLTlZj
Be2kPhaOKsLh/KbPcL5K/zXT/xZpdjRmjkO1ylZzEjYDSQqZpeIfkQds66GivtHm5NzwlubVuX3H
QMV8HVHz1M9l34lPs7KOIY9SBdl0vGheEWMFA1em3FblEXWT7tcysFCUx8i8KdWYt7ES7O1I0oAW
Z8c0n6IRz/ZOBukyS32nQPb0fBJtXddSD9etSJwmLBpX3KBcqamoKU+6+5xTZW58KNsD2YL0LHfA
rOM6VdJrPxv1Vb4YkO4pJmL8EV66lnnfq/WJh+LaSoaA9qzqxBrAAij/OPS8sKWCL8UFF0yFQpEV
jDdlBsZUKdEaumLwMS/0TAlfzXEe4cflTWpa+gMOX+4XSqYG6sCg2KdF8anYKKEPYnppmsfSoj3K
Etz/BOEbd5SWFMZWY2ToHRc6DZ6mEcPSMq6SUnCxgsQhkNQsoXYwNEINBm8Qz0wEZM2NSwiPLzB1
EggWm3jVudYKlJqE2FNpNBMnXFMKEZTeJNBDBrUkyj/MMXa3lFLZOyG2O9XTGkP8CruHDjOuTFz+
rLyjHKCQ7ui2vjNEWnRoiOqo9KNc+yaTkN8lzQ1lAyFaIS2mEXwVNvQl4gv9mp8widvKyMK9ut6R
g7a8gUW5uOq9Htgaes7fwLJQ7PZ2mNM7RAP922C5jS4wtOu6dRaq+oD+akkKEN37qRhO9yMZ5tIS
x6bUCWZ2Uu+8AcFo3oWH3X593uhe+c15uemDTtnblWuqBFwcVofd2/3qcN46HQ2Y7tSvE70sDQgq
eYC90JM/pww3bJuGk1q0K8YuwQuzf7ZTKK2wL19w7l0aaAoSblqIsgpYqzv/+xP8Na8RCr+CE5WT
WUtkpHD+qkCOU7DDZuRmoVG88vzmk3/R7RK/wXNSk2ZJZgsgLuGr9IuqrtuG9Bjd/k07Y17u7gIT
wEPcKLTg5K4f2gfxiwBI5ELDwE9T//9uL3GHkzlQPm6YIrMWkqlV0PIDIKPVKy6T2v2mTvzrlvEB
v2ZNmAvr1bzauc5cFiVyuf4yXm+gYfhtrg+3JAfg5C4cT+mhAUP+o8IUmw+ZyfgwLo3IZDxuv0je
nGadry3qBISKVIhz7QPHnGtufo0WCMc8gC0hyO1NtElEQqTAiHEdpNQeFoJAqqW9w2saYiyrVdrW
GV9UKyH1Yuhzqmtm3KGP4cd1zSTiniuS1EtLuS51vkY216zrs7uxxshczl52y2SRSeNXlSK9hSPT
BFzmWbh+nepBdNm2WwSiOv062jRTWMSAf/tVpxx9UPkRAHmOEa5Ht5H6KK91j3OLknlB6M4nAAv9
Ow+R5fQ+7bvxI/eJym7Qq31ckOm6bOuVMBPKepWcvZ0kjpOd15ZQw0J7vnS8xgcr0UOdYpVCQD/B
JKGqWKNOBS/8PsVZ9y0Lcux34skxhUgXDDJcEOpDzapr/VB5nBnWOme94Sa8z7jvPgjm/4ir3+A4
BoGMrtODAVDTuoQEFdc2jfApLOiCtTfKuV4QfBkhJiyVwM9pJjan1zkriRvn4k7BcEUlfRln0CUF
EVbLzGJ8NWn9ZGJZnFa5o0EPNsZ6EQbGOsmPRQSG4LN945CElkytyVOyNAJ9UaZb3BGYAHUNQW1j
JXBGEIT/agfGT6hpJWiT9IGDBZpyLx2anqpcpaO0yCtS2JvVrrAI9hQfwLsPg/5U4CPdBJ8f24C4
0I29+7hslUmwXToPk7WApjpiUomlFsEwoMDthP1TK1gVWzC3aazNKrkMrYMHA1GvASwIxh4VnUjO
yWMWTL+EV8ZZ03OBPun5McVavFupWYA4f4ChM6HG8G5hF6ymnUjdgX4g5jBzH0uudmvMC9iziqBq
sRCcRzELQJz2ibDme8M4B+6Z+6P/2+NKUte5tNbVNv0KI8J4cA2PANwxQrib00vDTRIkHLyFODwD
RtyMWcivpxLhEiCACY1WCycT/NeAUmWsxBpelB8JhgH/sJ2ciYBUQVpiRk0NeG/U0LyZ+YNRbVTC
9ns3jdVcG/IVUUw/bRwFHDnvHytw1LqMTf0GOOEGxagZ0JkE4mGt7NLaH+SDV4qFv75xHLCCTnH/
6GUNHekcfm9z2vsNNjKGFTg+8rbmSzHf+Oec2kImdZOg8ElXOEADqfNXvqCPwN2s3hfdVHxACFce
U/ceJpYrE960eT+OR5ak9+DyauEArIgp/OVvVep8I5Ei1CzaKYJToH0OkUwOxxqp9u5NcGATC+R0
rDvicZ/pN1/QFEvd3xkqJJH+m0AT2gTV9Yg4CH1ccEMRJW96TSt5sTJZTGfVm44QsBWmo8seMcCv
pjz/oeu7o0uNUPHMY0QiDg1shkCDWMZS2YZE44zVMdZlVfj1YF2YdxksZzYFpIGdVsdJGPsXM0NS
9Kacr3JOPQ533k8b1M0UCjsLs9AzYQ97e5z4+8gtxRxkihZHUO1hObaLZ9pgBzwI9iVkofy4bbKi
Kp3WnlqNpESqfcLcBqTO+bBPETcgT79rgqeYy4U6OyN4FTkzQSf67dG++Yi3C0QQEqrB5vas0raU
Zl3hMWrVjFWYy/tW1LFM0nHJH2djmr77D3wt+2DuEAcTXtNHgyf33qoLDIWQWANIc5TWAHhWG13t
eAueF1ZQqRIK0drkGwic4mo9ari6k09loZWnkTIO3bb62WOUIjOPEGqb3OLbm2fYhbs6Ia3qsusB
TxHGJhYMeCJ0X3POfcZwnL6yhXXq0Y59/MBMJgWroiNx6KUVGq8fIh4ULkSYpO5mrCUf45kkL5PJ
XQ0ky9MF7Oj11hYa/YG4TH2mW9LREm1MEbwaIBNTYNz9xTBryDuW59RzV40xTjISc499aeTASNc3
Ri7aR+9sjKQ2DJAh1rnFsUFNa7OIbjjA6DK/V0OdXokCI234U2CVGa8qjQd6yOkW8zY209gFUT5q
jAQ/g9jgLrbqIJrR3h5xDKKS4na/uQFSt6tnbgr0IB/q2pktCCEiuCmvkrth6I5JhMs8EJ5017f/
rIpt7cNKKmIpdKTBq7Wi6h+cM29tpVFcaD49NzvSjaPuwam+sB22AC4JhWyZjUWwv/QX+Yxx++Be
OvBVoX8771LRZZADfYU/jm2m8PX9rEWF9s2tGDOmCoP4UELSIY34yVxlgss1EoUHv/wXgf5NELqp
Ep8vlzqAlfyp2a+0O/Chj5y7I+FY6EOnDdziCPHjIOUWzDci6xEE3ZejvdTjK5FltTorgNICaxIG
7r+YwH/R1sZsdyESp6mYIuYLH1q+ZBbPETF3muTzw8bpHeC39TFZ2csO59XYtkRM+zT+0qDYoIdV
nGnH9lWTeYFjAwO9VTl7XiUd6eYjG2Fm4yDmYpccIhIAM6yd0rI428vpnez16jygzEapnym5Skfu
BSRYHlnB30+RKllksPkTvsJDFsx5zhsl7XmVoIFPBVuoTXXd9cKjuG5i8u4vf4Z9usCfL5yRmtT9
qyQUSGK+WRt7CZrWPQs//z1cJ+rF0YlWchM+SsX4Hbvg7lzyMHsw3sZfwVYGBhHw5S79xmb7YZrv
q9TzXlW/NlMYf/8gZNS+7x44yCcRq/r9IB/sqjWjvw3alCdNSS7FYDZsdk07Vx3tGko/OCvPFx+M
BSq4aYsILxJ1+lrZpvyVDh01snE5W6408G9C+6cfNxOzkAqPWaOFKiOPw4cDs3REVKXrgt4r1JyF
mgjn0u2gL/rLx7wQ2SW4UYOVt9ra61y1ILLjCEfeJX2xVKjJ6rp9lWGLHt86xwbAs8oKJ0DydDB3
JqZka6rv+yl+U5oKlkyP1LUxyTYsKqEFjc4k4dpRhMzKSvgtq/TiOYQWGihvyE1g6egA4HVn4doD
K2SADfeY4UyDVyqWTolVwUlOuMQQ9lCtEncPtA35iWdnUdnCAK91vhSBfQxz7G/sef9uKCEqE51e
pXWVNqC/PkQAY3EZy55+C/Hcmeukfjf6ZeC7YcqUmo35VarMjyB4ivu6a3Y9WEgGPUK2USoGwKws
uUl9nLpPHFYROROXIRRqUrIRs57OQgp+7H0YemQmno7ewpg49jaKdCz0G0xcSmW8fBg4RL00P6p3
MVjEvvo2ipjb2dMehua/AOa/Zy7emhQLOzTG9BQtUKQhjweL0AMxCqyvbd4a+oVI+boJF0mld+Hu
kyKM+Vxq/Id7cIhagGoyzTkGlVDEIK2RXen+BBoaAurrZiGZC23Qy+CXV27sQo11weqemfH26bvv
0nouETv+x6J+eJDxA0zXS7JQUlxNkGe0I9h7h0gliU+2agGxI/EZ6spvwW5/j66bSdrzWTSsHzHP
ewskd1R4o9PZw9RgTxDwCRjIiPVRfmF+IZ8QhaVGBF94bfPvlcF+BTRTgpMS95U453UNr0KfJwli
EbJiuypnQEWUJRvyusAvn0Zqj9kzMWV3YNmOVklaq+QYMdBvcKmgIcTL6EmcbEbge9IRj6bJuwY1
bX8n2itOfEeHA7DLD69OaMpFVc7Jt5ZP3+LTetFhr4cRsRP70g0cJe6naZAlxMQmCqwiY59qHA27
8pL4LsrWCJhUofleUAsZpVWlulp7tjry02YMLawhYXdLYFBaXMqkuV5psfAuxPOaQsk6yimDYZPd
vUKoCx6FYqlI8N5SfmYKZm1NW4oViKaLDnKtzCTGOSjfADvhNN8ONuOTtGibIiCj1qAVWqsffFhm
CrC1J4bMLCDTA2SkpxfeaLMW60ObPTELTvMWV3Gwf8G7sO4jqCZ+F0/KnQw24qidcCUBIodJTTFk
M9lMgsKB2oWcA4tnopkMtPX7Z0dpmjc9SEK78OBXpeQZdENX65/I+Yc0/YaoLQ83SVjyoFWe7W5D
CQF5LHN1O7mm5rPXNf+E7f2+9cC4xsQbJeIk1Ie2GcnssvMKWgh5SUbpJtfNg1dmdGX9swOZMbLX
YkkoWpIcvrToMFHEqImjBlJiXdozkk/m7PnXSHl3N+2s6/nF/5wvBLNJxSJa8lM1juWzzxuDrnZX
Qz60dVNzTbmDGlhiWXDgGZ7S7Zu169XTdOEmmBvNc2SAJkEBrGMYQHUWQkVnPnFeRVPn7DstoWeY
+ajU0ICv4Lnpy163CDInQjjjPQFdkzIRrkaw3iRDAtl2+52vmj/4S1DMq8Tl0ZaPgUOBB4nQNwMN
ieuNpMinhdu8dnIXUZGViDdueTwpBlNXyhr1DD11nVAzSLy/B1izGJ9sZ5xp8vV5gt6oAF93jOIN
le9g9md+ET+bs6o1e+N3LGdE7grF2I/YfchLRo6IWFWpzE03FSXzavsiUVlPSXLRVbPBzpbnYWZi
vIBUKhRXV8Xvel0g17Kk3KThuvDl/OgKWICjCHhOzh5C0D49kdZjg41P3jsi0TNnKndQMVT4vaJs
BdExuJZluHBE5p9nVONb7yQbrKHkzV/+7KyEpb1iAVAB/Xv41QztNPzHOeMTNLNg/srvVB2jFveP
w7xGZ40F0IjszR0j3ksi50zkW+bNYh354O29hdBTgJmnmnZfswCzDf1QNoMUf1lzLj+ZqvYynLZz
6OQKs07Iyeqt0sahEiZK8NocCixTXPPRowsUlEFikxkcyZCaf6DevKNCOZFwhOxzOV1jdyUvsl6n
ODuP6yUV7v7gPr1zw3lior3pi1Xgz2As5B66GfLGd+2rgEH3iYvFQyFf9+zG7m+n0cx13tnMP0Ei
v2gzrsWs+mgj21GmLRCix9eSmIWr8BgtzuS2wpxtuv9JBkFzhl/t0zi5PHhxUcnrsI9y0Myrde7N
1MtDqhe63nTQT1709R8WkxopQCLpb2Rt8HWv6PxEzGQTq/pRv8E3WmCctXOW1e7h54TtQjh16LK+
1ax+MOGGZVpzaq47qZnOhpI+epBtb3d96J4RQ7648+rqkkA3n6LPz0Uj/atjs8PgtcA72zahVUyc
UUDf/fW8wepHsl/vdCFlUz6Y8gzZAvztmJnlfwemvJ1jQHgA7fWHFs9ekzNcS/q25pnS+MRTOsNV
wW/0JCtrJrMdAimdh3MlaspyejeDET8/s3Ho4JcKiJRMBoajx5/CsmSvKxXLBOylT1ZpL0cZkKgq
IbQUyvlWkNDCfzCC69xthfdE++mBwaSFYskcNCq4yoCaN5xyNrZZFcwiVmxYJtaxSSZElkkHb8bG
jeZHsysZdcDgk7P/MdubUZS5pao3DUf7lae/5+OeZ98tLUnBy6WXHsQMxOJ9flF6xb4WzYkLSoNm
WIZEfbaGbQZPsiuvB/lfOInSGQS7zurUSZLn5yRaPG1bztg/m/uXb17/xriT+3hkglbUebTQgIM7
5JvWgFM4Go9xWMEVk2SvQYTgmKIYrMXlUejVEnLQyYSJAkAjKYo+DqdZg8cw8GLgWslz8hUhrS89
j3y24/AunLmT98w8WhpZvhnAHvZMRZzMJ+m3MxP2qpAF/y9mMQsvz9nfElaIqrth+ANzXTIYimKr
tlO1xa9AaBtFX9a5hvdToIFFtAjr4/1MfdVVyfujkhQRVL87AwdvClMPlN+59Vps0yDKmqs0RVNv
bYbrNNzTiHdEuI4bzHvCZT30GlGC8nlUz+HQzRg1SKcxYh0wDvNd1yzmxb5w+CqJCMYviRxyqsaZ
AUILAKiPZVuqApG8+aZmkJC2U19S7MoixTOztrs1c6u47e/oJ+K96aLe3H0pX0kTMNYd7Af4tgmZ
orXYM2FzqmkNetnRUlvz2Jh5lNA8vb1GS6/xrJvNRjvGlm10m+2f2BFsobeW4SXjkv8xB7hr4/Ix
Qf7ogK7ZFmznc0oi+i7C0kH6tmJ1aeeWucjk8BhwGLGdcqL4OjUgLf8Dg9HP6afXCI9ub39djj+7
DPIkvL+qTCdbUybWT72TTryUKJjymShnrmVXXdEFw8bvdqDg4vKAywoaqkpFijbD2juZsWz0lD3K
9hyOnULr/6+Cfnnay8qXgQnqitYQExCpmWnmh3eYOjYi8o6Ja2phym6I3KGS/KNpKQTQlTSV9zqR
szJ6knwvQkniXn4+nABKwKUTtGqgVk1GpMWaQQQm1MXG/cn30gpcxU2AaT7xHRuK9/qEg6VC507V
LNnGsXQ/I/JZTAox30GGgILHabVB2E37XpG5fVsJ+Ss+lULtFcKy8AJ3cgRgm988zOG4xAIPK2Mo
hl8P9FUWDezsap2+z3/SNrJo58KoNk7IkyoDsQpcliT1h+87ypcbXbkTPlgrDqkDyim4YjUeG97l
DWBFanKwR3+GEaACnNrYhLKinX4wS8zO5sziGn4Ckwvw1RbkPreMU+7Z1nSx9xBHw28AXcMbwWs2
oiMqOVTTTmZE1u5oxnZBKm9k/6Cvf5cTINP7Se27dREMlOncSvx3D4P62N5YMtJPerlVfDeqA949
JlT4juidfn7KOwukKQYJEWIxeNkPfRaNVWHaz0QLu8I6m6Ikt3gmUvBQ3Of6XpvX+BFAmHRsSNuy
SMr69u/c/yYjRwuFu99HqGqOMc/ZXs2S+Rr6/LLvRtuCn/vBQz8mjePCYrHyJUmz22gNe9rrLlbu
ANMFxn0FBNAAvS2BAHYCNKldTLuHrY6Gdx/ispg85KCYVb/nYatqREL7dk5+xAX0yh5Ol8SRqX83
yIerWyOlOXCHksAjMGQOFDNvBz+obj9Oimy+CSs1vagGhtkyoKGwHpMYdCRNafM3vkvL0B75uz0A
FANtuutQmXHKnIsEaX8DTttcghF/SRmW7Gupf7DawBEylKyTNVijZb5X/raXI9uFWu6ZNWL5x4wy
Mb5b4AETNaOoM6m2AhgctEasDLA5M4e2BNrkPNhG8WIZQ56eL9IByLuFWABi9LOo+8jQSs81KwpA
vOkQVHBWpnqAPsW8Atio8DoftKiL1TGPCLmer62Pv4gwyrffXhb8+wQ7ILri3ME1hyJhLeTYkEeH
9UDV0Fa83imoDrnWOHcfdbwEWFNCn2BM6mfoLw2VVFofqY/6d8ydd6TOTuODwAVz+PJ2qiVWM67b
9B+Gls2u8M7NlwxSe96Ur+ToqgPyuk+briZ1V1QFKaqzNsnkpdD1txdX4FnGxXmeLfZO0ujfHyH3
peWu+Z1JLNkHIWChxjvf+TMlIrOI+r+d9JR6yWHCjZPtI/juMPFXSB6g6H3rlI9vHnwLUIer8RtJ
suCTulDXB53IC2b6aSye/S/p8grVqQhhoDl15Vb1Pvs6vLshwlz/kQOIW4ndWO7ASpLHsrsek0KO
VWjLj0TSwVOeaXA/riw2QHKGoErdCAUlAOdWa2W2R0Ufv3WEmMkaElOTx1lk0tt/ImyEnRpaozJl
GlRqydmYlzDfw0oLwgOx9696eNR2l5FcwXIw0oc8xmf/f3j9GGCrR2F1AXH3ncW6iLWBqYpQFazF
oU7+/eBkni7U3AAMtwifKfjIqw7edcV6BuvzT5aI6S6J12ak5u4aXLq9c7W7EbH5yc7Dp1iFrQEN
boFfDnBGUs2xZP9puV6bWe1vmNC/sRPrvq8tduemgfTbnvxFoZAM4bAOF4XjzD5BynGxzpDoL0Db
9v0+hi377m01Y1HT89VT/EwnaiEZxWtwVzIqIr09Pr14zRJsTWrLD+Lzs55zTao3SJJjB8eh329j
SC1j6lfUCba0POneicKQIsP21TXWCCcoVhVMWBG2ex4IAg0VSS1FQZoQMutd+z4bPi7w7hlGOYQL
/NL+wVDGv+bfJJxNvM//+W3wEjiV8s0nBOpiMITHR6u12TcgadxbQBJRBtNcc57t37LFwbs/jWx1
tFOynStliZE7AxMv9/BgHeJDIXoDu4pOpWRrX3pn4aLnmOk0q4u113EwCRn2sTJSQDl/Q42vdqnR
ULy/Jflz6M7g9O5TDm90FhV6a51e1HJQ7HkjAPBca/o7+cMAchb1G7Jg7vUhKH6I+aujEl+rIT7H
wFdyFrry7+cYaeDP+PE2c2Cm24MJJ/2a7t6cg380xTTj45djb+KOQfJnwSbSshqZLeShgqnct35k
SyRyhzcEA2VnhQhRNb4q7RoU+zIraZwd4w2zojYuwM4CvFw9AHyVwJoz6ZcPZAKpFofBC9D8Jufd
N2+53pSVzIkCgYUteirCC7f0KS9VYoFtvdCZG7L4duW5TMAJUfW0gDf4r4mV4Jvhbcgg5eb7JZXW
4SFRYDDwkrfhIgseK4SqARL8Wn35b/GmbSzba6PcHyNoYUrYiqLt8awiz2Hed63OXm//a5vm6fJT
5sC1EHYiLfRTc26SXFCxOCP9r8MqZL7f8SDwnZi5rtmC5kvE+CM4tPaWqcVP0DKW0MGcjucRBZ2v
i9dEJ3MF+OuexPpR4mObj4MyOAq8Eh7y4AlHb4i1RqEik7Mnseg+6VwNWSqepcRVCZODhWA8cpcM
YLh9V67bs8DIiHnlzXHpGpIS4Ze6p/ZnB7E/6O8QfxlGW4YtwebJLrNOLOOsCuRURMCFwgfwdMMn
XTk+ERRtu+EqBgkHI/LVuofCopsU44pS9wMDuyNHUbSoAEP9PafPLgHATe+b7RKdatjau4QrzZMS
FXI6rC03gDKQSmYaSWXH680J2JleurX25vnXpYxw5lJezYQ4ggxPwkvvsDSXGdq70Sw6ho8S/WoA
RG3PpylJn+Bdo4gtSpFgdjahpGrjLQ/LsAC6MwqnhWX1GICrR/Mz7ahUl+nviWT7ly8uipEC/AKb
zjRdXBxJFy8yXteUTAhODPzhhXOAqBtC3DX9NKAd68kFh8LxpywfNjwAqxnIkZSBX2M8oPC0jx+b
ewe6A/zxVT9glLaU/nj6WrnBE/UPhjdvqH4Q0090mOdFbDit9H2oltL7hVNUdspYTlIaEDY08tlT
kaUbqkcmjd2rGbTxTbPUTTgz+8AwDSATBMiT4/QDwi43HUi1d56w6kYlGSah3b1I2PyYu7fR01fI
Lv1cpkE5W46+YaToPdMGRDWUAUIXrpAcNz0l81OfvxCC5b1QHRp2ZXcC+HVjf8Bvn8kBJUNv9weR
4ogzMP/R7EAjoxmR3L38XuVcD0OpXiiORoUicxmU+1PLHsLfHYOIgoOAPfqQ09fondr38cjlEo8t
iXASRS6yj6KSC3otQoEJnFxd8gnyY5QS+4OOzhKOgfRWlxMjLKuzlj5v9vZqzhWqr6DUZGMcY2Gt
acau9aB3lUd/rGuL/30KhowDFI9rM3dHPZ40SH0Ikusi722JUH7R90qoH1mgg0YiTmYtAPzqwcQ9
et7TSH54KjBbltj9ZDU8UsDDKTPbhWXZHkmD64+1eSWrBydktZc/v37JfrQ3g3QNews5MchjMEju
XQOcxvOIE0PbZq5ENr67oSSrmKy6v93quJCYGJGvQ+SlnDiW4EiB2ng0XNV2oadq5CrEMxsO/sRe
7ej6FvZKPpZIvSoOqlJCIJwW+ZOCRVv5+YHuP8A38N+wdIDj19wPMisi7a2znNGiMFS50mVnexnJ
J4JVat0oa97Xnt+BpDkj2CJJTzGncjTZvq2GFfdZbRnIUZ30QIRy2Epo/rPrN2IJOTbemp7jdiiD
vvlg39pA3Bp6CXxAZfk2OYxikscWX1rxrSyUXVfdVRuLL4no62DFuzUTB2W1UHJI/kdfBsP3gd4d
nkit8C1vgYkJFnP5HB/DGUVxx/KDqw9ke0igv6Yx7Kvpy4dHpgAN2Gcfw8jtjdHSlMEfKZoUBx8i
FZpGUijNnvoBTXD3xuIRAl9Qcrv03SPBRqEiqmc5ZZDc1lwEeiJmC0xUAlV9BA+jYQTBUT5PQ8iw
xPa4BEY3qL7k7AwDe2soy6e/XUW4yibQNYxxIa41a4+wXVwqqRTwoasPiT5FGJEd2xch7HmOYpOS
iSwoCHBHWEuy9SF0fPEHApGy3W2zCCHfjPQ/IQGfCVoQKNp3gll/NJ1IHyWgdE2wHBy9cRM158fb
KYHLWbuwnwvmFv+T4Cfw4V6JTL9Y8UekgL1VKUuf2O9sNe977F/bJXtTkoi8xO6nxohirRowLRKE
p1N0btvDbFKfmc+N3aa9Ge5VfRKXwNbuAIvcMaDROtEjpAdQ+PeQwHlboKrS5JXb+00yzOdlxYTe
xnUUojrfyBhuQNCkVzocZSiFC4QVYVf4Dki27w/RMZ8TGFgksiDp4rZs+vEv6jqVX0j5ydOmo/va
qZ0bbJKsKjB+cMDLyiTnlhD7yOJA9dwaiHrVKiG+Wczj7wPNMzUzjYnBtylpDczgtBd+AHFrMitp
YQI7FNfEvAQx+iYyzQ4S1MfwUU1fQ14allKowZ41MMTPH52Wxk1pVPdH9CN3PzKFQF7pdV5j4E3z
TQ4M/Z58nQyLCSaTYMAHivn16/Cbn3tNt6SQggKFgg6ncT9Mt/FqVbfRyVWK2Dpc0nNXbhXfqQPP
gRdCEY89/aqAGPOWx+s2n0FpH6FvaH/3AHFwRFJMaR95GAUC4jgGslWtgUVjXt55bb8y0iJwIHgk
vpwPIYH4Hra2HvNSudnZ9Sg/UF07UedqsW8XsHf57GOw4AJX25bzDkHc4DUo7058xSVRD0pgdvfe
49TDZwbWjQHo4/bhRiql6dDH08ZmkkqMac5HBCZoZIMdEaOiWxa7LSsDVLomgBragXUY4FGKQKPB
kgcqAx2ZxmWcMC8UGDf9+6jeP/++/aI+ZloK99/6tRMyud3zRlPO9IonHKxq9bhFGrdQBDNIaRtj
nUHYcXvvJJdlszrKCmhOTld2IKwGJZP094Acu9GKlG9UHryzLdJc/tdI2ySarbPJR5bZb/CzWRZI
l5romoFR7H6BeSkV1yezDxaaJY+7+iF2YA3KMAEvRJ7o5sM/+4qBQ+PBL/mSaMxpumqhia6jc5OV
zD7/FnFuHJ7GBsSRDowVNvmJTs6a/QSWqpdoVkUGpA7l1ToS2pPwe8g5gyTvT+uYuntChee0tRkU
c5pNgxqIlrMRVbKjBppUvrm9XnmjiqYOcQg90WPc5/X4JP/Hxft5+icIlGXVprr0/f6LFJ9AZVww
LE8nV6webSNU1WpIQhnu5Jxdu0DzZHqJZc6MJuYtCv1OVCRby+5UUgFRNkArSsBXtVgI1ax/d9L9
pf/rwW6GbfOeLILE4reYxxJ5uZvFdS3O0HScoIWchnFM036qNu8W7PlBYNZxjSh0jntnrRAXgdnC
VybKhG3XL/r5I+XAc8RPbnXuBG4L1gIUCefGN3K9GYOo5xONys6BKB4OTKoTn0U5iczdKeQgwn8u
y1LNED+33qeUVJe8oH6jjqqhQge+ku1LkbpdoG0h3I5rxzzcl88r6Eic30TJwfBNHwc+Szi+Qwkk
AXBtY+htMCi66zloj2qJC71Vgb8tBocStPWzzMftsujJDZmIqTVzL8SIaycc7iimOdDygIFSMWj9
MyOGUCcoTtHt3p2kuhyxCKG/MW4rdXatX5mrTtn4DYAFwLbWoLmAxTplpxKf66tOD7hxVXbNdrko
27++Sjdo8bBindLzE3EU5AuBozcPkgZCWEXpzJHVTxxY3fc058vJUBGOkuqpRSWn/tn5sLEt5Xxo
GMeJXj5ZvxGV6gNqlrxbQSKt+N5ldA/xRQ6ssHHLftQY29U6ZaT1Cl+I3wL/AILGtTodnIfCkVKK
XqlJv/mxnFFuin249p4B3X9XlPYcMzfcZhpdZ+nsgHPYr2xk1FsgwJDbfYi/a3x0bcpEwdBqO2zq
brUErjdlF3ms6Q1AgoyVIxiYG6HTskgZQziWX26CEfYk+0Ixn/4o5HhkB8ASwxTgX2MODN1jgHyp
iC9tDjzKu3gAOPYjk0QvBZfXBLrv16uu6X+5VhUfgZj2LWFyXHek/MxONMJlN8rK+oJMNHFk75/v
5gEx1Y0T3EfKnZJs6pR16lNDp+n7Mn6Bf8iMCJKMuU1wb9SAndSJ8NUNIVjedE0MifuDzbOa+RuN
I7auRj/JTlfEqNuCh6pQ1fXjuAt1PaAHOi98VjxYZN1979ldxUkla4+HR51E5pEOTbHJMBaIafbS
g57Thqu+TgQPZw7qI3sRI/zWH0MDawjFxX+3jvX5uYUVcSyfVbWXUrBfOE246l75wp8NAcSBAbni
7Iv5433RL1FjfZLcyO0ryHK2YF1DQgQ6XQ5+NYNQud3KapSeIdwgkBncEGI61FQskS0V5z2xsaRP
CewQVPP96Q1qblGWqE+KPssAGSPUluPr5q6mIIxIWarAGTxAqgEEPMho7kenQIlgMtykiKy0Ixrr
0vaKsNyfzk6ZWIiNb5/3UuRMXNiv/kMIZcJ2qi+4b3XGhMnyRsUkH0WAx4vCXhTXMYOm4I57FUvj
XHpEfhxlIaThn5vCTXVKHJvuYORrVb5RvZvluzBsVGv8MZGIQgrhHe5yVMrlQ7sr2/lU/9+LfWyN
FjZ052dX/JX3v8Ja1B63geResmhLx+5eYdCsidU/6nS6l+mexq1crGx2tBm5UanJLO3sL2G+jYQ+
IyME1eMvPiPJ+9G7Zt6cPiPeoMtU4tISqIJUx6bAcoRYkVeC2WpijWAeH5AKLcNajF4zz1uWvo8G
HVUDrtpQRWxLDmovC38G0cpsyWKRdlRAzStWPQ9Fm5hwrIMhB0F9aAZReVnAeAt1NvsE/TEolSpq
QJxBcFKXvsEls5lY+qHm1G1HwtxBOXA+MrkwRNKxVyrZJka4VBmU/qKW8ZlzVBU9v6yH2db6X4t+
oSFy7uaWzYzwT6qmTnmiUuBaIFw93zHir2BcG5irsqZTcPv8t5t2SxBDz65mGLOrUP1IPZpJhCve
U9ylcB7LWcxD5TPrbQSmRqEmXdBCkF0qp7FpAUYYXTGGorKGp4ZDVyeAmcnFzXThO3OBCbhJ0/pl
swVYpKDc+sbuI+PrJUaIV7cUILSHnGCstWNqWNCVgYCcKBkRPOzfTpsG48WYab8eYkGt32NmVCsl
7msuAAHzHZJr97A+CW1Vg9c1xAPEmQPzPDOz7d0+3KC4V/1YFcKqT5Drd7oU+vPTKbql1VihOqpZ
RNyGjR9mPmexcaUa8GM76oLDwhjMEtYCyPCFtEuTxte18xNtrAahJ0O2nyfqYMpfIUbw6qnzrp2H
VgqKdCFINWKQ8qnJNAowtF7Ye4Cn2tNmFVaBbl1hz97MFP4hYeWru1phgp+Hn2oFEBG/KnAGrLUl
rfrjGIRipa3lGTpjc3e0pZd0ihrSD1GrITp2H6hi36bT3wNfcItkKNSh2zLFQSysFqWe5BbLi3jC
gswcI0NcgtPfk+U1EIq9JK20VXrWbQ5llREhQDWPBOvN1+2svjsePsZrYlxXxsOXFpmGbNjHO23v
M0t43c93y7KhiHix2leKL2W1hf8a9HzIgPA+G48cFxa/3PGbiHdutoNijAyeNrSewlnlOhSOCHvT
Wsrfzv4unOB3PSMVr4aqKygxPvu4kltilHMBuktHGZGcnlDY6cG8BS475F2XxcdAFydNMaqmleKO
c016NAtHMatNz0MVr+iWQG5aELIMS+4xRh3tH2pjN2e43SR/TAHa00eof8Eip/sZ6hujx0Xb+Rpp
26D/algCYyDQLAtio240YSCBKKnAA2JRiyMcawiPDuRRvBbcrA0WGtIPVBlxDp6n2r229VLLyshA
+EMUhBBPPViYiATwVy+zOOugBe+hY/fn+HWzQF9UWmPHSON2sJq3NxXW99U6WN3mrbdRsHEGDeCT
UdCCGuw23rGoeBxyZTiCn/8a7qtPjEPEOn8JdcD1EzZ1+u2EsZNa1rIufAJXrSGdMqSPgYJOcKDe
y+XD3GNczt3lLGMYG8ykCL4ev/qhkkdxyjP4ofAblbcHatWo7zbBTJevPli5wWdL8Ri2HnKoLZ1k
QSFHnYPDYlvBpjy+uczKQU4I3FplQcmCBK2jfXpYqSL70XT6VUM6aMwPj6fKjLbQp6DhCtQIYWnd
M0VSVOpPw0/+NIRbbWo487d/SLjdixULmHMYgQw3XOWo57afBxfsbIhDopy8gsOXuyWyJXu6rkJC
j/FJiRuqDSroZnNBdUL+sHlesrbjYbXlPlw5LYMzrvHoPxlAz8ivqU3ms186qgJX+b42lu6AAK7w
gBMUNiE9ZdOR/MTxRhLNRLw3mIUp3PSQ38FVTXqqx8g/HU4ZYamuhtZp289IzQ1gVy4zEyPTfhPZ
FN5/kNztBjLBPkAXgItC94oqVIFakMhwcGfKxrqrBEFc8Pk9EXLxfyez6zKfu+JcMFXc1a4MFl3S
pDi03zIT8E72mYumVIzZPEqt1841yUNQHNTRaSbaRZyAQVC6IcCDbeYg9iuN20d0YGJc0GEb7MV5
NprJlgAWlJuN+NoA0zbnsC2Y4I/TOWy1rIaL5MIQgyhntQkJ9Wp5zj0k9+zDEtLJl0dRtLBgJpEF
JvA1QEYcoT8oCc4KanqVEBSSY0GZFIT8KCnMp6/PPPBanTQHAz39ZANfDvK/wXKTi0PyT7LWRiEt
3Ew9XiFy266jUMKBD3Yhdxyv/G4xd00CE9xde00wKqpf6KXM0JeaFOuXMtIy8vtqgYvVzDJGQaY3
Kvqe+0XKzb3fRKK9K36PMTgCa2QDDKlqabS+KGlym5sqFuBGBlB1oU4HXQkSIAkEeawqfBli0Nik
/NZop/1x6K7Er6Qan7ui+z+9/JXVGNIsUJsnrRSPuBg20IlXlV5BF//ayXF1rXwFsXfwbMEGMHaJ
etyp6BonTlBhjmEIgEqBmrSQzN72JlpBqIj3z/JB1BUIq3bphZD2NTireaZL1KfU/QI0hZJicpDQ
VqoAQL959AlmrO8We85ezZyve5Ae+Tt8kc1tWNDSEInXZXWkcK2OVmNXOwVFI2mUmgFNkvVPUI1B
cgAHZhxUugVU1YJHY+NJE7o9os//D+DufQiTJkPhsXkkgd1MvwFQRy2Kriog6A73yvcYFmQWP69s
eUgcRHGzgEw+zeZqCe6TVdirPg+tndtmvU96CHmviAdaPDqQ1PrcbqWHnQFJ1KHIeB5UinYuebDQ
+APS/rBc56FqRTM47yS/nXcgPgGvmMQC+dBPbuIt6gncqJMHMXw2AXmSTNRpc5tPreCNvwWi5rqH
PSgOt3SxyMN8zJrOccYbxlmXJY0FiEcRIzic6NkxebbGJC4QAN5X2FvBFURN2g3U7GqYxhNH7brV
ZgYreOLo+XGkOgNEYhxMBMZraN9KdlDVsD4Gps+WvjAWDs74gQHrMVYUqPvnQwrf7Sq+X/2VatvB
907FztrP4p+NTvtH6ien2/SDS1xQ+L6R9wIn9YDyVu1TcOS13MIei4ajPzICZSOdLUSoKMjyj5sN
vf82Jy5XC+hQJQ0CBjbEibkDbKBGUCGt3a9zjsliFl1d5e70A1djp1oAkom2VCCxT3rlmp2YnTlP
q+pC5zNpexWu6TuYnjcFeo6QJtNPwCYiGM/uW35yx//MRFhZ+MXg8UaGLSYjaKGmFTB3x77p7AGj
A1pmtqmsn8Ad9xX5i8fhnpombue4OrqKvSYaQ/kbq3HaBw0+bSSSOO9qIkyGIePZC4R2jMQGGxIF
0UFTI0kGTA2uJzdJbz++A5n5ggXOegxYEEfXicOZ2EpXtI183lXLVGlBlxOTIXFGwYQFdsUj8Dx9
IBH3jVjFbOM0QoQpqmZpdHn94HEAoMoxtmXfIneEfqTt56AZb8T9UaEvitu+n5qBzGUhe9y+d4Cs
WJWwAMCZ2K1L4Wjv50ps6poI5jv3OwQuxnjre1EZIszngF8ryUeN7sMDhBabVTRTGzlCdcHCdRvA
XfruiRNdNAwPQBeLjKXW+VtEtUBNCm/oC6rSuUWqD/g9rOJVo715Gc7kNL9skC8DDI2+pnSQtpEn
NhAIYEs67e19J6HllKhHEVGFtoLVIP6DgbBew+oWDIflo4weTd4UBHAr+yaFy++AFWwSUlKj01qB
ZdePRf5OiYF24/xBAqAfl+cGi6AwlU9OsbOZqW84qW18LOj1aHjw3L6LU9lhD8cKx8zUAd1HLr6K
nXyNTTgzI1rQp+5/RFiL7iBh7ryaKRICN7RN0zwu5FCUFKdZbpDBegrmNC4XftHJunl0nF6uHl05
CNzROthrHDimfWP2aeVBGlodGq1NSpj3sAMpk6DTNYokT+X/mv8uSegYN9p/rcGOsPZtjqFd53sq
pQQiiyPfFcKOvStkpHdHnRkit+7/eDrCzypBVwzM30hXFMIuKqPMSWO8yG7wZ0/ioDTcOYUMicuZ
79icGMawaAKTFSnqJvmSwZAvsSQzTco1qIl46adkd8yJZu8s8I8TZz9h3OcUX3NVj26x8WB+M4rr
gfATtpuN0vqdBW/QoPOCHmxiEwvHtOuN0w5b09Eorfnb618aObMxe18RgtlpF7ZBAxYybHawAaHV
H9k2Nu6UA08852aiZaNfyc4YqDeQqi1YKrTu5Oniz51fF/GEWMbeRKRI4UwPjFSsTGVt1pt2d0Mn
dZ0FQvaQ0f1DxDJMB5Nv4u2T8lC8EbPPjcjDlqthwS+lFevr2JIyfDBwkaXzQi296MyKJjckFGPH
9d8mimES1C4tifmpHI97Hem2C4Xs6DkhvTK4v1mDZ+WYzJ6SM0n43vfGAEM4FbwhBk7nAO9CB0Y4
a9m36wmmsD52vsSAt2VTzNdWZCaqH7pGaZkpb495TCLkV8JHgaBq8+yrJlWsCOQfyIKPRRcNBvU/
z6J82G4RH2Z12P14Mgp6kChHtV7slq2StkCRB6trGIk94kxg3ltL22qKT7NkvZNJ5z/DhQeuxNWi
QNTl5iYZIb9n6/8fv2i2wJYVFTnGUr9Xw0egcQ2GBXg/HbQxS9GijQ/SwYyNGkUabcN4bvFhROt+
KWUCZ73y6aXZ/k50WyOwuJOWPRUte+yzwKgk3Cs+FsLOG6d7KT1EbZg69QFzkYFNTF57+u9dO69g
XzjZrAG0Lu4sYjdMChgMsi1uHs4eW48nKeb2VWbQLp1GwIqc20Wq/17aBHdmrTTku4/zT54UgFTv
Iidb+G2pAahUj8ZvIvDx8CIWm2LumFkBsfI8V5bg5KwKaCETC/L78Bi27zBfYc5UVBjFEklGLGwV
/OA2blLAVns8YIMkhjcvk/wf9xv7UntO5pgF4Tz016fAc0bv2jVbDSFNZx2mbzlJeQEykat4u2mR
MUz4r3aiMFNn3bCS33/HTrvpeRr0pWYq2QOUFlToB+IUp0CRbj37IYfiIANTk0m5InKdWq9CRBab
gGHmDh1JQ3bJawO3lziErro13e8Uzl6VMj0RcdidI937nyf+zTT/mZt0/s8BvEtm3rE79QsKWXWW
QEJ28pzL2oTkeGuYAbUOlAP7rdxXRYAPxj4MAselOnJYJRtBkZFX+ufVWX9yK9D/aCBJ93l9ibhr
rD2kTZ4XtlFohmqQLe6PvuNz1wIyYJWGwdlbkh+Lfji9yUf1Az8vHmgrGLh/waZBZB3gw4mOmc8j
bCVSj2alp/w9DVS9bsPppc3h7+e7fBfGXs849IdE6v68qqIqqZkL/0KVznUiqUO00YuOeIxGNH3c
tbZY3cq8CuRAvlZmQzmr518pJ5+s2j5vfIog2QFLJk6Hws9BI//0AEUTmoXDszpQMZbqKp4zJzW5
YnfWic9/aE9yYqqMyNfyxthR/if2juNEU4O4zYEcTRrT1HVvBMV5CUGBz8Uz5drAUA+tH6vJMmJ1
X8yGf/24KuB5ZmOCPlpXAQPNqK19k2A3WLiALHMQ1gZFRx6u9XkeNkBE68tlRFSMMr4LV21rX/8c
VopXhYLq84xbB9du/1lRasjcReQO3ojifz4GliXiF17Nd1QjaXxbZHSEamDUPsG72fe6COScP+MJ
Hi/lpaay7n6/HtTiZHwXpVSiYWH+YvfIAypSOPEKxPxPeKmP6grLEi7D6CEmAPBCcWANCRTAx/Rr
EVUCS2R/JVy4YaJqheURRmtIBhnG8M96m5KxmQ1FBzpX61bWMDkfzESf+H3eAKJZeFZHgNB/SHXN
rs3dKO7Bc90qyoWGEM6A+hNx+bxTOgZxz6t/MpJzZz7hET2TWh/Vd1+3H2ktRKNF17xUapq8BxSJ
nDDxB5tLDM0YtmJnf3RE0HmNyeBaGfOtE33qgzig3UWkQXjdi1i/gzasPRYGOJLzyKH9tnMPCSUs
FQCxlmnOV6LaCVoqq0KNNpCBbi91/4FwrdBVlxdit6toBrlXO9nLo7vtSA8xrgT5edttDyM65WPm
GKQ0LUbu8ygGTqh3ecfSUco11h3wq4N1k9Zl+QFVbMo64HI0ws7+3LolFxkQXNa5UPesP29nryaG
6YYIstudgzwtghpT43TcvvvYz2tJC8zjE3Izmu4JHfl1q8sxKxZFr76vNSxi03xt6qxbf6kPpUqM
r9btf079L/xiWkULo9ErtIYucURXVht4HZQbj1kAv6gIqfLfDLvsnjaB1LAqW/1S0ip0Nba9x1eO
3vpln+YwxItCs/Z4aPu98NfE28GStOuSNX/FqdJIG8to1jM6ZyfQrhSf/fjvhVShI4gekpwG1uFb
+VnZqklMvc8eFcFJPiSKM4BRSIDrwlZTPHZLMy7oDmVv5nrpSBXgLXZQMIiGHkCDTMm9MZ4UYkoo
sj8h7AKy4opYtTj5To9l8ECQbMjRiuNxkYs+FZa4yTXgqmGq1tl+rYO2VFH6O2fl9UzZrviFEJTo
NnPqzpcK3YhMu6L2LgUgP01lg0BIMWvfgFFL4+XER0LAlwOXsSiNoLrz9/7zNeykAZS7PKoZ9YTf
ECUgpvvHpXlqAm4neSjCbQyrWxJBUeu2j+SRg0Kp5sktCuYARXunxnG9g0Heo12BWGA35nfpqUQ8
O2e7V1f7uCxxbyCDiQu5f03vYddCbuiA0dPcMQq1H22Foy8juFFiooN6aW6Atgh3Tun4v3HFPwX7
1XfjlqgCAd3DatX48ajhfenEUnl1T80J25ty/Opa/qp6dcvCcM1VcrycCnRDZGnt2tJYfuOtSamJ
RyYGch1ZChAEn+54eZBtmhrjQwMyankFhf9PbbwuZ2ddrmFTmztersMin/BylWrPB/AeCdXh/F1q
gi8d0GPi7rvba3T66nGdGTMAvwhRRjsbsGo1wyS95a1lNJgVUIrBPFr/NQqfEaTbTlyKF93R3yTr
b3+Lw1yvLlu4xUk+TnyJ4q+pGicroUE6Anr/JHOz20NnfQLANVw5XROnNmJJNm9p/x0J0O8u9IaS
t2VCs+JFoq3ISePIPBdo2cokQoX3lj7c4Bj2r1yusQHQzCEAsvDByCYJSbK6HdrVZyAMatxBEZpX
rY8DgG4TFQwBrw8+1p69PR4o9KbNVaZSuGAfdrvqLzzyAC1My08blT2UyOwQYKm4JL1Tg2wenm2M
gsu2XsWPzd/FZ64+q3s1qFx2w3FUx5VyHYuX8h6bP85P408mvuvHd2vJqrHRKOybfxvzot1wLCQ0
ZNDEA1bfl7Do/lkey9Jf0xZrx2a3Zefvq4DXQdZoQXqwoxUlgkX4LoBuJOTKczM7cPxBYnWAm6dp
7id1nxpAR/pRF2ICU1HVW5DF4K/2UEXKnH2YPd3sz9obya03AvloCYnkdSV0eEml+7JlhF9X5RiJ
1NoncwXG7EfEzDSuoca1TkWCCzCEfugOmrcBezi7NWcIADWkydiSCOOOBU7IPDP9dGslzzUTlm+1
B8Oow5tCxJ8BabyeBhS+UkwzDO4TC6Sfyl63iYOl8un1TUlTTBE2T10+816skXWKb65cFMnHjfXX
KhnGnw5w9OgIp3LxslLhjW0pnmUp8tUJfdTEGIBxB01ZwlleZmFTCba6WzTokBXrFARu8Qw7qt2b
JW//4lnb13th9txTVkX/H3SLodDV+CDaRUFucCpswARhSADjvDYqSk2jxftprbo9vXQ9RyWrebPR
w6gn5pbLEZIQtavPoZDUOUqh4eJEr+4lKmZ1yyymmgflE0o3RP5C0mMKoMMpBalFc2yzZTnZ7iyk
GyC6Iaey9pmRJ+CUKNocve4vGSIrUUTwjDJTsxqPaqLBYanN2Btqk9FNTV/EhMlR1zDPIKN+2IRc
SvyWsdGmrIL/lGSs+wJPVoolSdB3j7wy75khwW+n1pWNe65M0NXRYcwuhDKYcG7joHom27kFSAhc
ospDG9qMRwiS3iZ6JHzROD5+d0zbCDUSHLTY5ZTHQz3VIM8gj+vKDK+18x1B2gsD3KeYn00lWmQ1
x+LrjzVkPmjKyRihflH7lwsLbJbMYVzZ8pCIYjiePJDAZN6qwWj3roLCJUkYYUMu32U2xndAAgKn
OEmSA/EAQlp4wpSIfUZ31695O1vIhKCXt1x/fKo1+P6MKWsuCVMJ1mZ87kjR3xEXvVN5M9Gwd0tD
qby4iQ9RIIqoq6NbBvHPU281IbAX18diWI+qKUfsn27LErIVVfNr7yFuJ/JKnRSGMtTq1XQqPEZ6
8WOcLMwd/VW5uQYeY4k5ynLkCB1Z1Fhn0GQCNdcbQmbLyjuYKKxZP2/1kpqmi/vOHIi+T4OImMCl
P2iV1255l9v8/UbOHtDMvUbUtz6o09JgQ8sd+OmhbqKJ6rDteYuE+/nQ1B7qDBRL9Y51WLAoX9vn
KmHhb0rhpPZQJEfg3FIOV44x6EimGNUHtp9aFG3iV2/CT90FyKD5GtKZZ3dJqcuCRXtVB4DGeBey
zZPh6PluWf/F2P3fQ20qazxi0t6ZuoKI45lj1Jx0qh6/XrkR70sVVqRzve9VmhEfJr/YKrKRwc4E
KSmhY4wHC0d8Pusii9XJAFJhS121GFRA9VmIxJisvPT9zh7OScyHEoBk5usvx2ljZ2mRzPEhyT16
LKVt4jCFSu3TeQCdRc8q6lWZruQOJ1JEP23/OdHDymYJThBJfqz1wAKzM0MWdprjwimS0wONBd9d
dupbWY1TaW1J+fzCkwMMiqyipasJo7CTnvZi7CR/VDo+76Pudao1qpIpbWF2Mj1UGd3jD6RzqYIP
DoknhuYqXTnfiWmWi7AXVq6YeW4jsOUzCBJF8gQmTMiOTHNOuMW0W0yeG5EGwPvGeWTeJjMv0rcl
lSEi2hqte4OUs5f+A0NE0UBUmqlY+eIQwEyI5wXE8OANzLxbpk8YsPFAIFCRkBREnnciqOrNxMFr
/qSTsDpBad/uBm8lNklestjZcAYsrv+YVwZ9kxy+cHiwfPVzlMPwnN+pyv+DwmR+zvacZ5P+pEFp
w6fcbSFcd8n7ppEPfwDdwIPsxG1V8Pp1FQAitsjBCVH9UdpVBCXuN4SPQj7N6SgPpPHeHtfwhYwr
meNSZLWWrbNwMXm1cW5k1X6OyRexzXeIDV/d7lVbyZqcvsQXRn8K59ge0mQySRiEudQOMJnO4TWV
dlluwxu7rVcLi95ws3sX1CYwtxvOqBZQftjK92dVdI7BpYZ4IF4AZpx6kRdQnAOuYpBev4/C1w9S
HxT0NSUzj6Ihzm0PSpsq8qexM++d8SGS4DDZKZtAFwnkUbWR+dtAcbMA+tWLnTnpSdFg6iFJ0Peu
hX3zKWcxuCh+OOTBEGS6XvLC54oEjdGp0xHMirPdT+PjbgEdgsFI0XfOqah5Kd1Agfejm1y7qJri
XjnmICs4OAYKe17ADQWyZeSgjEkvPwThiyMC8ANXw21wNc8eDF2vpKpvDlIMGn3heA9xfUUInsdS
zn0h9ZmWuDVF8Fx/BuPtHAHG40gFeMtNet2icXePDWPJS6uSXruvv9N6gh8GTdosPNiZJrhbwSu8
B2i8SMtjZPNFvwkAqe01f+KxIFmOWHhPsTEP/lEzfDLFNyqrp1I0pzAG5OYkjsMX02pon3E4jhj8
O84pbMbNeTZdj4dj7A/IAIiRFC1TPNr8u6Ao1tuyLG7CDGhdXD2kvFGnn9pX9Zg+GgClSZjEkYSx
+BaeSv3/ebgKvA205lkF1fi7Uu0Xe/ugurI5sFD+PEy9Bu+e1IFBBXCtNlVI2aMQ5OezV3y7yWyC
JRf150DegsquSuRWaiePzegbuSaB6Tz2bzj+DD0j6Jmc94wIpefIHJp3+phQK9S0aaofvs7fipEn
SL+iO+OfJfF1xgLk+U+YErZoR2DMtqz/al7xB9PfSmYDBMIIvGq3bZpceqYYQ628d20F7livynGR
111gCpY8XaB9smYzaNyDiprhV9CSr9V5DMtTDtjQdI72+yPqcg1zMRmdWG5yl4r6jGWFsK7BIYML
iTHpzLts76WqbDfvf3e2y0rx0MxXwY3zJJwC6Aui0X4U9vbA3NfT4xoJ9t9p8eG4ZG0AIVh6qZbN
/km85uRcgPylbtgQB7328HomN0zgUE9piepGsOBhRlkjhBrbzX/tGvhJLqoh5MzNX+gH+VN41a3H
1tEIYYjp9arn8/A+Xofsy30KGc5AVFW5tymHAr2syNtqfDG7ODjfgBYKULHl1XPpgeAwG+9Ie9j9
C0StV8ur9BROphV+gRF/rB+l4B1WWW19FexWLlozgOOVj6akkRQUI+u4Ca1vmPxJKqIJgE2uLORm
wN/+BnQp7/lIsY6h/h0u24KAMx5VHaJXutV0VShBirwkiCqpjRLA7i8kf091wJSzQPNfJVkTNZIr
nBfoDUvM+7sqMVF7NoQKrUl+KJSi54FvHsJgBuzUPw1JEcB5eZhHfuzf5cjq/b8FIIddNSMGizoi
DaFS54yg9A5RtCSeXqCPz+Ix/oY4sWwzRfjHGgMJDl/3Hh9wbmaRfSAMMB8SfEap9CiIFllbN104
2GAb8cv7s4HAQawBeAEfxoaCy2hibpvaPMiJcnHG32VprgpQe9m07TI5dZU63gDIgEM0E1M6clIi
gFc8dljypW/R6D0TqmDbksXiJ1C8fZHQgvGqPXJNhgzfVf4mRUo0QrMm0zk9uUt5QP/dcK+04o26
EkHz7sWHftCQK5G1rvbMaqdbVRCAJjJV2X1JbPAY/ePyTJkcRPV9yaupK6pE5/NGCUQU8KQNu5Ld
slPzVO7iEeZKSPCk+ti3rKSEdlcE+sFqzRBP9Vkvr3Fc06cDQYh5LzIXhd+Kqdbh/Wm+AeXNMO9Y
QMKQRxWiL6N2EIr+J3uy1Y+f1Tnc4f9Qk++k2W9viP1HbG3/1d0R+ep9ZK+7Eb0SwZSoIUrnQayn
mWQ7O7CnNL9lNftaM6QtpQxzeW/vWRezPgdDuCsBLzBxeu+9cqn5+Nuq576V11oKxpO3+IB+IsWc
32UaGfJDQFCJjaybpIdKownp9Ak7o5wwCSdcLWRBkqbHeYEjBZtfzqmHke/N/iXLtWTPSGRkDAVy
Lc08GBt69wBZt/W8w+yeNZSTBCop9xjBpeWoQu6s4pqLE3ruIVCseUv07kv9kRO40e+Z/qQhsJCz
7z57tYQV9zzpBwJX8WduSR/5WDisCbIYX056Rdiqpzw1ug+002egU1lXk96ryMCowW3dnnJgLvDw
Aed6eblxoPhj8yoVW8Nc6GHkM6iJT94dckLrZzJ8yLLC4lLEYGdzSLSxT3OIAIdLisnhwchtnH3r
eKxXfDUbAXvfPyP7PclqgSEcgn1JKpz6CE50STh6MyreZFHTU9a0FqXmcT6kT5QMSLCyzfJ4se8G
ocE6t82aEjc0r2frsYxFO8GYsEvahCmUy/6TlZEEJKCnKscHL2fLMGhFVEQ9Kdk5uZmDF1vKDSMh
qwqvOTA2s8uNwamVYC7+MRQSR58rCdYIGyUTUANDLYg97tkM4Li0vp7S21lc1tjbGOUjLXg39sAw
14GIQRl+MJS7Ryu8jkiSXytZfyxPVWWfso3k+okDUs/0VtCa18/2sj8eWaNhfxNXrdhPmLs2Nx/+
5nuQMZbYPl3Ns64QniI7Rl81ySLeaIN/Udg2giBCLEoQ+EDSy03vEjUWte1f4+CQ286gcNmx1YEJ
VUmRNDleN6gQu9ZYKqgClyF5TZWPAYvlVVV+PsmoGOtk4GrYzkHJPHVQA/nEyCUboUmIEZ7qLpQx
IK8Zso50y8NVAHXnnJ799prfholpO7nXciBvjaOURxUURKQyDW6BsTU/uVOixsLNoSHlz9qxuttC
divIIbS7SD6RSZ7WETvLhUKZBzcqP0EPm4E7I+ppRkbw1IyzMd4vliyeH/tINWndKJiZP3DxOq33
dG6AJZcOjS1Ak5Riu0DIXx52hI8j53w+FHCoUeicSyX97DM2owHCCxhBvywDWQP+I9GdLnxDnPPt
kWvtk9MeLhDhVLU9v/r5YUes9IpgapJrPsBm1zq2iOrTGvPkwL/uEW69ibnDV5urrM5IgYAGWMjT
6a0QycXvoot6nla2lKJU8v7lGl0NEhfYbiACTfbuIa66yTHgi/9s0lChDxCwmPR0701hmts1E1EV
pa4/WkgJdOESEXKom0IHTfE5QIwN5H0Zmox7nV0cJJawxwUHbcpyn2UF9d7Dpb0r9kVtlPQHoyKF
KV72QmaOrqul2+o1sUdcbKnILALkfyR2HiTOgx/jKrBA/55oLQeIcBvhKzN9X7bJNneLm5ctlXpP
RxJ9R91n1wMoMzNgrDlu1swXV5lr6SV2rzuMAlZvadvMsnD55LtlhFBrYwKk/XtnypsFbzODRkca
vpn96b4aB0g7Y6TdUZrCfOs/N3rPCLXQHoSPEMoBZLntpl0k0WueoSJGsJQfD1Xl8WdpktTPjRAP
m9hXejhGLCidcpf7r1bKF5LaBXg3RgwO/QSSuNOLB1G9E0IgFouySdovinbUPjL9geBFOJQe3xfS
+6jIA7r6RKW4gNzrhAmPoQXgL3bE9a5jbeSyC9y/jbM9LN6bY//BUShJKY02MiPA7NrlEMmFsA6D
nnKXOivmsexHWezfcOuAmyhpQX21t+LrVEJPbmM8nzb/c3O3nYtmIy9ZLba59TN5QiBDKDy5R4vm
dK+tj4tBenEItUYNiKzHdmpBokfWk8D8SxaLE30/fdW5/pH4m3tqwRdBPQkhzUe0UkD8btFhzq5g
uBe70vSHxM0O75ChyesS7LKZDDgF2y6HHOakbFSJssl1W9pZx528DWSm8XpWltVNypIfqU5NdQkK
mFrbFlwgSCs4odmKgFawFV0bpi+URd7q9i9/AAVJrXsZlp7i+LmXyBQ24TUPqPw0fac6tdfLak2L
kehiWBKCWWrWEN114QddZHsZPPobky4jge4oNxFb6ujqNeEytUkYXXkIjl1Irfu8yVWOoB/9jdkG
VkISrypWIZsGxHx/C99Fc2IADWoUjkkxqtfN4G5/x3S6eCICUFuCm4qbDFk5DuK9oBcgdj8I9bJN
IwKXRawY8dwp6O43jFsG11Cfyeq3Ik71K/efu89olbffoViO62baxzKzDQ3T6bYA6rqcQP4f1CAt
aXwxVOduLOsf8YHALRrSsrEy062a4IHkWpgnotc6K3KtFnqHeGd4BgfQu8rnVrokr+UfMbyM3GRi
M3yoQasGX3fpUCt3HV4ym7lznMu+y1tkMi4+ScoAGcGwD7Hxtd2OOCxDEDb4fJN6tUgNeNktd2l2
aeJ2QU86pX6BVbUYwdZxfuU0i2R3Zkc8cHGK4qf1Ny+ulpajcDnNRkXR+qnj9bR31psTc9U0AXGq
7Cc6r2QXOKPB7kjmKc3EV/ykWV9oEH7jlj/hVqvx57MMfShgDNjg3gO/E2cS+68quiJBH4P6W49w
WWdnzx1haQ+Z1zum3DgW6/LY+Y5B1XDnicP3UFgZSEfrjpr53Y/98ro4hw9lYVqDX2kUzUIPfZVV
ss2roGp2grprmKrPC8XdNNf+a8Uxso234eO+G6Z7pKRyZ1uG4x6MvMu7fZmVo8s9IvmzY6pFXmBO
mJq+lc0HPz+5pEXOTorF80uEJx/UHUHVTU75sBRa2sQvXZ7ssiYuLLLhSIKJeMinryVrQqBzWG41
mJBLiVJYrwtZ9t8ZBleO6u7ccUIPR2U4Hq8Ki2abETYgGAIfC0Ks3VI/+OuVSWbDZa/1t38PskAy
UHyEcnq1rWHXZQ+JbODV89GCJwwaNsUoThRTJjHXEbkh8SaUcBst6awsygSChikSlUdrgsruOzrB
qI+aiVcFGc5LJ5dDFFUlXIpez5+17fF0XBe3yZ1YFHWUlx9drmLmrQDqCCuItjWa5GgPdtKFjHxb
zL2W9hRIn/F0+068vDzHqh6VCytlT573jr+R7W8J9F0jhOmz+IqWlnbSGQG0JaMtsJIvDxn1dQ19
Y06+510Ds+QiNEulvhgZCh5JWU3BrVW1XoXHCqLB/UXeEY4PKGuWmlOud7YyC2m/bfDAHEgjNZlg
Xm4P7lqCLs5eRivsRJxBiFEughPwISCImxWdxEqLm93qK+uOa0aA1pp2pxeLV4qTXGU3lRcdEXWo
j/aZriWqcrBwppPbItAX6xbg12phS3AuElW96t6ZNlIDGvqjeTUJW77yTpJEy5wL0tKI7Yokf44+
FDFi9kqbi+b4fFAveBl9oWhpZVbkrZvrylUqyOAz2LdzcHQYk26+vPoYsCrs7yI9aKKEcw34NUxc
sSbMfVBP/udCBJN5CMGBkeidSvTNY92gq78eIzZ/m4Knj+zuXclj77aAD5RRvByfkf7yYXxIBKkf
Bf9yXy+aUi5j4O8BeRv2EfiCgjo+pCtIt+e5SK2BS0gYre6YhPdSln++zpPK9++IxoeNLL8GobtU
+Qz8Pb1ZwOmISdZn2f5nySPDzjg1mKgUNcxb7BtA6efGAj28Wq7E03epZLeEqvoLHASUfTlZXNpi
BnWIs845fH31k9E2+4P1Vrdpu8s/W6OH/aHiWhk53zzqna6aAU16+Au4jL68+6u12w4wr/jh55y3
UAQPKuM1ARz6QNBiqw32w4DrTfqA0QcGyB9hx47bBY4AfOVmwVgOXvYjqdMvnO+5RIi9A246s/M6
TEwtIwUPMN5qFbW70OJaXPumBy2pyOli1krGbAHNYKZ9Tfac+TKqFSTnNOpvkrIBD1gTMTInZdB8
/iiTO/2oFeoMzISXAI1oSJzx1j82f7AoP3OJCmtlviU79YnPjm0YY3PimyxxBMUuuSRUbOS5cd2D
kuNMtg+S+rYiI/MUUWVBX+XIk3PGJG0bPTdbZEWuItnxwwL9VWq6mt9Woj5jiGGNBZCCYM97JtRw
23husLZSR33q67QtWJXYEGceGjObqc9YuOF+1Y2whifuDeXVOfXckf5UOfm15Q5+z9EqpdKGVu2P
Ov7P4wsCKcDj+B80dzw5XRRfLv7SKkJ3syR5BQv3Antj6xL0+D4+rNHCGo8SjZKEc7yN/eO5tDRa
XaiXMG1MwmZA4OCRqgsVdacNRa8fWuqoVYhVQG+VfY745fH/N22yHQn7xisAQy61i/OLKTQd+20k
kwogFfx9p03nCiAnfJShzu6cOlWUYJhklkEefNXR2P1m6ZLslRqQCuZKLtnFvA5Xp92FWmYsmDEF
ZqcsIGxmtSbslZFWHEJQlIVJZqrOnFMH1Q2PbbS21zkDjqi5SYf94GW6mf57wxwosBqjI4AswK69
SRxUFRcrdNWNN2lqo5qV7offHAMBhAgLP5YO0UtiqbWylhkaPW7e7tMUTo1xDDhHgBeSHg0uX0fC
fL48uTy+ejU/iwciYnc8jgGxlZuyGnWhLHfuWzFYQQxHT69LQHOao0G0oGjzS89iDIsujpvar9PA
QQkUXg/7KhCLJsbY6Q1S2pM/nZly5gGE0cbD/LB6iHNdRxD8womXen16aEkgs/LbLbq9R002ggKs
8t5Xf7KvpDH58MYgBaPupZYYcRr8WRYf+p6zR1Hv1MYnvjp9+xSFULAENIJ5QlsO2G8joXfLBW5Z
NwxAt6uOm7f3ZOLxTnUZYtArA5KUHnYI6foblcvaJjfSuHrhQd20tS+P2Wv9YP66xw/yefEAp8Lg
637/lt9buxJLMLoRHp+ojHEIzDByXj3/F9LQxpQFTUlqfCvbXOkLrUFXnV+ol7mtsiahK7AZ2//K
6N6A/wIY8Fd025kTa+EbM0oSVt0RCEPmrh0mztuU+BvdUaMOY3CJkO8aSVIyPgn3IEkVmf1ixKIa
NMnU+qwRJtLeUp4aBiYHR0/ociQpRxSI/7HwQMoa+WYwD+TdxwGA11w5MGHMPkO8fvCttdj13MkF
rJpebVvgrnKe6Mf5e0YNbL8mn+USplDbh2eSrA9I+ONh2gmTOcoA186G8/u5EXux2l74D3gKtQ8s
S7J8rA0bLOJH7buBp9dOVtAwcm8XdQJjLS3Dyc52hQuIImVgwF8kTqukxkyApvafEl1DWHFi5HlE
b8co54pJeGMKtOKiJUJDJmjTjaTEOYV3oPe6fNQLA7KF+Ovo/JrKUalgw/JelPtWkqmytqq7hPBp
xL9rPuuu/slJGdEAkaT9gkQ5g7NeKjQwVwtzc1ofzLIS7K99uE/e1E5id6jTbIAp2wBCddzjoQos
Qse5TwV9GuaIopWu0ONvNBna8XmvyCLXSln7tyClHbyVhXBlq0DPHg+z/+YiRT7xMaZztBqCALyo
5T+CHSo30HqhcsphnSF9SCFOUgzehTHO1EUXYhQaUxH1SFc9yhXUsZT7KEEOYtrNWkzzh2m/SIz1
NunaGs0039meMel9W2xVY77EnkICtvVSG6mjHVpdc5i1SOJB1+n2A4LmIGNxFBFuStRNI3Kjyldm
NQnVfRVZqz+e4ZT0UjrbRC3jSWsMj2ixxiC5T0MAx5aNloOhNamm9m1ZmkHHoiSgvjTzxjpzBmMj
RM41GC0tJyldY9P33ZLJ3izaF+diDQVGII2C6hjscvWzSSaZKkYqFArCE1r61OgH6doomsiYnexa
pxdwmKhR9q6Gfy6vZ0BxGbqomlllfGczTS+kXF58iue9VxjDfHgYR9TNnS1w29HiNwR1xMcBUp1t
loM3lcytpHl23/HiTduIz3eDvc3yj2ssn0tCzD2gDQg3U18dt9jTFpgT/brxSbgQbvCMt1CLbuRs
VKwkmmeuH9X77uGuIRZ2yJxX4aVHB55ctxNfrPBfcEqpeJG9RVrJLKnHGop7S4evC7vUb316N+r0
mz99a4G3C3+urd5SzNM0UPdy25nPzpwwrxp4wkAd/kX2UIs+B3hCFFDdD1mCJLxwqJZFPCLbNXr4
zC2g8SBxrDB7tJrdpxUexMlt5Kh6iYieMuLsrfI4OZTSXWZFA8In+7Re++3/6BxgqFsCIpyGxz8t
72r+39aXSqgHFCX+cALB1zg+hLFqWlDbOaEwEF41jQNxgEDXM20oAPQVOo7ZzSf+2m63QL/ey4aH
P/GfJQyhKKuvrymzP+oUSQKfwr/DaqUyl28IsRSBi5ktok3eXjtg9uxtWmW/mATQWL3XrzGvZJiy
OYQ/B8qAVKKZeeXbpLwm7fJ+hVO9+TA0VjWCUiGbH2tj9HT8ZO8Ovd1Ogy5iO9t+0ERPV0vZkmt5
LpBXb64X4CmzahYpWO3Z5V1JdW4b9mHcmPLxfYvbNJ/XZDe5uYfIVLrilFxTPGpHh+4xh35p02fa
kwDsexLU/nyq6/jREl496Rb0tAskh/2k2fX9ETz80RhTgSx6G0Q5x/lGdT7BBn6weFXTS+SeZi/L
jfUU05MmuOTET+6cpcUlxcmfQR4jYGExwc6rXZl7aMWRa2WRjLgLMdvaC53UGKPWH2Gw8hH1l4Lr
jRe2lykgFcz0xrd8OBSGlhPe7bqhhL3pt/hcFzgjnVN3BpNBcgWDPvtrAeEJjtWDKFGqiuH5bYqQ
lr5jphuWK4axCHfyuRJ1SRZS36PC2zmVQCNlusK7G84KOXwQgzLhHJcv6eW/mju4Hs5AFR5O+luI
OoRIZAYJG2hwGIPn51NGDGrigrjjOXZFcYgj8pWXsaY2WMQc+vKNWeJXEsi3HXWP3xUrO13Hgwo9
Nko9Fj/LbLuuEvvbX/pnwsYNVYZatG13KYeCeSUoTE1OhFrYBOHvpt0aYYieDJ5xK4nV4wDLDs62
tY8op1Ca5jpDyIe8togk52gAsyq8etWQg5jSPF3NXC4Ec+WgL5N2YJ9XMrzrPRX/TGcUYQIPT2zf
RuM60gIgfZfot4q4++ZqbvxrwIQg5/EYX8q30M+T7GvpNSMOATQWGKEMq7ZVAZ4O7QZqLJh8Tplp
kBjR289x26sgFlFQxjVo9ycyESX59/TTneYomovUiIV4RP0hvREqc/deNU/jnVRWl49k0RA6HqWU
QaouwzOwU0YbyBeTzOf4H1ly+T4o6XtsvsrSUN55JI/cTH6XIk3GXTm7oOw4jWihTms1GpfbT9Jz
WYwjBK/YaBB7WoswAZLms/RGZxbH3XH8FY7doqtmxBy7op2cuYGxdbsBld1BWMadR1nNunpWZpIl
AQxjzyl4le6I0NUU/o08tBWF4Lp1kcQqWXsCs8p7drzurOQoruo8FQzTFhHU0+K7KEKztjASvPUX
8bIZ32affwkC6iephHSDcgfcD9wpymbK9yTY7IvUbj6LYEHawKPiQrl00jOC2833U6J7+GeqRQBA
Uat0isxfN9SUPsFzkZJsmHBBZAczUfKwnos9yo6t6dzMGhtnetpnj+rx2lOomZjQhhx1i3ObwLcl
El7x+LACTL2GkM7ZLskdWY2nVUFKgXFZR2nUDzjvSsGL1RwKXTtcXFbOfc5bTmQ4FO/omebzdBHR
RbzMb8+MMB9JaRa7OfB4tn5wOPy/IxKEBB1DrNNhM1/thH2XbfGxWOPHsujQ4DwI2dhkRv4W3M2T
+gd43YLq+oYmHn+3RonojZcol21f796/KJJiiVF47VfUWjOcSX83r6zRULDfx+YPcx8yTV/UDAz4
Kkn7FS5pzMs/r6H+du/fX9Irdw4JtnPHjBUVQWzjJVx9V4d/sg4fsvNfuOy7LaVcoFI1GYAxs2Rz
tPhKJ8822Nd1PocNM5XMkRTlz+8whzEx/LJPpn3+pYd2On0KKeu2Yy6kSo9MJ7bMqEk50cf0uFKd
ggexT/MJ+d75E7URXzUvfaqk+j8WTGmGOCkZlgO+O5+SkSpNzMT4btEheZqM1zTxPq4qID5aQx2K
3cmeTqMdFQ/yPGivwJ7s2LY05KYSl/LoR7ZMQ4i4M3PmyoVFrsKB3tDSTplHXD1vCHx3DZNvkRJM
Wm5yKDkZSF3V1itAA/ticf7D8UbxXUSX0/EHYCvuZovDgLuXagZcuz0Lnc6nh6x6IT/j0MrQc7Fx
+CrzkqSREAAREgtam6G/45sLFFGaHTUvFROZN9dXZFZ9MyqvfzgndDzaJRmJSIOobCTRgPJij4A5
1RetZZtKnoBuu5LPDaQ0Wannh/ruq9Hf36eUei5AyB9gdmpXrKJLxqNbhu9N732+Z58ofpEerLJR
8qb4xiI+UG6N0G79Y9cDcm42frvF7ZyaaGi0UrOMNcgp/xwDUkWv0+2hK3OhNwW9LrkUQBaE36NH
1Kdj7PAtRx5gJztElpQ6FQZM4PewGhumigL+KsZqvJJ1XrNY9oS8xaZmkTRFuVCIG4WJOi/eeSrb
2qCTvqqqj0yRQdSXeEhE/B/GZKtkzZFhwC+VQiH6YXcYFskknGQar4OqPbpRJrKiIR0ABUWLei+k
4ufpkE6PGdZw4awoAgJHJ4Ag6J274v/g6meUqZ/Gik9Vdhtzss+eBoF9xE5zKSh7q8plNS7+cqoi
G5WSoKi9zEKEa+t1ts3Cwys20xwOGuU8nsuIrJAjFPTsLpQ2G1u3B31k9SDqb8r02DddOsZQCgDv
Sk0kOplmMMH+HDdMAzl6jp1yIUVeSQtPTJYX56uPuaEFxiZ68+a565A2goenzVuZHx9VVVIuB99N
MNiE9iR6UIhWzVpAy1rA0coo6A8TiziR/dpHcURxxlC+B7+BFEuUclKYz7NUObWVnuBmK3cEV0P7
Miyek21848C4fq/Cnj+AW603OLjSQNXjf1nSC6fH3wGN0LwvUYgu9yE/VZTR7IXlIvpTlW9n65Ox
sxiSihBkB5UrlXiTf0D67F6du/xd0oxUoTxwU5eHmFn+OXRE1RBkK3dKyYb2KcKvYKQGe2McSSPw
3erQcl5hU3Ot5+swtMFK8GER+5aj7aWsGq7SW0DWMCUPXwiqv6Bxs/OFRkldqZUtrE0wiUHn1/Et
3/6IO18S02nQIhw9bEP0eLAV8KKRj7Ia0/7ZId/MqrWin5AEPnxxlm1dF1HhepRPyh8e8GzrTrYF
/4TVQal+uPyfP+V7QzMuOEFKGd5fiCDNqBVI41/iGZQqfHekd2A/u+Sm1lN7ql6tPcn+kMU0RDCo
ZwyMpJAtV49mI0m72aDHDxGvFj/EBqA8YN8GWOF+TjG1S4SzEG3hp84EQhRbul8gOpinZdG4Nhvn
lRaDiKYjw3eTBovojdtoBIfeIXOi/Acc2hkrrlo8H9LlDY/Y+xXhzfRC0cDZOylHGtPMcIcuG7Bn
3wndeqaXs3FUIcTcRV8FNGOwVt34ctctwL5jiVpQVRuFo6ZEqFEAq5t8S5auKr8aHrm1O0tOKH8G
17txNJtI7LiAo8b5ALpEGhfkOUqs/zHa9YyD5xCLfYZ11r9dOeFvjSnulRm197fcysp1Kv1/L9l1
0UPeqjuWMeM3yeJvdAgkOcgkQfkIGjIvsAxBNm2Io/c1AVVGgdhfeMU1jUlsZWD97/T3veYHjguH
owCdpTvDBzkcSdAcPegj90PwaJQItFRIGhusf8pszAp/LndFtKFayE4MgRw8RF+XeCamwxQj+/OI
MvwEFpqW4wMr1VC3pbhuJf6UkCPgkniHLFc90OiUQEGoNDuTRMsLjkqM3wAhEF2S3S/3uAzyiQwL
/8UML5COaSIemK1uH7doxh9Z2dTLZXBGc0pHxWX6MBfkLgpqqqeko6djAGFrht56qznVTNs2jBGS
Sfh0PkHh4btpFK4/ov0XZwK9q/WJzTHJZoWGKw7/QTsoxkA+CuNS19AL6pJ0i3yDx5zxS/k/O2Ql
l61obdIuwA/F9Nd2JuhWQvqIZR9/uAJk8OvmxOTf1iEuLJOx+ExfKldjYz5fcjufE1E3TxuNzjDZ
0TOfqAU7oFkJSyXnPfVfwmn7+KNc28+fT2YfBs0xFMVsILHpBWMVA1w2eGcUhgUywevh0wjZH2Vf
AHiBWebYnNxw5vRPdVmjf+WoEQFNx2dBNb9p46c4vnkqHTp929UgRlUcgveYaZaRYvQ4TCiZf2C3
6RB0xxhKT2P2brm8tTSv4DYKqnlj4t2YZlyXyJADjt9YBYPzw+nry8P73HNJIvlHB3R0gk46W+Je
SFuVqYAkeeOZoN1TgrQzX2/iIm/Hcp+aNoPyKqz9N8e4O+g9VxQBzzgOKKY+Z9yMK0S7wrzghAAJ
YZR1MbRe250XnU7WeSOFUHecDkfUIpbaISJMUILd0IoRMQPMJhPQmdKNjxNVCeqsZnye/fYblpXR
FXHg6ee/kFGCuJS76dXS6kjqdlRfjZWx1FLLmfEALAyL6hqqMgtW/eqkAo69Qh+JpMQnFqqMuFNt
WqP0r36zFU8NByYmngx1jpBTY/Qkciv4ilKDQ9tBMrrv5PKsDjf+uYI3DFHUYStJ7sKYj0dbQVmw
RNEcm/HRQxaGP/Ha4PRgGZkFU+6yBxdBhAtc/r+bW7WvclQwI4JhefzNYjntbfpYZayYinP/LUZ6
MSf/wJJezRAWojXqMvRkCSciRb/Pu/ia2VzPH7ac3zxLU4rfs+rOxAnxbh9o1baL97kega7x0xb6
1dIyHm+GLyvqImpX/eBoywZ/azleOj5ENfAgtdY2eq0qGeY1MS+dhkbpmsGI14A9MlZYVb1Eg4kS
Yw+ILJDPv+7AjgGlXlgOj79wk4SoOPi5JnW8QuEho6kPyLsiSvoUtotqaB/Aekv0mpXBM7m0DNA/
g2/CtX2xwEAz31HxbR643ealQUKhSya22buPF0AWnbxdv/LSj/Qi3zsfrCcgtT6fyeikBQFGXlXE
Dlpv85zkYKQYF1bvGsm25REZJcH58El9zfLn0G/6yopEUGqYSAlgTZp8mpubS755qxjpT7L1vPz+
o5yQIL92zlGmGSqYMgxq6mxx22Xc1p8QZjJLoNeGNPv80iNYKGaqR8XF41kmNCc3h4gcgQ8MGLif
JECa3UScXhAOXiKfFiWB7T7dzr2Yn06VaxypH9M+KEbJqEl2H0QtHJpgZnJ9HB22CUcLMD/nTi1s
rWuLhHR4kYscyTJU4RHkmpNeetjOzgNRL8xGLFTFynmYa4f6GVFBQ+I69ctJR96oIrF1vh+852nM
ARaTeIE1ifAVzcA3LyvGh1nSb23Try6PS9fHhyDddz2Fuidl/HaFzmqbCxJI8x6VzkeGIpMZCnT4
tyfuZXUVK04W1tl8GnduXuMm4uNvi0MsCKHV/9+xjOGRcS/u2iOuu5sgGv9hmkKXl6UuIP6E/Hw1
y2TQ06uPDlzCTd9Ly5sWDGZiKQUy5cwdK0ZBUymiG+ST1mr2JwKgkNP8d6mVOi1jkzw8XzFe3Tsw
d0OapTHWhJxzBryT7r1TbDCEj/xczdEiKCTPaBmL/hxWGC3ah9UvaLfB4Tk5BA9pec3hrqend7rf
ItzC4nm5obxgBPdmVPMQOGsydrLKRM6McEcbjLeSmNNYFmJ6bfeZ/y/rjzbFKecQdWLibf0+mpC5
UGTaRzMx8mttvtf7OozQir8u1jArF7MEL37zZTxqzUVvaBHdJknkcmxmGqef8buTTO/2Vth8GiSV
V0DM3Z3wyY6EKe9p9hDAAYL9/3f8pjA1xcQIm7/Rdh/8n7e5xnuBhELqJLjP8oMuYUC8q1sUz6W+
bt2MxHuUapsOryuaVsfdd4Bv16MHnSOt3JIJwm1PkVtkaqxvyP8ay6icRdTlbBt1fUNW7Vpb3XPk
rysqHKQCmt1W4oFoLPe0/R/jH+/nYwlrJlOHz9iqJNQ004KTE4GIPyyJcurn1i9jY0+1qwy8yaed
ybqkxP2JkwLBjezCqf8IEZPGb4oqbtKBuWH4fvZDHKatcQuBydEMHJ5tXNPDLBh5lDHEQRimZMGv
rmBpYGyACy6IZ3CfStOINoNYhFYCrVCPtPGtyRD8uwUr/KowzzkdvyjE3HjUzhDG0Qq5Y+BM1lWD
FuLUqAm2DRgXsvb3X/F6CMkB5q9ipts3FIWgJro1FSxBs1vTa1AqKC2C2QfkiZOiE4EGEyL3T60J
VoVC0zUyfA0v1kHAyEOKbJMD+OzzIlzTGHu1n/mKYYvnwlAInIrzDwkTQyIaIPOOt0dHzBo7jeZQ
+AHnDAayfFtjNeSAyRQoeueBTli13Kkf6IANT7m1daPTsr03YDYwAJpxalcVWMCdVb/JdU/FA8lf
NrZeRPm1uzcM06Hh8URTn971Wc0n/J9UF/fg6Jk6veoFrz99PH3Dha4fRrySwED1TRBA9DKLAnq2
W7bDIQGOEPLn1Q83exniyzuVQzml1ML2hGPW1d1RGhy9h/YL8drWG3o+IVJlExx9Y7pHSn7/UAnr
IdVWqsuo11BJabP1i/sG/0hB22A4PpgCiA3BWoJ+cB5aVY11vqO84MO9cEmX4iUt9NKLFmpAeDaz
JIaZwAYQZcH5nmL3JxXISA04xWlwFvJcAFoaXPMXdULUjZNp6lOHiWkEU2HM0QlkrAX48z/JeVf7
GjouzFtvm8J0Wa1I711RabmOYKIDZtidr53VruNQOOuxV+3TXq2BF7sCnWnQQSsecBQ9VSxsLKwc
/yd83Qjy/7dxG7jZJZXP7fcgWM7Alf0uEUnKqgatQMKjs5UNj+Fgx173jbd4xiixofcaI/Akq09S
vioiXJQabwnVo1IuWq1XdlzP4nEOjwOrawJ14y+mWRAqxA8CiK9Ul6/3GLiGLDReGl7jD1SdDuRi
KSnLl0G2k0Ii5eUrimVj1nF0F8MMwaFIHSVIvyl+NC050Eizslf9Zs/TVRLRuK1SzJ6ri0OKA5wk
uR4PyDM/JvahMn5Fhn1BrUAQVUK6uLtiQtkpJ/aQ87qjiIsnSHvbCPMPHwzKDjnulSN21d7OLVAJ
3/dqaT6W78JbIPHMkPwGq+fP2QR+RHUG3zeZQ88B4AA3dsl+g47/7MqOtNduLS4aNGZRJ2Ydr4tV
Avyel9ZA9selR0rvrFgf3X90mmDQ34Tn8ZixkyPeoocQHnTfebCcM1jspOybQWV9PXbQU1Q6nGE8
oHh5B9wAXw3rrdE80a0uFDdN+9lZPCJKix5gv2z1H2OiPY2f+An0+7ZVnJUgr1NNT4IFGAIgRVzH
o8jyJMz+LgdqMhj3Js6t6r5ABFfH/tXdeG+Ytf3q5QQuAHTwHYl54KMdE5o1mx9rYTevVWj4r+4n
PVVuFLcj2c1q3xSQZN2GEtBaQE/LKeHnTh35jR7ZPG4rnWwJNY7Li9tOgxKUpOl0Bnv3MArFAE9V
RYd8CZknCkP9TPYJqlBOr5UwKQ+P/cGgx3VdgAp++00glf8B7yY3VgPEPufGAX/5iHhvqtaBmIL1
aGC7jMte9XZyMfew68iiMNbPrnK7oOoABwlw4HD6KVqEHwwmQuf67bgM9eV91Low7lWrNULSm78U
fZrW7IzuEuLIPRtofTkM85fFuNI9KV23E0BP9aSc8svbQy5uM2KmkSTA7RIbVzf8aNZX7rmj2NWl
lIXUpkLADodckk+htBcg0uh/LcPDZarEJr4VcXzrpgwuvP8nvbW+7Z2Ok+xSyUJ3Uo1rM2egdrXg
6sF77ojh8SmFuvhfY/GCnoHNU0cX6owcfC61XDGU/6yDN5GTU3lS8uO/IzxZLnk5rTld1LTbVBwU
l39qs2MQlewCtB7Q5vdAtM76E9iU4JSx1TaMmUk10OhnhWnFDxHcOEfNcaj2Re8Ff9iRjvLsj/oi
UVOVsRYzT3K4u1eNGLi8p7GbTqjYpzLB4oXPPvdNlYU/qjhaQpObjG/aBIJWdaBYk4A2xPIIxfmI
h92TrLJSUSir4j87O2nIB367VGaTjYvPuopJiH24JWvUw2814N2AdBThEiSNACNQZWxzqCq1l8Co
Sa6g9BpV2Zlh5kJt/QszkXxhWqhjol2P+ei/yQ+XyNDjfQA5XEf8jVyEom3w7y9aSvej4uGlTro1
FGscWft0Pm6fUuLpEIihjUjF+8WnO0BrJnd8QtJOSY0zAfdic2v/h7qDuWeNvZGql6cUp7aWY19f
Qv9gcQ/OjPD50bqFxV2G9iBGsIUVcU6wsprExBo0wHm6/mmFqS0WGHAqNPw0HcsKTGAwARnb4kBl
rin11ez/Ll69CoTIzpwO6ajuVn5HNy0cvEdpcdtFBsKqUYeSnMs57TnHe7KbpB/W1YxnUMErKn86
mLfYawNdmS1YbB/YFJNS3SmOWa/hAEfxfdcXXuT5NcOJgi78ImQwZJXLXV73MXveLrZULxazmbqy
92LpIbiwOhCOJyt8k04j95N0UIB/wUjsGX5IMEOI8qJ/XGcY4WGo3N3U1HbKVLQNSGsgpQO42hTJ
dkqlRQt+CbNe+jdP9X2I6ZrVeP/9567mWqZBLOEB4Q1uS7vDLP89d9Mup0m4V8cbA4wY7gVXuya9
LgY8GaVTj0ixNabb04rg+5DPGc37j3B36lZoGG/7x5TQ1Kdc//tyBv2sk28r+61Vi1ID+ZmkNA8S
cUN66uplxL2VDXJPjHN6qZ+SJcfqYZShIERt+mE7XClDFFEM3DuUeWthDG8LuAyIRBhxqBN2m9do
30OPyaPfT4gewQ6MxY8kxVYru4vWafbfzAWx8ZFMwj7KjGII8MTKgOBYi1hPGKKgTVLOXwq1WJu0
EKmZbllIsDhGVGlC9YAUsv+0yuuGuPg2bAddQ4+WThaC2tmYEAPnzUF3J35g6tS+mqIVsoY2S/j3
Q76n9bORLHHSoZKK8W2yJ+8aJSJ2lL7zNEprTnE4UicDXYB6FJdDD1R46ho35WpKvDGi9RYq+vVZ
B0N8+c3r3+UUWxlMSnywpC2zvfWpdmlxBj9+VWkohq1eYhZqCQr2ozs5KJICIgRw7afNeeMsC5WB
fkkUi1fi68adkR1jgk2FwM6yTYnuMKIhApE034TQw1QjFHsOjxxkAXM5rXQGavXtPqOXuHJ794b2
/q1jMOatbfOfin6uPFp+cBgFaKfv4wB2lALyun9k/BvVDGOaisvstG2rDWweBf+hwlK81oGA+w4J
f5V/S4s2NBkDvcZrlIUWuuTWI5tbKyiAFIEjSBUlpo8TiC8D3ay7unll/oGhM72P4xNePO6j1HIf
CjIiiFsHRV13gOjZczAuDOgy2fYwhErxI/w2pAcZIwjx4HzdyCPhe08BEyMmMhuX/vFZXd9q8Uk5
VbA21Kf8poqinlfEr+1hzPkJW+gd07U3HhBHZn2X3nTqMvsdZ9BaT/gpZucsBc5ghLupOyXk7B+Q
odRLxwaVNus8KYN0B0rYkk5pWzdUBEN0NztFc6wcaztxowGLAjlnFdDemVySfMuv3VkGNdSyK8br
6aV+PX+7uQPYMRw4iU3bj8fgf3ek1yWT0DQnhp/DD7egpbNt7SCzsTwkJysUAbzRYhO9n1RDZcAI
sZT0FfVYnDb5UGUYRBLMoJFFX06UoPKdGgXEgTIn4HrK7kGO8/IXmGCzo7Pf0R6z9vqxP8MoRdZP
SUuFQNUPmp4ysO0pl5KUyzJt0SUvgSZ2tijuSMuJU3R/Qa39q57Qb0qypGR1M7sEoDuF01hU+zLQ
dqws5U6M5Mvg9tXIfPl4KH8+yxkRJXhVWx15t0A2p7QvZPnjNQfDBEId2/rjM2emDBIgKyFRH2pJ
Zw6FK0I/yHilrSvQK1SLZOnOwLUdNSO4hHJAyQQJXLZ27+NRf+f382xwLVCtUI2RHbQNqgaSU8tJ
+YH8aXobBtAzrM1seB+siIogKXDJDA7uztLRAV5iSHdnbpjxcDkgYGBxyrDuQkGs5yR+qlS2B4aQ
qtT9qqz8xvdR8Ud8pLpVEFlqp7p3vxDLKqaUjvfcPxeYUftQi/RORubiPwk38ONcjv1y/s6XjADs
01hcJQfzSyTEoPEmLm2wIavb5Tgibb4atsl5wZJJiNUnJtF60zI24byAPVjF+JINRysVktDCoMnb
pDbqGfNMAKYdIJTEDpRfDc5RDfxnCEG2yapk3RD9RoHuGOGz35Uyzp4usiNDmgK7YFX6KDtCI5+Z
fhnd+/2k8qhsgjzt3z+5sQAeeNugmywXrRqP8SJTfL5oV9/o++Wj7riNXznBdGYuPUeycHaGTI2t
pdI0jn3JTw7eGLW+Psq7H6/OUnwoMb7EV6Ix+h7yVKcgFeNkcP4aKqkSjWq4acdpu+fPw+hbcWkT
CUoAy2xpjv5LMUGcbtdHs05Vw0ZcZ70S7VXwAiS12U4WTi6hLMEUvF/XrdTXn1LgU5pdk7RnDSTP
yODV0w7oBoUBaUXWL/ynCC0Dj84m28ASj7oTpn0Cb+7HbJ3MpNCR/d38SF/1HobWhP4SefvYQDY2
P9H/zvTl89Oh/1NNZsrAFsmB8gtCTEX9UHGFp+voxWOvfI2Pdk0kl5CEJbnHbjwyoymNt+mLHPnk
BrdEmYxjaqK321tDm2duCqjlTdbtdl2YfH4DVUuQQ74kqeLDg0RpJ6B7myVfDsk1Tesv/4zaaF4J
2UXKTplX+7XJshOqCPujSibun9BixZj2+d2uKXzpPrWQZ5D7MgsqikA5k8k8v1J0T64DC/0aRSpg
K79g8vimkKjU3NrxB+5AbaqeE6gAHbVdy70nCuN6hyZgv1YGuQURzjQxiKfVe5eL5FsxERnlrDlG
GfIqbsDCpjcTyVkdje20uaDWadom2cLdk5fL0LVRB3V96Sv6jmHgQS11gZSOLx3gAMvVaxVSu7Cf
g9c5rJQfDMgwAPXocKmeyauu8TeM4y5IOhkDum0n3OhG3RA4F0K3/v2gKhlwE910r+Do/NasYKiI
qiXxV7vTxsRZY9PQ7pTCtEhNPM5tKrPK5KqGpCAujsrNBiTOTyCPnZQ2uvXLI/ZskJorCyDs169p
AWaJ9qLEJgyPvpmTbSdVuUW2/UpHAF9UKaB+mH2JzXV19hL/bB9e9NhRQLTw9cxXSsipVStq/u44
nxmF8TlKLyjPQIsykdHabV+z7EaTxFA5/caOkgHcZrKpyaAUsVBsnT9A0t40sJhy8/nRk4D9dg6w
1IFmURVPmuDCNr2pywospQxDOUnlkV5yCm/klQ6FxhpVokeeias16STtkROe8Sal8D0d/mpbBPK7
pJXnHkdMd5hOYc824MaNyzkzPI08sqW1vHExn0PhjwXE0ufmH+gSh6M0d8i0fP/CGhnv/OISf6zz
HRoEj891uhGn5QOCB0D8NRQeUhEI93J3MSQ/tpXKhrOr/icu0q4kwiU3Ekd57baUH1eia7P+PNn/
xUxvYhCgRH7DMAzREB8vOSSd8ODeT8gNm2y4hEi6eIS9m5YF1C4EkPzocEelddMwzbyw7SjPh4pP
TM3CLv27VXtnSv1z/grx1Feirnh+HEDmUrkJOizutmkxhkmwgeA284VVlJeXHqTOAd7jfTNrXz03
LkY05GGw7CW4W7jMrSujGsZIr1+j99aeP0qaQ5RTwMNjUUccDUAnzi4xsKPkQ7vo9u8NXkaUYBvj
G1xkfrcRaEQBlBRnY68XkDarBJTr2+DC194DiZDrGCFB1TMh9A0rowjgyg8+G2OKdT4/9taO0s2a
RcSs8a8eFqUu9Ed4cx+WSvLqpge726jdPw7mg/mp7f6ewOgEboLKSqiWO0qwLNVz2Af7KArRHdNC
nzBDk/fgOL9UocAslguiwV10sGqJ8lfuMWcenXNy4Z4LmCfZbVdh8TfSMpJ1znyCPRP2CV09hZhF
dZMNMbBGkh2/O/P4HPSTxAr1wgnaqzYjhsI0kHR1Ke1I6zscwqzAi4r8AxhzTXtb9MWs8bZYZrJa
QDqtUf0U1VFhLUQpxGO4r4Ag4D/AKA48aO6oLgojdqDxhRqmNQFMhzw7oPEEVx9O4dNdMqvOljsk
r+jCBW9L0BSdN4MP1ljKUooFdeFGWW+M6v79B5L3lJSMZULmd4Pq0fUIfvgLZrMleei2g17taHX1
P+rmBDJhYVu24Ks1lYakp0KshuTQ42DrR1QDz9N1S4spQBA4tlWwc1fE/u9Qt2YzJm26DTvqCspL
Q5Z7a8QVBfXMKgfhCjSRzyzDl99xOgrC25cyBdzOXxABxIh8apqwH2C4iMcCF+kSDHuU3yj+A61F
3apld43Bwvn622SewbA2Ls8YzI2xXHlWgKg1ajE/QzbkVPZ9GaMCx11Zgq7rnwqq26WaBxo+fB31
c1aKxoZCgDtKx4GlODmOuvHxNdJW0mZWgzwmUTHZxHF4G59WxioZJ5nTGkvjx3SqBl5PqT5ZqGFz
/vAYKatXoGbdznmBmUPI2o3YHnIAMbFGfC+PNvinHwcycitvsyhccnvNS7ymKUoCoEuDQdyuDOls
/49bkmd17jDE5WZ3OlhlR3fXTtAKA4nlT7kvKrk2S4h3Xykh+B4YJS0+N2ZJkQYgMUMasuuTFH+4
HHHwfnIp2gzbZWtcISUoUlaRfP7woEF12jLMkTzVstnLZgyA7tBDrx0m8LkqsW4nyFXHXev7EdiS
KVIXiZJny9KJJ77krWiBhQlRzPsK4HmOh5ooIWrAm4WGXVQ56r0FDhr3m9OcqfwD5oIuQQRNvpaN
1nDjRMcAxXIUHmWYVba0JhrIJtBAbrIwETRf+DE5vJ1xOPw9OwcWWm1Ezqoc374UbToU5ifWej41
8T7WlIw6Za4B79cjCCiR7gWdqnSo7UxbsPSeb9ciDUL38SzxGkXzD/I23OQ6zidsw8gDnrAsipvA
FHVE6qu/mb/RcRBJ61/GW2YMFEdroUfNntlBuGcvzMo8sfLkSfTvijJa/Xwz9aMvGF5ifE9mBVf8
h3+PVXNqrnetNrHjQOLB7uzoC90Ma281uJSD9pzE4yA+YoiS/g0y2dAMrz6vDngJAq8kTXvwmue5
/sSuRkVsQExu3SkS0mAKvzjzuO7Y946H7wZsrGQ2PFV9QOejfUlugDqzM82Oti6Ts3r0YEeG7STg
qRwtPVLQ8SRxYXYDXtnQk7BUC9auPUZm8Kcx02ObE6EtlbKIettxQWhxbSMPaxk3PXA6DeTKykLv
pGIUbYgcic6qFwfP7k9gxGRnOI9XGg3r4CF+IxVXNKZaoU+BBBZAtohI8miK2BZ2/l6SYdoWAizx
VHH1l4AKTA0PKnq4Io76QkOLYxf59FsG3Q16A/DEYucQIx/DSCsAYBTATeFiYRYxYIHLvdaED/hS
2CWz4tvT1TgLO5H9S0BHPP2zOrGGGV36TkNyHDB0kbNDok3wGV664xhdw4iT4CM62icFf0K0ul+3
1fUQdSL3RK/NM8SIVWg7HZw18JJkpl881VSbEe0PQqgiSrW2hBY4u44Mbe7btf+2NtcB5DczEAnj
QIyC9N4wKaEjd+q60kDmqvdweFBLyVvkow3XRxXlETOJWMhBvLGaSGlIJf38m6whOicCMX3+cmQw
/oX0Hc91OYvPk3SPUw7wxgN9W06HF/Ysq1/sQtk6ioZBgI7EgVLF7ir5xMq4aQG4E3odWgvhsFwj
cIxWU1Nrn3VWDcv7FHbbu/7M1BJq73O/tTSgGqNg3/vtzS43Olr3c6H0RqlRDYZDCCsdKyWxtkkb
SEcTfuM9p7Egtv1wUS5qkfUoWGv/7RlhHbJ9Zi73BF7eVWIQGK8/qmPwGjAxweqVj2x/Ln9RDsVz
Gkbao8EutAU4pN8kndzx6oS9sKvglodygBBbRkJYH3XbpbvOjKblQ6arLq5X0NvkVvP/bQQpLUz9
YG2uQLtOhrexSz6UWiPPbUdM8BzT+lmRZ96zOnw5/CSNJGHtPTuyJk2DEt9mt7EpRTdnRniuqoET
9jrBFpt1OgHyiPjXLfux5Z7vthLwUXoNvXq58BIzY4FFbROKVk0IopoPVn/njvn080cE6lU4wFxA
z4sdfh/LMLyJIGZLSb8pbFZMcGuMkaT2SjEV9wDX3X0RNGUW2YnMEZnUvP77kgcwpmRB5h2QX6ny
Ne231vCQqtl6gJQJUyWu7MBag81DdhkKnMIzHRVDXia3IX3XbZALDnWkQwlhxyh4veSgr0Jtf13A
5KpXxyE5TdEvHXXqtnfAZ6NI56XRA76Rkt+YSqpWRzdEXU2IL3T+EwnObPMWYotGBZk3LQ4a6/oz
p/AGOhsQf+b61Ij9pDfMWnJ9e+MYHkIdShoU0Xc67lNRl5A8EdESFOKYHory3v5Xy2LeIscSLmZh
++5d5GshjJRAMmh8Os5cxg9oKHgiTc8fHHB5PI4bYJyt8j0OBxoGOFuFa2cdGzattmvtZh+P4fAV
Ba63vMfD/qABGlBeBQeLIXVwFFQEK5v8FkW51s/fmUKNlt3+F4K3gmzjmOf42qtai7uLlaA9mNRV
7qMl1qNYz7+W6gGXsrKsPo97QsAjdGokHZoJzgsPAeju2WUS+j3kR5rspT3xFpoNY1hUJ+Wq43LI
aEO+EuNrWyYgGaWXa633rfApEflfPU0Bx1CIZARvfZojJFbWa9QSGmPEH+gKYPdgfhQ/fXlqok7C
RnJGKkjy4AGPJqR8dYPO/vFloJ58YPI/m2PKCLOw133m5GPgzEAsdvLm75x4qMRQgomTfLF7HvH+
QuYH9GaL2q1EfdPoc3QLn5+xPqyZal6kMfLV0E0edb+455A0MPTER+xQQ1Iwsy8wjWi+z0ex+y+O
B0SHBcBH02bYNTdQWqj5vK+D20osyfTadPF1DZycbP1Tjzcc1APgab0Qyy3gNaoQ8C9MqMB2AGYA
HX7v6X7FFkbX/b8sOg+mOdganC/TfYryryfKF5eWTdZc1R990Q4bzONowD85n5687yv//Vyfrotk
/mfQTXFpcpXKDTeSZGfUahl2aHOoQg1oMP8UjfdO3b0iOTQU4JGy6jx4orU1SK0129yvrhfXkFgI
u8rGgYHBBQN0x4Fxjgta9G8Qij0RUhrFwRYd4LrGOESMTLVyo1a8FXzejp5iDGO1Dz0SiPQRIEje
C1F8qCuPlN139AN8GcmmYG/8Bv0eNeRfad4UegcFGs63vkVh05IvaTUbiEB/E/rHOt+ABz2N21q2
ImddEW/xGa6iX/ZN8HUOLxno7+PvGbUk/zrtphl6vt6chfmcQlRnDREbxybNhXXLSqkKjL/DXeOS
pWFWypsmh7+8GErqphofCAIll2Effygquc7LtTKpTyCUkciFpzALadaGOREY6zgEDTgwdtyxk43y
kn4kOKlK1ZoGcNuw4XpQua22SnxcDfHTVYjbLKFQM74kvhfjo+SwnzaqGlh3hmx/YW0IvIwPxkGP
0Z2uGIhW9+pga9iybNxM9lscwcQsCtX6hiukY2yzxvRVyFghno2DXg6aTlfO1WUHdhtiqf4Eqrrz
eRCDu2JSWnnyXpTAMD/MVV5GW7/0cCe64QeW65pg5EVJth5QeULrumGZx5cDwUHgIznwze+oQmjB
F0E77cKNGGUwrRZ71/UBsKnb1NnzOzPXvz9d8hI4M9NLVmrvHAa8o5xVM/DsTeQRkgbhi1ovW0gG
Tw0ykpJj2yrnXwtKe5gcPO9lqKNaZOKYxSuCrfL5UAouHZHIBKwFQyr5WjMtTtCDFTwqx2QY9XLa
Sq6eUrQ9FnXQQxTHqGv7HKAv2R0IVKWpVT1F6m45sPRBjIShEp3XebhMuGM53HvDqgzANC5aOjEY
vOViJg/5Cf8WFQTJSTFSxt5gPIuj8NQw/MDVT7wcW2qWQq6PGQthNZXrvxD04Pz/W0ANoK0HqS6D
4mxMEUCvcHqzNN2p7Vt5SqlpemdQzEzWG0SpI+rPplTUeBKQ/Fp6iCXx9apcgGn0idJNjsAci1OY
p8E8cuQDaItjQu4yiEZ/Gecv+cdNTmVAnqVo44qAJ9QOznmC8woIR3U/LoklHqCcJ/mJinWxHw7c
X+LEjBWQugzSCtHJqgHufeDaq1lVtGKy72jBi3SdU/5Zc8pwiY9DzRxl6zXdAFaZILAgWhkRWUvg
b9RTGXX6hCmodWHJTNpP0uZ/UIHActOV2tjuz6/M56mvUVxDsHhuAs8Yo5EZ4iT/DXQKtAafxdJ3
h1aS1jpIzoMA/FWG9AEW1s69HOidXe7IPKx7IrQvIyoZfbVFBMLIR2lIcA2dN9aqr1C2gPusms9r
E768Pv987bWCmNpU3rTHeJDNF0OnrHtnjWq5jiRmT8sVz2SbYitTNKga9NB/0+MK5zmmhjk2aX4J
TdGXPQCAxYQ0mbOoFIa3zcmGd8+lE0Oud/xWMO3/B1FiBUi+0d2DBGZf0+1+p0TZHH4pbMgUXnUj
MQMPcGhArTKo1KYGaRzLxYymQmWwDEuu8Ko3K3ZXSmfJjo2IgrD5yUb7lIBiZd4RgCjfPheKKdbY
n0Y0DgD8wOK77IKnEUrSu1GPUVXBS+FR/xCnwOJ2keSQOcpbnmM2Cj9cFpjFY8fr/bZo8XOAmVJO
0LNBHFprYzgOeHvMQwM9MKZbEC835uMCQGJGWsF1/cTIpXYK0pt/7Z0WPqa+0GbfGmJjCuLc3NWS
ZNmnsQvcUULtsA9f+uIDZZmTH3n+9Nt98cvL6UT9Kh3LtSL1OYSSkhrhyrgp6ah3PgDjHXvye1X1
ZoJrVajhQDhOs/ejRG6DprSYOZXKNNp+mj6srBSZoBiGipzrHm0+X95fJuJFHfhIEjq7hbKwlhOw
yEKMV2zo7gvVrFUat2w8Y+VrGJX+y8b89/c0SCNylWGl+riroi42hSoas0E1tf0E2RAKh3ZoWb0b
VInJhN7eoHwQnzkXTfGvETi0cGJlBOfcXvYSQgTg0bh/rytHOw8EDhQGmkdsIMIYIlweiQlhPWVs
pzXCamWO/xm88Q73Y8A0MRDxrQHb9zv41AxwIhO6En4ofPTqI2pM+IZstSrzBSpVcgqdZ1DdkRMI
9HHcpyZLZpzqTJZzkpvnLH5Kdug2CkFUqtMp5URyyZh6c2rz3FQ8iIlmzAkrzA1Aa1fu04FNLnqd
hUpzX8gNhxxZ9a8UKIDRfH3PPILT4R14yYzLhDTIDciUPLkdYR7rqG+/Zkf2/TsY8XfH/6IqMeZt
ugFCOEQ0fOezMbgRR+FEInWXRlhLQRiKs7TjM2DBj8QPDEIBcw19rieIOJLOHToEGRn5fs7h7gz7
uNLR89fowpF+humyajGe6u7ux6Uf397X3oPPX8dt4jHRFKJrD9CC+w/abr43wt4NmcJjd1XV48V4
4w72SeQzZFuRbIxeHNH8PDwNtNASciFwTXw6gMsj34pQ2fXKP9aqBOemeoj27iaeDQSQbinno7ri
Jo45mYEeURWbts9eaHwcQBXDGI1eMk4bNCEWJrhzpxOAXzxJ7EBVlnfcdgsdGr71VrtqqkbyMaEG
9YdpXsIbnRUSRk0GuuYcmWh9QHnktPNKJd8kaQjcnC4fhw2jjDDY5jxrDgEra/1RUYqJ0+lNQe8H
aMGF7r+75/yFctCIz6hF3wHb7GGYB0jcByHp0+oM1+yGmgJlp3kwd0l2EAHr+KOxyHmYWgxeYJnN
EypVUsUuVU0dvD9Tr197zBPQdiEup00i/fjyamd4AUPrQHidc1g7oigshsHjyIqpbBesaPvEnhTg
KjWt60xZItlc63Eq7+tpFv6KGYoEGI4tvl8EZ7KbUEkgyTV2iHnFUB6Ox2FFjeNihVmMx1xWnPtt
utj0UQQUiS9IaQenGEnIktgdp+E0RoYLFlv1zAVLaH1z/f5vP5b9i6QeuTsH8XzWlB7qiAvZTuJq
6wQ/01HgGVhCJ0tuhbL74q1EKefO9NJBk6oYgPqs6SSAJMXkxByQcPS5u8f6B/ubnBxR2paHDun6
GzlD/qF2hC143poL9Pu1RmSEIVzx3Ku/esPWVfet8j2UZM2ijd/B/9YTEV5ZxpdZx9YJOQUods1V
KsyCLgQ09UwhhTop8hOT0aLdtVWlNS/ZCfKdqI0K8JctSevPXIciB0/a9TfVOzdGWIEEfWM6Wskt
D8Jk1MOJu0Z2pggV2/pA10VT8TbbptfgBMKIMMl8it5DRDozlEjwl1s1yBkjXtCx06OiQI2Ju+cG
o78xGGQAzHBtxFRk/5oP2Z8fNca9yrkRaYdInFoYomORmH34/S3/sVD9ZwTX+JCBwuXvnpV9ky3m
aiy6+v+Q1mB2/A9DgjcJw06VQ5Sa6xbg5bIBBc+OyDBXjUL9AmyI6uFrkhmLe2sRG4yv451+cz6c
JdcJmQ0Rix3F7dniz+TTiEOWPz8o61dDAwkKVWg+kigMGt6sUjefzi9oFdqwpnmhNEU8zKS/uZLz
dFdneYDEXcAmVwwoNmCgL0ozA+suQzxgtQEnNr9bXW73SCY702frZ8Tb7c4MlcC/tOyP4Ty+3NJu
9RgyjUCD7F/fq0iCfJWViXw33L2zcvSpdzhIsiV5/3Yj0uJpfuvRFMp0UyUt+OQ1fry1ebOyZHdm
JaQHhutuP+QuYCVkXJusXLBUaN1TpIW5uDcum7FNPU+ZU7ngo43C6lHzB2lzFKGIj3K5igy0DMJs
FNJydIqnG/FKw62YpjZKlFy7jS8ykoN2I6OBxCY+1dePIFgzewBMmZmONAC0vhKoJilx1iZ2Ewm8
RgvCwYK8CsUf2ASlqeigj+m16q8hcHn9HYiGvSDcvzyQjngwWP5q34qd8FMFl6Z1G6JX7+jgn/kU
mshG4N82z8mNoPzxnwDD/t96WI1J6wiWtAR6HCAmLiqKf0z26Y0BlFWm5zKvc3hgjFgbQF9CmjH9
QsGVBFPKNKfETPICq/borJsSVPz62tGLSoi702pwev1aru/oAQnOgpIC4zM29clMxV0jdgNjNuMM
e06kUEjoRqxY/G93LG1TiwudmGwu/ar9uMxLnCalgkHRSXSZIyotNin+4RrKVnAQswNsD3CQmAnS
O+4oB4maFPXhX6b2IeeGrCgwa71+TUIg2KIe/zKKzarfBJpK40f33S4UIPqcJe2bqUU81TOIHd3A
46Ma8ATwldPaH5Zu7lTVvSYUL2Gt8bysODPO26wfSuNgBZ2gZ1+zo4DjjyDZ5i8cyOWaGh8A/rKc
Gh0UpB0J2cpXwnbUFKbMHY2jS2NDpZp6GaWcn4N+bggam45PdJlI1YTXwBNp2orMToOB5e53k06s
Kl0RXKdl+nNhPAN7qA9eDAYZPmCyyARI79SEft+DZGTJ1ywu4jk7/9lcYBFtasPkyz4dGEELD5RH
HpMpFXr4AcYgfPRxaXuNszg/ANzISsijlhC+/e6y26PGpCgP6WZ11Lm1L8I605pxvvx05moMqoJY
3TY4osrcbdNgbmTyZ9Bfh/Y60rcKHDWloHiOv+NK7q9zBpBIguE34DyXdkg/Eb42FfvCrqmRgwvx
Bj78qBM5IhYhFZaMFePG7uRxbivBdGewFF+aac+a+IOAUhJji31e7IDLwHZlp/iaFlvt4xgY82Hk
QRp+JRF0650s7GQpwyyedkVNxheDO/aFviJRqiFEf71Y1LArmwZtrdFg1hxzmW2VTt//rtY+cVVJ
iaUEuvhyFCX2eSsCblyCisoGxJ6hGcfk7QyT4SQ/pvY7lNBHnAW6sD/NxHVAlN1sUivwcGvMgfNY
/vYQuduVKh6A16FVnIwxvKUQYhOPgteKnTppWdwy9bOHKWuDWY0YB0LSCDAhiUYUWlspt+v3OFqv
++ilLyAzR5/Q0BjgrRT4NGQGSE8JquEKBrtIhwDo/scv07Lm104aB5Sodyinjlo/7EmUqME8YyGT
RBhOjCfpMV7kkNw42xoSfHBpglu8N0ZMD9ZZiVvgBPv3MZvfLJ7XaSnsyAB2BN7qvUODYtk2dBUd
bQN5zowL5m78FOxHPwSMVP9pDs5gYYCRCNnw05vkzVShLAXO0duvNUO7m0C6kjl1Q31hRQas1HoM
jUvTXoAv+6e09CjNfKPRciywhHo+/BgJxyTf2RiGc4RP1dgsRfoKbz2AS6a+c2cL9d1l21Eontvw
Qj7dN9RzWqdV5sirE9zYpJnb4iP/b9DMtoUo3YteQfxqexlmxHNWAjCIlR9Aho1TJ46K0z2eFkNR
HAmvYCpeT4AQia+A9KIgu+qLrIfFkNt3IaIwwpkdWQaB2JDFS2DweuV8VuRgZRZFNMgYuYp2IStI
1kFbnjI0D14HqhegHPWT+Dz99swmeyDYftrWWZcmw4CBorBADHoZ6LIELZ1wwjWixFkQFJRR6wfH
T8J5jZc30BplOwzsSX5ZNtZXIjwixHosCuDkmX7mB9YjXYXorrWRDSAbt5Jj7QGVZdjvmXc7IUAT
kJ6urNtdlym5j6T5BxFKG2CAPht3lWPPfDabL/HKyBdeZx8u8tXz4ygO1ogd0X4FOFyLcXXHACMP
Egqf1DAlQ8zNle5K5j9FOhceKfQYveFioWgZeYM9pk12u4xPUoMUQx7xc6GtuMNtsShdm5Fb+KnM
chEXyWVN/2ZbdX8j5tDtgJ28/2QYwp4kcIe06w7GHcROKRgom6maWEc9EfK516vrRxNDdw0AQgxp
JpeWGZEFidmvxqNa33nAashkMUqQFkWDrlPEyhlSiyCFIMzpaAsknJ+3rQCIn7Lt4TNlJwNCglEG
tYSkdu1aED4XAFm3JjDYmopeA1O3KDzwRECEF0TWN5YpMsuafPUrAU4bLOPy1SGGQ/HV3nN0HM8M
gOZEmyKPmwSj+Ky2dAEdFJti7yib4oqH8pLasLCcat9qCz/iCMH9XPFofby2JS5NrFiSdFFuvLcJ
HpC8OrFgO9/1iruXsVhrf3dhB0zjThNFm/+z8H0pxl4NsbQ+N2K4vnawt4rvI7cBLblEX29aQ4TP
S/gFRIFl3BFU0T6whWwZ3bI3rjYGiq5y7qldaZ5orw5P9O7omofPdAbJgw6gJeyG7nnMMkMK0nI1
gR5Ac4l4WbMYMRIriAHPZwoUJLRx7sHdi7qaDidbVHwWDs6hcXRba9xUIzQDbezeFAStP0M4HNku
U26nFG3Dpq6Cl8ojaV3SFZOBc+YWP8oLHHN02Ck0i1BHL67KHxDoKgsCINP5ucLwSyTgQvqnak0/
SfUWE2f2sQdz7ciJEN4R49QN0byVNiLYlmh1BD+D2ETi61DAQMcRM/942eaeYvbyInW09WtmbbzL
9CiGMZVY8qnw3wPO2hbdwvepsCw6L7p5CtzPZLGe9ZeBOJM5KecUY4Ah69hVUgNY8q7mlvqcdkPA
DoIdDuIaN3Q81nXzehvhVS2RSVcdfiBNAuPg0QsLvIfoZ2TKAlaRnhvHpXwx1d8kzfFmUuIFfijm
GsbWxgBw0fLSWrowXPVY0IKzwiZ1HM7yYusTDuF4Du9Y+pWmgvVpcN4gE1uZymyykIg4bozbiH9H
c1ORgam4Z4JX1E2VvBFtrK1dIakYBDV9ek+RjQsUe/mFhkoZ50hqp5VotnMMf6s/DrHkHTRyOAVX
F2mytjeJ5k4oaiKCWUaCcQYXewOHv4QuMG0kB54KB992jbP+iMGZkMu3MNZ+YrfJvJKW64G/49XR
BHut4lMU759v1joqHoYCERgVIPaZImJiAqRJkFlNhluoZ5yJwnJeFYfnbXVrd9YsnbfygkcyoHDE
dP3aMLAlI4YwEqeNx2vAvBJxr4fyG3p8z7xVRsok7DJ4ZeoTsWJbjshELRN5oTy26IeHbtgegR4F
mL8RCmhP2Y7Rw/vylF6fodWy9JyKvxwnwdkDcy+Y/NrTmgq55+L1Pj+tup3Z3S9OQ2SMTrXj1kpt
lbPkMABh9jGwLJ4qHAa8pW7rpEVGFGRE3DS9cqoXDrTuBcuyVFsFz8rsY2D95fECzs7QmEKT8srh
TwQxn4T2hOGfuG+u91kF5hdOsZdnhKkD+HGj+ZSeicPoiQsh1LZI7wNrltZo8P7PeD62S046M+0s
FlmBtzduYrWahyRN5tUlFQe+EJIDSOda168xPe4Tusod/4Wwc0H5T/1C2Fy84BimnWHD6R86RYUz
R1bNmqY63TqS0lrW2rHCr16CgQi1qwXjMiVMs5O9TXRHG98/I0i7oLi9MKUJyC+JPcs9s+Sa4NSI
Bb5VUVogYyMGQ8BWI+I0MsjL0xDiY3E6Jrm5xvZgT7jEUG57wicLufAt9wrAa6sjwORcu/155tME
xuM2q28XDh6VpyY96oc8FQKd4VG5oVhNyGeJlnQNGvCFo0DBS3vKTAWbiGZyteQfbMcxRJL0jaYz
B028vt424hZPokqBUFWme/hY1/7DnteRdcPA7lmi0t0EUrooQD1LZ5ejDSIhD/CVE6UN0foYSZ3q
G3sI3XiVfExiD2OmUTPwQG7n20cVk26aD1duytSFI/NiDLjtXqf+PVlEWkUzLW0wEvHnyGaGCAKl
q2ICbzDbWRqpcVhNybDgwW77VcA7gFv2EVkWzpkxnPNUKmOZ+UfK0CGokzTAUC0zh9wlixuv62xv
Iq1WBIHY+tLBlcZ5MFs0IljbK641yf4v/npe8hYsgRovN5Ljj3P5S+Bs8oQfDNvQb4biSd/f6yeT
r0FUY3AI6ppos82DkoHocJn72POL21hzOsxi1FzG78B67XD7DxDXTCXNsv6Nrztuc92waqLkS8Zq
6ZN50UmCyIGXul0o2WWlB03b+RCJGcSvpyMxJe2FZzR1fysPDsTKJkG8b5NTSa1ncrcwwcA+cUS/
kplWVAZceFMg/QuIwhOgcm2LEJaTOQAxZeCgiGMokS7bgGCLNzMaP0WCUOmTSgCuLN/j+lAjeeiM
O4LTvl2kyOOIRWzm7Bl1S7o0aldLsCOrDon94o8u0n6a28yMvUn0SpsNr3jBrlR/j5EEJkZt9O3s
xUyXokh/adXCtq+1UKHIEOq7RVJy9n2nyDzRqGEK0TBV8M+PeD2ujhmMBpZFmRCr6tW3N5p5+fy8
8OtjPaUEqozEZRk9k9CFv2L1ZvwNtgFDu5CaCnAqJeYn2I6s2tWpYF8RDiroNBIL8y+loxYhhu++
SFYciiTMIrhUillwqgv0CUsm9oL20+S5J/ciE3RhLNImBM+DMpVDrahRSu+gB9pgpt52nEvfXqCd
PCbBmGij+JU6YWbcEDUjjNaZzswLcDuxF4AEbCv25KpC7ovsFJh+B9Slm+rfBRzExbiGKMvzvvfy
1gmRu9RcZ7sUhc/I4CPlhpkelwF3+aPH8Zim6iAYd8O7K9izjXf9XOX1kRtrOYr19d00tGIzEXWY
48Mq2NAJa/Cv27pX8kZueIIL2gGLe8m8fF9SUQ/YFjFjwDrGdIpKv01cVofTcXHfTNe6p5TYzNwP
YqeR68yI5vj3U7TtFevrPRpZRVFbH97q+a/eb+X+iqxSEEIJky3Gk4tNQYFekDSvvG9Um7iVPKdW
73vWKRWxNueiVx5V5pbBWc6REST/K/5LC/RwwkykRtR9el7PigQ02WFnqloX+JGJXNQq1j5Siyc0
uTDV+eBN9yOIp0/JSt2I2ViiSP3HraGS+p2aTYueNMfbSOC9c3E7yMtHDZNc7FTPp7yfnAj0LBBk
xIp1Wpi9ZvsZr3tdMZ/o+AiAjomjCaMVOFnYuIKqVHk9xotddqi8PIP91KxliiF/FxerzPxb6DF8
R5Di0fhjTxWhwmjFnETITOIE6WIvBLlTw8MoFFCNS2uwDQP5Ghm6Eq6E/4XNO8+H37OIyq1BrwEU
brbdA+DoeyYpc4Q4aLeFvHIxUsIfk2nGz3hE3Sj67HAtDZRHuUsxik1iZbRyJt4P3vFhEgcwd/cn
5VmmWR/fOvRwTUPn97QynAJXqNDKFmopg1//wke5zBS7tm12M7vCWbOPaXtH21bTE0Wt+6G5WKnJ
qNyL1Rnf0w69heXHWO2BTDiQsEhX9c1EGClI2VMTgps/XyRVtNLmIz9zbS1bIUDCRHaKqy7xANSZ
YAAJ2p6lrKi6eD5R8VrcAMvnivsNUEgHdwpQOh1ya2dNNPaF8daDl6Dmf3DwETHmuwSDha0QYrlh
6dTO7h405PMB8TzcVF2LxWbRNWPCFZwH2UejAge++IliAZ3DJWMWnHYRrLTOwJFS2uF0HD8/JHxx
hcXpSdEIwER+DzFlI859Lu8gWlODPSOW5CAF4yojCbo+Ko+KBYn6MrUvC3sfqGmPo3lbxgoU9nTj
yBFY2aQ2WwrN87ZtblQlFPkfSESy13kY/C58+3rqmciN1bNwUchyiY2BoBE4CJ33qACuGMCEouYQ
qSWLpjyeQern32x1oq0YPCRXrxZsA1puOcWeT1EWqMl1+oyUT0uY0YgBynijWxSe9xUy1XLfiSlm
ujJRVfEaPm+wD2bWP+eLUkq9Y8nOJmUkuG7sC2rvOtpCX8hvBq/+PhaXb56rK5naOsmkKGNBMW9I
CgdzJecez3YauooPOrxEVBU2ZJQR1tZy0fq+iQ21DuYQmEDWj7QqS6R3hs9F1JNe8tLmNkUpXsk7
kmyYlw+mGrufkcvNg1Oj3emVR3pZNksIsAm5xr55Ar2FKySevtbX9ay/DdqXqXfxGACvfHTauo8B
pjTa2L3Mu7osCBbjI50/dwfAhby1kPAirpBcSA3PcKgaiHtmns0p2+JKTCm+6cpI1JtW7rZYFkZY
l+Znb00dnusKn019pZsNKvy6YDXyNpifoI0KzLuGsp3hzIrtuYVZU4Ds1KKkGotI2hcZl2YSHEMi
w5KmOEY6KQUWTJd5jv4BJA2DUvIGbf9Wt7GZ9CKdkaoDfp01aT7BVU7tRp3G9BUvpJ56wDixQqfy
ACQknz/V6ZzgXo3Q9/0TXt+qpWbvaw9S3ED9XqwmzlgM9Msk5PUHx5LdTydUSTWWD8XGQLZD5EvI
rvyalZ00Phr3ZiiJXpGuNfilv6N91TuYaeE6v09rwn2w2WSWle44MouwB1SjJg6LUeBMvDHlRJKQ
rDNfb3XKYfLNEcH/+LAitmCQEtuWJZPzHus+csZIHy39FsOAP0Ipkx9L94X4qQ3GsUGfsamSPyQh
zPYfZu2f4YjRXzKAX2rYzLHoR9aPyEY2ob3WmsuV6Hxfxd6bSLzMDH06So0K5/OcOZFASUBYMaxC
xPH2PzEqjYtJ4h7Xcj+OEbNr3lUTzsGdy7ZqcrqfaQBRBG66/LfA+cFnD5EbpBOusS1UgGiJi5yW
A3beo02gc93vSx94FkVHSi1/Hu16WctjSGwIhi0mzPiWqDqM3SmekfJctJroDDN8N4vMA0Xjrbz/
Xklx6CC7+lSKc/eJJz2zdQ2bwvvxUitYdQ+Jursb7nxaoM5G860B67kJS48mqy2mV+fJYF5HUSVw
7qcbhVPrxZZ1DhoTXQAg41d2j5UK7EuUswvrP5SPCbK7O+swfX8NH+O8RLG2KBrAr/cE9V4KHwUa
jfpT/65c5Uqe6wzADWp4xJgdCGLHENLJ6V/SrggCp/pAjZ3Iw/xUKRm33SjOVB5QZ33o+PseZVeE
LWE98GNKEKgpNa9mt+sCdChSIiGH0yJh8qj+8ly2dabbB2CvkfTCgZRMJsaFPZqrHk7zrbDBPjXL
eALnGrzuTa5ulLCoi/xTFrGDzryIgdEdLjdDwND+TewYG0dvj0MALj3b3fkUG4VkX2/adU46kntf
5/Pf8+L4RaYuHX2guzt1498yJRCGgPUF40UOlVmsPVRPnK1pzVhu0+NbdS3VQTyPowK6OE4vh4eP
shvrODLyBsxpnZHFQkV0+2sru6AHAFOONRjhe4bL6LVEidb/io/QNA03yf0mQXTsHBfwXt+mwszc
7c6Rncdhk7bnHjIPy7Ogag2MtVr0+5Ij2ymi90ozTf2FgGCFFZCfkggB/4/igXJBjs4ht8Pi2Mmm
aNbuHXVSYfrI9T+KDwTwF8bmyv5bTQR1yzDd6PDyoyqIwk0cfX/iWI8DxwQcxOFBTBiBk582G97u
j0zZWIR+WakZ0JubWNoJF+DMB+MQ0aGL+Kkjis3qHbV/eaiADfMYdo0EHcyealSCtM1V96AVOtMI
YGbEDXEJIWTE4UbzPAF4UuHYiuwE7TfA06VDskp+/Y7It7taZs6Bv2nKGj9n40Oxn36CIQ6+2eQK
pkVo95Zwgrqr2swcnlOATnB4CK52OBvlkiFm+qCNjUxc9CIyFY550eT1ptSKaeYlU27BRjOlQSgX
kJwq9tiZEil4Xs/csR0FttPni19fgrY7+CdrLt4ZG5Fmqe0eoKjA/XvETBh3qLm71EWtQcO4QwQW
ZCn3PRQZ75yzus8PKI+YPyKao/qi4emTQs9qQ05Wx8StPQcJVrFcJQKN/o0cN0prDFfTa6VIS2Jh
2g9J30uB9435CE/1gK0OlGsV5MQUuxzamvQ3VeiAV9kdqrchy2zywb3I6nUPmNW4BeG8l85I9LUD
lP4cbmi3mN3wA0vIMobeNRHFQfuI20fm+wC04w5t7JJ8ximCYKMo0PYOZHPZqqkH7lp/bn0iVyyx
3OJ9SMW4vsOxDs2RE0+g3HKi6VU9M2MCjVqzTakBJHavllmh2/RrBUPnBul5yWd6zST2852oJnwd
KXMttp7akEltoNRJqYhRqhKmeZ3tB5fa2pmT3OGun37WU+6zEdvGTZzBa3kA3KccGGR1vOfk2fv+
x+RL8kPPcjEbGLCDcekN3wOSzvhwefNRCkZnLmzBXC0e/Y2PqBBxu0XIbxdLXqwe+vDf9e8lvh+1
1a+MjOISzf7fqtivnjUh/cAOZwfaKQcm1Cly/KTaV0dtpDgUfkZvG7+GdpfLyZ5FXQOhHbquITKL
LdncWAgrL49LfZf2C9C6VUiU432EHip4tx//nIlHIbz8M50Xk+Ppkz0S6cfFZJG9Ng1U8HN8eV4v
GRURh+tHV9D0DqEYCELqteBH4tNKu5/7DwK0bpZBXF6lEPJkjfd0ofwgaAUA6POunSGuZnLhqWul
8F85VwmzSZYMSK++p0N1qLeVyTW7/AAKimWL2cPkBmkMZYDWVSjUayge6ch4Hc4mt1X9uFNe2l2O
4ygvX0gfjXsX2+ATZ5ya9YQcBUnX7srsjU6UDPTIhCb2lKmgBJJWHDpquuw2OZae8LOwxsCEz/A3
wN1uDe0x5leNnRY2BssYz0iBHSAeWdCgpkW0Ja4Y0xh/LKe/NDLXfTgkRko+A9Dp4Vj5vf4Mn103
VwSFgk+wOTVaShl6FxLHyBly8k+9vrFJe7sq1hdYstxvcGr2rBRONL0ksSwk+01heAP0CwvNoc2F
iTTsbVfZs897rFLyT6KaQNjV/+7noJ73e/92R7iRd/hOPKUs+h+BCqLcluKJcDKkREb/HV203yFo
CibV0umY2mGkIKV+sPC/Nf5gC+XACrg5YJmV97DVAj+l3BRPY86AfQF4za+Yeehvvw0WhCqf0xJe
dWxVETjBhoXntndRUfCJ6AQ+uhuP30IN3SONQkW2vLGhhEkWjptlHwEMm3sdLiV+i9JLv4kottCP
In2xso1xShSE2lSdLVOKheChmzQKoEXdgY60uVUcJkx0XWB58dFYcE6ZZdP6g2YJD9HBfb8MCice
iKfgr6kU4NfYARPnOIduLcXKB97QwdX63zEOOFzQr3D5UwcuuU+U3KpypadPTQF615Dfuq0zYSys
wEydpYNU3HsPixn/Oe3fX8rZlfJhYrjAa67jRrJL8/vlHpYTnXUYCz9uH7FgIaPFjPiU8OcOR58y
e0e/ZQIGgR8lphTD0qRmoHuf2t6BeeN1aIoMxqOEu9rDEd8IGdcK+O0itPTpGqHOXx+igMa500BJ
DYcKVP+L6sl48s4qfHhsRbRywCS/W3gBna8eoiQcIZGKWu/0KkT78n2duXERbyq0HSs8ra9RdmCr
Es+4duAnVick9eMjouMRssieMnajkmpHl4BNw9dtE2KU7PkVzRM8CFfhLw/rOEdRa2wqU33QGm3R
x9MoT/zInu41WsprOznfVnUFxqxfi4JloGiYuND1pD2ZmrWjtl/KBmPAYnPPYS675DmQhHCHbxq6
s3XUy1C5TuoCY9K557eSdW2sD3NQy8LZFzXIW6vxWeIuZ79iLcBRaJlzb+6N1l9Mu1AyClEUnSsy
Pnea13TzBIc40xq0T9WD8d4hhdthrHqWMfxcJJ9yC/h+OLjjVwxK/VvrriyZjhGmL/K3IsTh1ndJ
HXV59iVxqEf5w5e4vHrFifGx2TU/WGeDMPzcw74BRKF9m97mqJ5Ow1AmPSh8lx9jWuXrr2hbWEQr
314nTrANNLVQsEy7AIqu5wmMChMrpuKyfwJhkkajDheTBUqF6kWiSbR0pcnsgBFOstRbVDyrd5Gk
azHlEa6c8P2mPxx1gSkjCCRZ5sFwhVmvwtTOsnougepeHt8wvfqH5+zg2dCpNe0rpTLIy3OkWa4U
5+VR7z1KYBvWO5p2Q3vdYFAb1O2qwXqwJyA59xZpraEXKwFL0Vq5CU6ghJoG4rzRABwL/mGujslt
hGS5t1HE3xZ/BS8yMnDQkm1KCPaz8O0O8kZBcr1uE1VfQTLif6cZ7tLR3JptMVCMBvRTxDE1lgn1
rQNW+uVkzUudnO690VcNLVkI01k3YLSicbh5ueTfilA3FxdJ8tcPVfCim3tg6cASNAaQVfY4NGLV
CSisewBv8YEVPpb8PUOHnzG4HHSSPpn/0nM9LU3yDTaWrM19CGJ8gFrOB2mJ1pFDH4UUj4dctEvS
5O/pwcCvAmyAip/ur+C0Gs8IsT70gY2MikCXRj+FaXVwiyos7kpUBEXOIzlmUSNz4e/PXpnq/KKi
tIS01tMEOVTYCP/vHiShBdxSH7CE4iMv1tYZ0KrqxKvDuJJEj0cGwlSU8bSiXWUKanla085JZNc2
ei7eJ6kJHs08CKQffjlhHW+lFNtNAD5tbMc+mqP6IPzHi8ipyixBWB2gzVVB8VELJpxqW5VQ33+5
XcY47ebzvfytfuBxlC5rYiReVpWOCkGtxrxW+d1cNQJKSj66w938WPYxbPVLerb5ORNtuL2P4RgH
BkWb6RGecdI+QIFv1rslPyyZ7i4G49P9NqbOwN8s7WdAztXa2xNAv1X/9Y42Bag5hZ/6KDtJXg0L
EcBPXtRxiIsKbXXtQOw6E2Z9KypW+8L8b36TNbsrALhYoZuswOcDGgaN6PLMfzIC0yZ+rMJ+5g3+
haISJlRO4nKDELoLSxwtioK3nop5dofMD1/hxlKgeEgPKwH1Ra4TkAg3W4uRBKbXx8WvH01I1szT
FiW+oqqJxPnylzTiadUaNN8nXLfSIkTdxkFdjereAY3oNxfsrRCPUH6Pt/ZszLaRH7hqOHfX+1fO
Kepa8E/EcXF5OSXw/gLIHTy/s2F3cdbY6ANJpqFJXOAMeZb/6+C5r/iP+ugPPaH6KFcD4smjIWsR
LTVbqFBbZNw+aDbRz3ife3QAdr+wN/R1bjv0z3laRUuHtJcK+6CesrVPHbDsx1nF12xBU9rWMgpx
qD6+lX2LPotosZk5LL9LhiyPpt/ySdJM7T4dYTP9qbd5fWAFMDPmPZ/v94WoftXXyqEETv3eJ8Hs
/nBQ/vty/vuu1X6vV4oJyXLRLlPz5jWzeTVNR4tVrfTcLpQyU4o3ynPy3C/G/PzMGO472NctLBdL
auHS1oi7Zw3D2Trp5NEguPORyGsaBiCdJVC/cxfyEpNIcbq61ZHl8fnB7CQqFqgG/YmiXPRIK4Qs
aEe7mfa3b7rr25tSUlJh5LT7bEUtDlwV0UCwhv1SXnrmn77dTiNQ0xZsO6RgjDSwKpd2QlVGAqHv
MAj8DouyCkBsq8Dqcms1nAXS4t+c6RlfqTmf01eSxdY1ZXkr5wtrh+YU5foBXwhnkdw3LwqburVH
d7lxjuLnsqrhj1OGTH4qIW01JXEZHDn2G3UrQFfBKlikRKrWknmySBCfpNUwpLaQ4A2jXZ9K/ETY
hdc8vmTcpX1mlGaT5etBMvNczym3TOiz2f0sVkfIDeYRyNJY/mjqMLiebGF29T0e+RY1SApDdJbe
SZn74UBLFWZ++sijr5fQIsoaConT6eZbTfyMe5e19qBvpVIbAsKtNxhQfnr3dhjyg2vdUtdR6DI1
0N2RCGX/+b2ulrWrAZSglpfEFxQMsZf2Juj8VwPEKGBPN2KMbL8dE8c2/Mnx8vt8ricz+sexDhe4
oBNPqgHyJegOi2VgHoO1DokXVniOK56WdB2sSu9RDdb96V266s1orFdQ8jYIc/nTGYIbjdscsbzk
Ect88uvT2shcG2jNmhGKMauiiQwJqof/rdybHz9yT8AhBWC7SDIJ2MsRHjGX0JuyaMgu7AQ3xcBj
YnwmEYbP2DhsrAgJ83nnYAsDpxOyi7kHuXWFt+f81tgJl3JNJqY+68zWBXrkEN0y0AHeREw5tNe/
iGzjyQGRWrVdg4Th5WQFhVI+pwtz4+hFiz+3aSuZV8ksp0O86HVKgyBQueUWE/ptte4XcCQU8r+A
7RRJEc5PWSAIdY+3blOTlQpseb3JWFxiUf2cDcaoGA/EW2dyccRuGZOFFj3W3rVGcgipjZP0ECIW
ugRuV+MhBLCIwkFKTiUr34G9L+2/auBHik25ijEyMoX+wYZ3w2UL14X02CKtd7ArQqGkrl9mfBPL
ed+zOcckI64nUy6EqXPDoInPB3k/i0Mea5lB5/gESkZvR8ZvWhj31AtMXso71ZvIciREj6zgslFA
Gga2HFHHtykRqEtBFYmLSH4tlXLE8+f5X7fLNUM4ZmLZ5fFY7MbESQfzmwjQoocFBy2w/F5Fc0xL
tAdATrWlPeBVfG8acUcE60/QiSflsJKzj04+Z13V/AAw0f5NX/TEs3SlGBxmNbOemqhL2BbFeMBn
Q8J9rvvaOuomGPsuU3vUC6n9p5a0yeJqpFlF83YawcBp5Br1eAKMumBJg21Sa1SHmGdT1fViBNqA
wqLbqTv4ZZMq/51+8FRcjVr+epgm7h0UyV0DmpgBmcloduospZKkFbQmBtNtwZ4bbF7VC1xrKp7f
0mxRXFwc8tjoW93+USF/q9rr8V/PBfb2EkYY8ExDuBkDSst6H6/TBtlZwYsUAYLc3ZTeV0b1BNxX
n86MYby9YhvkmbCPm8YpLM3nzlyobaU2WTE7FNIW8e5+q47LS0gobMzdDbudKVRFkIKUTG5n2ebg
8ivYoepV81fF7XGmqrRR119rSF1Lfz32NRX/ffqYYItm4SXW02uUnntw1znya8b7rJdONa5F53ME
7kxavTLuwcTJ7WaNjRMmSCbdPveOcdRX+2PfJ4zbsvnyZmqsYJH+8q6HNx9mzvpUsA0Nnf2KnNgP
CUrNYJqPUbyuc5OcGRuSh+J+1rmWaZzXRXxT6gdK3TbfJD+6DTfQdZu/PHJkR4SHvd+G4JeDxmU4
dg9SgoIaxFVGexI0nfnrTVD+HvtEjBMriCCWfcTTwxdVE3zgt5irQi1UALuA0hSW41S/KwpzkP36
A1r2Ekqfh0NMj5i8lgJG4lkPnT8lY90Y+nOz8LSJ7mR0skYViMIw4S7UUI/WjgQutvGrJTl2wKx8
k+MW2S2pruB/5iVFCJZTRTYz2tTcyo+vbpFKbdp5LspEsLOhD7XrOsI+kOLtTiXPDOsBTQZ8s/Cn
NEGSYVhO7j9tz7TTTn+wQA5a+5RMdmI4D0gj/vNjfViB6MlFFFwtjy1Y2BpIc34bRbvbg8Aj+uTF
Ke6q0l8bqBKdaYwxGDWOo9R4s6aaxZE9kuY9bqde+KB21KlS2LnHe1WWsplGtRViZ3snAL1734PE
+G1XPpyiQbdK2F6RVU4MVIIEQvcZmkf0SRtbkMeyxlc9CE2CCrKU0hB7era3Vx8uCX8rHJZBNlTQ
GY389JRFXfG+jtwEKD59atvq0Yq5VF5vRLwQ6qvSYQxkH7ZRb5aPgCL2E7WWeEH79DR+3I+9Lqc5
a1NWIsCgP1MwQ1+Asjs8DfPdr2EBVL2jvDMtcR72KX6T2e/WIChYdKKd6xCAMvHzCGlOYHZ+ri/I
ohIROIrNqOY+LYXCf8eAvlHgfVOb+HUnu/NzuLL1oAf/qiZM9FHXhmXmNBnRhup4llMwuzNp+n+f
Pj+7utEc4vONV5/sQohoVFpE/85gYj3eR0fJPK0a4rxQ/DiMzVNi38VgC/1tnBt6a3T1csynKNqg
fwjLgevGSghcFiOahES8GaX/s1/lJdy1T/nxnddXhprzII4RaikVwFO5ECB3YRn3mmgRqdB8b1GV
kliv/Xx5cjhmQhpbfFWdrCC0b0K8hSnhEfZzQlPDDLigBPRcPdhWKg2r810g9DxBT+nHuxW4vBf/
U7gA7shxDKvDyx+S6Td4ktuq9Qpy0mFhzfUmaoVq1wJHNCwqcU21dATTgTBXqrLFO7AWmsn+4hCI
c92y/WeLCjOVaVaxl9iFnJXdDh12F+P89SGgE7pFh6jV75/rAPT0Xr+zGf5uLg7P3AGe0Vz0mX3n
R3UqwqWY33JALsaG24JyqTCmeBbHbWWRyE6bYrTkMmZzktqIAC3FrFL43xlRNJNY+11a1R6L7aLp
o69/gJcLzq9DRstGvrIiLGGlm41f0Gd+lu0kEviZhOBkq5jWGnaRb4OqDUqaJwyFaOhoP/LRTSrM
Y/r2YUIZ4Iwqb6gPdXbo/ZAwgwH3kYLNv/sJBmh2pADGiRMapzQKtuC794b+QhUsXaKc/+tbI+3B
lY9XoWWGrKTUVUo3cnn7clWz/CRbNnoXPXZ9+2QfGShSWUcC8sBbUhqhbbqDjBNeHoJJ/4hg1UCU
yd2QW5yNTdOnsQVLHtlvciSz81xwqqQavuGMw46hE1QoY8GCgyQhHzempGbvS1l/k71qM+l6Tnvt
ghmRI/1eBzKX1JM/36xACu4GV8q/JQ7i4sSIjzuTW3+xrBk2XUBpwu33nvrX+/v0HQd4zDzBMvwf
q4CQX6fcz3RvxG6ZoibX3MajO1U1jyFsWaLxT/LVpgP3nQs/whpx2pFaL/EsX8B6p1Dr9KdjfVCZ
k75Q9wT1yBFE++lCZIu2JylEeIEUypO52i6UdBoUHbOR7NuWc1h9DtW9KiNYR7sfWRqVi73ms324
8wrtNpWyQHeFfHzTu84IqeEU2E6Y52MLnRyjHQdcYur+opOXZ1pOdOUSV/zIGeCLFmVlCNt8xjQl
C87wcngkfKZ9W9+UhLNSPthc/J2gt5pRgxcZYmOm4KE+hoqLJyvIRoqyuZI9Xqw2rsSH9MbfLSQN
5M5Aoq3vukAYNFoqkYF+VH2y5Zg2lMnqLER6SysFGdzfs8ZnGzf+qCHYpQxDBpFvkhq0kApj7yFl
ZBaJ7jUhL1BrqKY5zmR5eWzqshcy2ddRvufByTaX14f4/BbF//SpXsxgsHmVIjg8H91svI4l0rXa
dTKwSdRBVlive35aB0AZKAm4cG2eIx7ylHJQAlPjFWxGzTgoUqU8Ie2L5ZLN7gaPoA27vr5+TEtg
rfax2gmqIdHukcB6iMA8dYbVGefAAKyQJCnvzzFCeKE1VYDdrVuW+YywXIUorUjLgKJssa88zoMT
+rf5hH52E1lQpy3FgCwum6JDQuf76VUhpOO+Hw7BmOEo2iSkg7NrhIR7wpxfTWSxGBZf8u1sV5w2
ELr4jTvA1g4tp0Vd3BSAZvbcfPJ4x1f8WZ5xx9iEjZenEo5aSJYaIXNuMdKK77SejaJtI5L2k4eT
Q45RTS4+pErxLIi0ZTKIEDaSYd4jUXR2feTym2Psnttyl6udGs8GVXVjQ3p7jLfxlsPQ9FUgNNvz
zwC4wbZ5nzJfSGt9V3K1ffTXVrTcQnRrmd5jCcOCfC+yoOs0mMSDIGpfBgZ/UidFVkd4X8CUWyqK
4rwuz2qhbLfI/9o7eHH77S4C4NkcZ622hrcwsHRTYQSyiePjJg6OdgKbE+jo0R3NREdC38Ib1lZs
cYkYmj6Ip81OALu28W2jgSCAzJAm8TUYVscMBZOpHA29BCpgZiGU+MMiEM7VJ1BbeQHVP09EmfEy
sBq+qpZG12UGWLs1brm2WYckZNHVGtOGerw2IOCrPdpXaMM4JFOdWPSkL7fSjBFMyHTXjSz3HxwL
H4EbE/fe4Fyh4dGJ57zWj8EVIU5CRVg39pedZyCknL31+U9hqarcSM9qAROT0jPoV9yImg6gBFLk
xliSJlSbUwE1HB0Z5P8c2cBFcMln5oAwUx4YUIeEBHLAW3kKBUHYKorCZocFX8Ujwez9hlYnPvZu
jn3MAIIre4jmhprk2xfeU+m6xhf1AcYC+6iKu1GVnv6XGIsH43XB0OHDMEfAtSYdWgg3cut6mABk
ineyb5HGGCI00qtCNVsFbzggj1S/Dgi8PL6FnFFPSL7UfF711XSyPyB8KhOGNRNUAuimJUh+Mpkf
CnsUbI+N3TkT168pBieSPcKZbGk7C95ZVgAjhlfvEOARA/M347Kff+Y1P54Z5yBu4ku4rJM/RxzI
KfvXngAJMWYPhhbLHD2mJcRkmCTROPa+SuOtMpilekQ+CnUHzfau+F1iN7op6CdZDYRlp0xad+qA
AXxx1hME8Gqpy0+IMpcklKUSyW1EENBWkpjnCj3KneRJRUZim8c7kWIg1qAAYa11Pl7u2r+f+6U+
By7LANEmtEg0KAa1jh+NgD4GFxAM/nNQ7U4e+xr64a0id5ozjaKSMedBBkjitccyoeEDiOLo5cby
nGJi40thM9ClZftDBOdSxUetYJrCEyV64VPy5tIkNsbQaHLych+Qhc2ZZ3dSo6Z0qDo8FGWUTLlx
QK2s+5bV5rv5LxPuWYqDlVldMfCAB9rQ3wzz2dh/OsLTaAmlzV3/IH26iWscCo11amv80928Rtj4
L6855XUNvJlbP1euLhbOW5/4IcND2mfFDmvrfjR3JVK6TRKZnMA5Y+43GQQUMdd7Ls8Lw0CR+u9p
iaeOuoFVTpphiNMwjAN38/dIkpmp0+ZrMnGSic5MR14cQggQSLttfAAwlbFTq7HiP4EVBP9WT/YX
CIlfOX5rtDTT0j6t8ieF1oFkNmJdKaKKv7t/MMpEEGNg8Bp4sSSlHA6jaTUefBrzyL/yTFxJPFfG
asR98R0fNafyI7JbKuRv3sOxtAyAwjnzDgCJdCUQc23tJTe3mdIvVeg5nA/1IqkWdJwJQwHW4zJ4
Gxatbqky3klh7hntU8cZyvF+EyyKJt9Pm+1m9JJupvAe3Mulmk0oKsCxks5h6Lmj1Ut2Zx9QFZag
w+E4q9tWtiAq1RGb3UH20abtYTCT1c8htUMKGtPRwjTFUxmG+Ob54rDoNY0gCwbh+Yfm7J0iR7u4
jFTFpwW5P35mRjUpGlHf5d7+U8IgdmuPt3pezQIvRhDWvWyMuDsUhvRTGTYbZ3m0jecdD7pGx1Jr
SmYR+sebjQbkMQ8HMsesJdBIkfNU5R+UzCUpyaouoLOt3MoXtwXOOQPvHzTubUugT2wHMb7YpuqA
Ury5gtbYlye2HxkabsLN1NAoPoxnHBnay5SmdkU7P4xJ6H5Nxj2roHEFLflEw1+RY/sXIHO6geaf
nKskMZ+uppY/u9XUgrMQvZLWafGY0tkSB0SOx2hY6ly1vN6BMdwt9mFSYhjIRhNRsngVaYgmCvW6
lM1tQ0luVj6nL6ZyHPgu6ORN7E8hmZp2gY6Pn6djcPP8KU4+EPZP5fH0ZGnWwA9aPfcB3S+GTycv
ddGI5Azxv8AQes6hFFi81B/QRSR+QXMCgMDpNd3aJOn7Mylvd+AaVPTVq1nBRRxlhfSB2o5/V5uk
jFcwLgQlWNdFd8xtFt7uPHVPPFFKU61QBqfQEOUtz2p3wcrH8/CJ3TVzAH4flUAd4Ggdto2L2sds
3/7CpYLlg1RfXQr0tgCFE/SvT6+pQ9KzY95vn01y/6vTeS8LGeGAu5UNsrBUMyQaY7WZTrCzPpI9
RRdyYVH0K7ctJ38RCPKdLQQzZZeofHz4Tkk62yeITJTmHw/ZT+34/2Q7VqIpZG7FETjYEQSMhKh8
HG2H5cbL2gIQ5iJ1DOP0L+akkC/3kahPqTdv6qniIYTFDpihi4ydmpD2OSJnIcEIChsTiTN3RDpu
qCdmAzrOSj8Z5afKQduwNEGfYc43HgRY/6EINbyv0TouuD7vXab25xlNYKT52mdc89CjYKSMQBqQ
ywXhLgulAvTmRXnamynoJv6MuZaSYnUKbCptVvcbQeiKI3DXL/er8vM7z1Zmt5Noj5b9Lj+o99Uz
OmmOzqUVeZKJcwekOQzba3Ghq1b0Vdpee+gssbe6oUz54O0qSWbq565gc5RgfIMRTyV7dVwDV0iY
drfazOLRP60buE9xCXm9Wo8hd1GcT7FxlYjzUEczb6yP7FVmuY17RDGCSR5C5YM+V9aLp6x+tvOF
EF7pz1C5siH89lZsCp48D1y2jhRSCJMlMNmCqg9QE/vlBdPxQ/hpptN2PMuTXPjJI4WpyakXMdJY
fOGO4GqgZuZPodi+wFYcb/hIiELOxFuIU55yP54qiFHfM6g000j8dWnWQf5YAUlHlhWUqeXwWvIV
XXHbDlWPmbVjg6ksaN1LCNkolbUbF875HCs50siXON7mJbm2+ek733WgdjLAa1JjYnYzl8hvQQPg
Pu6czuqmMjk5IYY39thkfI2s53oKi2oRLYcTVnRAO0dhamKJJZoHPA0IMwMDoR0mqcquDKehWyHC
oiPXqSAEk1sq6X+ft9HievaGjVh//8zapqRSRv5n7KOO4khZiTI5kuI7VYG+bOfPs62nBlyZ+czu
cLTcywVxuuJMIfRxdHyyBk1zNpFPZCtf2IaI56H4jUbgL26VkVc6Ann75tOOpuTIEuem8x49M/Zi
N6sf1qHaJEFLqIzOsJnwoPvPDFBngrMRuph6WFPL84g8gBJQEnwW79XyjzYrnsaED70H17brgfQq
5OIBxWz/DMAV9EbCLCv4uaNWiANtF8GOPxx1MSCgbci5VngCZUPeIJ4hbA4FD5ZusOHQ5lHIdy9h
inlUDR/cqyxt07pQR9c6g49ugI8Gi425APB/6p7UfUBQQ8Ur2K5WbXJDbAl+ZuQsrexjnJypM/su
5iH8pMlDUCEFHq2os8QGVqeWqz9LMckmBK6GFqdEdoSa+/BvVrmJ/VMCysVWPCFM1Bn3TFANLxwU
3gfrw8QB0OnqU4vQ3O10m16LPpBxOt03Bsi/+VM+1wFEqWGT/2W6H3XDcpVeoTTxl8oD3A2kksp7
W9hOtx6Gbzb3mnM1K8/eBbeONY98j3AkEZuHW0jwPSC4MpYSHun4uXS1SXyn+N04A4I9jcwZHOK/
aA176nfqN68Vh/vvTSqfCo4dMADT3b56dn4iyoGVZANFOT9HQUUGKVBRcSuxr1QcEOoXmg+o04Fa
vE9YIR+iTnAJvMTd4yyLbHbN9ggWXN17t8LIjlWdPFiQ4FjaztEBy8D85Knj5yVpCfwobpBy0TFn
fsi55DTQsJ2b8SerZ3BeS3bTJsjFrh4x9l2R9puVgf+KKaCpgTkolocsIDFXaLOTbVNKJP9V5YqK
3V7sv1B4KkjVaNJRlXk9pe6NCgC4EWCOzWXBEZjaUVgR1SMKtKl8xHYW/zatTKl+OjPMq8Fp57oO
8qhIISJYh9P0JnMRQm1ghEcY6gz7DPKlAJRyQ+j4m3Vw0rSk0eYjjMUUk46Y9vtl1v5lybVxPtNV
vhRsK6GMMAFd3sMsV+KuxzfqLK3vXYTQbBVX5SGv72TyfoWi3QxBqWGjSUtSeLxl6gg37764Am8A
uJ4K99YsJE9QSpH+g1gq4BdS+SWyZejiauaKDysR6jJlf0uRzfuCn52ETrLrqQ6AfoYEJ5DAusKt
S6Ls9OuyHTNgFjLugdiH+ypqAnE87f3twtKSMZJ78sGCu/jDrvdddbTH0b76+8s+pZx24tWWbMij
3sHDFkFN7oNJ4mQOC+mwSxd5ketNQH5uWlZD2E8D3oABUHVNNEGfUNgrrIoc5z0Io/8zJRMMZi8I
G1jd3naBnmXERZCDQtIXORqjdUPHD+p0xlSa7kYGKDehtS+K5XEsE92kTlJnHkehXg46r1NfE7/+
pFMoKyG13BRloRGdDlhZBZlft+6PrqBFiCDg6dNW5kOHZEd6M7JcUngz6Al6gpiDl0UggpPjqoN1
8XRWnDo+NKpmnkmbedn7tTwamfChm+jtUxEDcnE3E6HAWMfYyogCKDjjYiiLMd3tHD86J1jPXzvn
p1dByFgmjMD36A01S+r69ISpSVkwzjz8pasah5nmd0MT9rD3PEWcmZxya9VqzxMpSvN8u+R6Dxha
4xrQ92mEKhY16fqQrTDsoy0aD4i6Ja2vAZsE+QfsDhMdY1hAcX6+WASMx82roBnKydzBxhuS2Ljj
GqUkRspo/RX739FbyTQQdC74izAKTEdgPu5jPah+vaeMx7qZXoZX9xY5N2vWSbys6BX6oGphmbl/
ZDFerUgw7QhN5o+Zpsd/d9hKNAqgyFiQUU0iuMzZQ/+ajrpE2SGrMU41QECvSmdlJajJea9CNXYF
F90iIgRYyJ5DSjeg2hVJ6v/IuhzRPkqJEV5U1lZJub63wefiz+sFEJnLBD9N9pLLK6tbkrx0cD7H
h/7JWphnnvaMa24gkyiWekWwrmbueaNOWQJytNrbro3O9qJYJPbV6xZkfxOH0HmTnPQBBlNXC0nP
kiYZBdQI0CoGCKS5jk2ROVgh2v+rI+TYSVxgfaQu2b9nfIkSay4pHNK4CaO5l4RWVjUqJseUW3SN
Z/hSPqsQ/E+yHpv7uYzPP/2r5Wyw1z9ptc58lLmyghEhWG7q5JzC2URADTf+NvnUrEWkYKw6QO1F
8x7GJu2J+urxADewELFlbKK7RrWivXTGowKjk1VOcEdfiuXRG8CbnVoktW1X3KZowbbizh8tzH/y
dy/XPTsnoitqKpRcsEXgJyU8pEPeVNdB/pNVgYUhZngFLrhgKJ/7/HnyGNzev+XFLVpC0zg6X8Qg
wPeqzR9qpDukrbaJSU0BWfRbUrp3gpcL2Z4JS0+USpZpRacufIDtcBp5wCSXn+AE6dxPPAydxjJX
R1WtQCkR5tX0kVYAuailt66UyKw29nrkLr97wV9wKzgrhhFJTPBt3ZdW8Yy/BbUbtgXSHmaDinf3
ccZWUe52TvrmSns6rnOzW7mclczWTDX0WhLItrec+yugBN7iF5iwwNVdMdA48Uj7jKY7EleTaEIQ
MLHcntbXiwsQaLKTyqUNv9oRcTc62S6HC6SQQoc2HLCBlYkrZdJb7AV0jtfbJtbtHi9grnoObtFP
wq2/DeQT4LGSqum84xNvFtoad9d78VD/fHySyhkxYd3ZksRK/Tv1Rc3gd5XPkGpokdOI6xGIyQjj
8CPjAcz/cFSBZTnbnw9iYWDqldgRH2T80Dydx4jNxWw0nEQHnz1jzWc6H5vNZsKmCH3++Jn8CTp/
PZjfnmff5wUACNmkxNsb3lVnVIxu7qxTD6x4uSWrwMBt/IbWXYg+0xW+W/wkOwXQfTxJNACniyA2
7hPqiwspnk6B8k35eolpkL9IokmEqvDtny8G83zQauxEKkgwqEZWfKe1h595Z8KutG+Ua3y2MjoF
C/6uGFvpFiA1vsUgR6KpsPqGoQscGpbCvVDnJSs0Xmb1KA1HOjQYm/Wrh/DZ0AhsXk0J8pJ9yhOz
D2yo8tK5ZOyZT1W3nWI0JEX2GCHVbpN2LzlY96Meld/N9Vm6RUO+KK+ad5G4ukHqiFEiuQEpXTXE
BqplcCWNXOjGltBVaEF6JxO6MtM9LBGJlMn0jF2NxeT3r104IZBRMfaggkSvUR3SIjhMXF7GpdEu
P1Rs9VUgONvAURucldQZyeUxRpfCq49RnUQp0+c4lr7s4xYnONITrtnVZ0Wgoh4k8gdMbLV4G6U0
GCIBe/miuvq5uQCOXWuNYqiKqoq0RPNIwVXhD2lxM4IanJ3g2tLuXwivwqoDnM2LlVB9d+Iu1NCl
VH194D+dVdM4q8AtwYdNZ8oMvA8ayZ3ggzn6n1AKJcJBLh4Hk3DZG3Qrv60WGlnoq2aAavdr9HBi
xKZVRoWRXgm4nq4H8b1EPCDuYK1onfu4Vwx3KkYXakF4g7d6qEMKKQr11oHeUewI57J8jJYEPN7w
la2Uz70MXVQ8xGcW7OPGZQyzQ6QxP2VeBrKyRgIGujneawodM2OHshiqB7F3t9qb/zmJfUr0p3CU
m+GqPL+a+E7/hsq3yCCbB9ogei6iIIXFVxWT3jDvlW2qdhp+QIGieCsUOiDcS0+T3gdMnWINJly6
L9uSRkrcN6kTR6X6Xw8AHvOhNVdcBuruKKNAJDkkF2DAc8BsCJK1e/1B+h/SP7H8iLPd4+zlyRRx
bU2ARKBnC2JbbsQcJKpTgTVq9ij9ykN5zQ6ikyU02+uIYUsCSk86CecrpcXTS86+9J9Ta9Czh96k
3jw2vb3FlshMoR/KFVCPwSWUhTRfnYBxkdfjbETyuDz5zuaH1xOs5wqZgcjUZy5M9ZalMWikxdYW
UPJiUsqG92mXheZg6uKe2cNIqBOLp49OkV3e5zP75Kdfe/EJDxbc8IOUEzf/95cUl4t9W7OGj4vd
JpuvwqhZsw5R1NGAnbmLr6XkhHmO5e747fiFy4d5IBp6fskN9n9E37M7YcAXs3pM1IgkxDkgxOkk
p3IHft0St3Sie9oJHn7nKRaLw6Co6Z3ZtQbblhbUrdHcFXwOmMnpFwQj3nHAOSlTphbsc2T+yJ5R
RN1+1xcPSyQjSI0X490Ffm2KYT/DHbYQWXrhYBHewsKM52YNCOzEqWRp2Yzj7v60INRPe8lVtjjn
Dgb7uWubY2k31WW5TMzjHrRDpN8e7ApYbx5IrqAj29QR4vkOkFXhfEKTTTsekR7rw8wq/l1RoMBG
e9fZEAAerOeJdCNvOpVEySpjlft0C1OuY5AaJVnp8H4s28eckoWKMbVp8TrbN4cr8JUkBRIP1PTb
1G2W2iX1puOdIsOEOFFIfqQPF3HQmMqpUlIDtScT/wuWs7pCjJv2325JkEorgUslxdgNuliAV8cA
wBcSyExsySdwfF+Ty3YIcV6Ha/lB7yr0qrZ0sMvubIZuJ3Gf1lWWyL3AJuwuOZH+bEscIf4HJZor
xg+RgQaLz5UE+9Ue3IUaiYI+Kl/J2Ga8t11AzbUxo5Dc2ZYSIngorVvJpkIyQaagAhVlZEaPKFTL
Aoyfy7FZ/uj2hLCaYTMKPU8PStGSOTMF8vrehFhuSZzZjBHPE+xvnZoLi6TUClQuEKCk3zR3SyFQ
m2YALpX9uJcYznaYBg4K0Ek2tcuH5aEVbFTT9yWK+Lnfd2d6czPyo1VN6gEAHKpo7Rafz0ugyFGj
m5VU6AC5PIF7hFcnUCuEbWvgV+jHsp/RJ8G+xB+o8s6G1yy6ta3X9tFd31zrM3C0xNUgIbjZjiPH
lCNiGbyeoNYVDBOyIQ6tcPlo5Z46x731qzF58Hm1qGIvguX3WK9XObzUbZW624fJ3BQo0i9Ed/D/
ifzKr/tUiigi/vFbAw9Hx6EGs43NeoQxCrgRLrSPNRwKdCT87rnQ+V1LPkARHodmltO9SEQJ2qTe
9d0BO9fiOBcFPfiexHBj409z9BqCsU4mRBZ6MlSqLPHWHjMicKLqKf5p/XTpxX6W4EarPGCnBMpe
pdDa9sjILpt3X9agfnWFt6pZCq/PrN+eFpjULDFCcy3V1kRC2g7+pkPSkIBmViLRXlcSpWcldQAY
9eji7OX02FtR2uwImwdQqiafy1vGGpFuu7CDf8Qnltda2jUwPfIwX3lzV13u1usI7xzuZiFFwja1
dhjU3bKziYtPCv82UGtxxxcl/nk6RWpvCEy9dYnSVRNYHXHU+mH9v8DiRSug9Ri61bcSn9YpCRtf
2PCZy6ABnalxUEvBy02yE1b2Df6zPrS6D3FhnT/hEZFUo6zKAOvgV93mgfIONkqikiPkFqO3NeWF
Ws0I6exzr2Qkw+GS7d+/JvSuxk6fP8WcDbpERaNABWbbIf9A9zfL1Hrwekrfu36JcG15BSEqHBfq
GjEwTy+Jum7VuL3QCa1i+JQGsR4s6NdrrG82BSLvhuBejrJ/Rd+j4SJPKoahcOAUsMWmybhl9UkR
s4QXRc3I3FOHX6UAQ5FDhFtf4XNIHuAPfP6qzILpz9aOFgAUZTIPbRhFmVUq5tIe3l/UWLII0X8Z
PSLli/eLy7hBfoG7kTm5YFfQBaPJffDQHu+O5DtWUA46RlUORZKjR4UcayCUxuUPHmurUdAORHC2
nv54cbqqDb0Q+x208HYYZ886pLFthcAVhavOQxls0zWcDH05Jj1Yrqw/lf/N4/KJtQWZghZyEIyv
d2qUC8joPyOjJxVH70yDgQq68PzNP93IVyZH9Rd/ElXKwJISBTlM02XPTjRLjD5dfSQvNOT81KAn
ns1YrGKFj8XhETFRQY/RcwnhTVzWFNgltZ5gMSijltKrdLWApNx7IIWnMwzRX2mSuPbz7EaQ0In8
s61td5J2uwGFoR8OCV2S31OIyDpRDXNxdOuLOP88wJzm5xmCei9vfUIBRNP/cs7agYERxO+f9kHu
tcOVc3CXjzS51EbsAzlt9c6cJzwtaNtUrH8LjpgGzhk+FnFhYoYZIuwjdP3mHfjKRT4341r8IL2e
vFiKD4eBbx/QXPv/chk2xk8x8YrIWhZn7Fg70eoDeiVbyIhKHZjrsnOX+5V76i6IQC9IKY5QLWAZ
/4oevrZtjwMO1IZzCXAiKsphCkDGZ4MU5NKFvIbXNIH/3ysZ3mhSS2rEcRSEOeIDCg/B+IpOE9f2
KO0ZDtOfcC8lx2SFDDkTve8fs9a0ekXW9dzJnplRSo1JSEwz9qOFrOFvsM19nbRA+0z/Dijw/dla
4hqjRDLsUzT8F/wXjzM0C8ahpHP2eN0A2tNbHHG0rwun6cdaY0mxvK620BQoEJ83ltq7eBxkssc4
JQKuEI/Ueu0rjVGsgqg5PgEbS4euRw+7SLKOCu/3fTLvj6MT+GBcXUzJ84dYiNe2oNsEKB8ctzcv
yhKFj4owhceLszpWJPBI1W23a5IvrYSMdCHwzroszmxRerXn3jiyeFDvYS9s4W4FAYYluHWFfLW5
0og8We8T9wkg2hv999ykuza8hqMaym7Sp/1C9Y98Ex75VWvfykBMouMcEuYxbfDkcjjAmyXMqnOk
2agJLHvhhq81XQztThuockfDvHz1GQFGEj3DTKlW4D4NER4toEbXChwaFnlA9gVdX0+2uB/Ze49F
nAV+yxhRK8dVwohzm6sblild1JMie+3s84UDKFGo0BGdygVnmEWJqcR2bWBF3T/3H35I6YzgmShC
z5RsJtkHV9GtzgspnljIpJURxmUfaCvKOGJ+Tk2Z/BqT8D8BlMQ1XpYrsGcm/hwM0B8l1uRbXFBc
QTwJIdBWuM6dN71P4Xtb7PWX5f6Ki+/tezxIS4ZkoDYcB39S4pJs+ORv8zxnDsTIvxum5HzIHmMx
FWo+qgaUr3sjvtAm5Gg1BGfzlYxOg8Mh0nhch7XaII4qfUepG59TErvM/S+Rup9Rq6ILpu5nOaaq
Q41OCmsQ/FF0qOwM6LfXQ3Lfk+0aJGtA8ZWHF56Cb9iwkleQefGJNlM4cXPSDBRu3CBBslddsfWs
DY5+PLKwQnVbs6asjjcpdbHGQTQT9IxCHhQLRcBG6r06OL2ClnQ0yxGx50wKLraki6kU1bUBtrLG
179cjLfqhkB+MmOEMvjWzKoVZ8IUwbSXqHJtIraxEW3MiMY2NGbApvXLtJtI0GPwrhxY8Dng7lj+
U7CMcL2jMMwskLm6JWvXDs2JkxKrDoXQISYwx4xmSAlGdlKBKxKu9jk75wUb1mv5hw8TuFl7xc65
5G13aJ/wgqAtHOEi41tatfA1LRhyo29dSIs74evDQeTJkRBbn3NZWTicOcm9P2k0+dJ/UNwc668n
uXFi+wVal7XGXCdQzKz/v1lzuJQKyQ+Rk6b3cPKvwV4w0/3yGIUmG8NG+m8GN1cmMI8l5lrWcLRf
tGjnqKgstWbxt4BzDfGkOaI1PWeEiShYrPrgNhVFtinaXlVhfvXDpBI009uKPJwTGEtOS2uCYKkZ
0KScsRRooyyHfDpNrKuWjSruNzv7fMzsSp7RGsbTSspRu8yCCdsHqPObXmFU7cu6PlmqlnAt9gmc
AA5PUuXg1LH6k91OfykX5me8Fpxc2SXpWoCD+mQmR6WqOV35snYQna8e6bHtOiNgQcQY/DVtzLOq
REwP7ioX+FvfBpkOoR56gd0R4II/KtpT6J8lobpBWuSN7UKBzdYO8TrvkWyLid/km2aUDe8u+ZVF
4ZQkVdb01FdxsF5LYBuUGN+261w+rWV0k9lQEqvgimGAv8Gqq11R5bhJYla3ZLBDtYZM4VMGqdsF
aZP1qqBq8Obz+XV5KoFqx2b0rgHoeyHSqzSTTcUJKtr4iSsYBnvSdVjzp/P9DGve435g21GMjPF1
9oo2aZkqQ0PNJn6j0dkQBxABUAmSaZGObyXcnsND/JEa1ENhHNNEtJ09pGGTwNCPy3cWiaIy3QM1
WzmDhGyVcJnnovxc1i3Jnv/B+csP077xwSplUEkhmD0uSIjm/+54KNCdOoctisPizNnOsFyemGT4
wROX+asEkAgTpG301I334SUW+EZPtb09x8cQ8LVRwwWN5JXYeKjLmedbfVN+IwwSy9gaMszlOmOe
nnwsl9PlNyqJnX0j8/w0oTZyLkj9ubqVx8CgfAwOpJLO9BFjShB2qlTFLLmc9TEDNkTAwHxCQOB/
G63wVBE9jpwhv6sMvBy0c3liIO8HMVt+X9W7pqe/CHnmMWBsOP9gfGSNp+jVw2nBQFlEalzX8gYm
+qq4MCVJjYDqvGJDMKtHx2Wza24X1Yg6ltr2bvO586jchmeHyKAqFFsHHlZueuB6NSO/RoK6IG0O
WExIin5XvUD8tADkYW5MQcAZOSDN/PH4VsHn2dmasXUVwwwZa+f1GCTgEjJnV5Y7TsjlOYXFqGI9
qYEzP01ddx/QD4PnvWbi9vZ4s/1waMmiZ66jNx/tS3HXKL5cty8/BbfeKHLD6IhY55DqqIZBHSla
4tfxo2IAtZtJNIvIo6Q/KSXCjv6q2mGm064wSU6syec/AhR7eBTkh4YPyecoQMsjxaNIiZT3Lyrm
/PlT490zmDAzIgn6Mde2YB2kgGsBGCMlmIMCVEAxVbbwlxnNKGN6IpCbnNhK1mfPM0w5+315m1QQ
dzLndElND64tmbs26RcL9wAQaTYhUFPdDuXVanK7rsQNOdlDCAjjr4YbG/FsJpk8fByli/fAkOfO
pqJBBpky7FXV3SXuiDFxzUhRNCHVXEZaoMqQx8enbKsg0pIxFR/J+XpCbucZRDRKp+yuXZemeAth
FAmnjnrjpWguQ/H5iFIPF+1AtlxL7eV81O0bvqyyMwKi92u0d3E95fZk7C4338x/ATCk91cHccZu
uy71ycEaD+ZdkbDSBiJ//vYrVIdUorONmemePkB6pCR/UeTL8TqDj08ODpeZZEypAldudskaQfYX
jQHBA+48KQ9JjODDNOVtNI6590uJpOSD9eR2YOzfm4H0E0QBzjrTDE3AdrPgfDEcmJjS8XPTJM98
ePHsr8OWegSrUbGMR8OHLVFVmiA0AFA0ArL9Ek6uGX+QREd6X7pwgHejYUcrG/NtDJTfSZutgtPj
VZv0089VI5A9EXVOYF5mSBW/EYvs0XcwlkthC90kJv/Ol5gk70DEYetey3UV68iPNidp1+D5zFf0
yyJfixFASaW83GAQ6pKGll1JyJejfX5h638LnTl0c3VCHn6ypvS/Sl3NgKGjjYRCFXASwXSFK1b/
g7uFZrsl/6/rCGYnV+KGc8/avP76EFcfW+KGjmfLDmVr5cnVG21Epv9DhQ/IaQ5s2uZsbRYYip/K
2rh+olYuEPzk0FSNYI5MQIGlSrD8ZPOLRfPCpePRJ/EKSioWTDxcsTU5YrqTmelQhaPJ3DRKoRoq
hp7z9k9n+/m01TpYwtMO6F/LvtCSBQndv0ySSRyMBXWlDU36f/DPFbdQJVAsdtUO9sljiF//zKen
9z6XR/0CxT6RZ4utLX6WSDTvc+ULDLC0bD7WSUQie2q3TGGIzM52xNAPuIYY8clhoOnNmlXZxXVN
NvtcSKpAEvqugM/WKQPbs8B/0jRFCY+f1wmwFI7OOsoxbk/9se5RDhv40fpy/M68c7MgzEsamFDd
KGQ7wonMqF5rOvEP1dh/LDDc3Waq+34S0qluPsdlsphjodbE3U9Va3GOcuwNm4TO8Qb0gauGix1h
I9qkuNEcpUDABUXoOdiSZJJZdirui/xCRK/AhNUR5McUoE5d1xp5dQyaMEP1Va6J0jsGFk1ajnao
O3fdc4yS+wTVbYXjIN2OnzMn9dWgRbPkEfosi3buOSv7Ky3wW/xhhNBfji/LQyH+F+dPRTnqODTb
ppZsNdnNiVxalqv0dn8Y2DPKUsHQrKEd9RdcXf4ZtEVcO7GmlNeH+GAgDU/Sjgsrw+9/VFvWi1uW
DBM/eoiYkYtUPGxSHSwj0Oxit25EdLHpOmgSoRUqIOyS3RxYZpyMmurVb2jsc+FvQ3WLB1R46PD6
ZuYaynsQZO4u7lYgVzYHQPWC/QaU12XUacMZHZmMLBygrImBilC6yZozjIZ+sYaQX5+ZMQsqSboh
xMT67Vku9powxGpHm3MC194tEghH5xwChAaeCKOI1bbagzKhMzbloC2+DLHRekIpPLpZME40GLye
MHT54PdmezasJy2vIt/i0tioc75vTJcDwXMkSecxw/ouPF0Ir1XyQqZHDV8wMEauwu3fR4V1hmh3
XS37xse7rbAj791ILKJTsj23We6bUjU6GOcfeB9k679iVY/X/nnlRjEsuVPKpIrpNc8I9/JrrvsB
TGrVb698dktWq3TVm3uc3w9bcypYiSgvtefdWTm1pFIeBI+wVNnCrWVi2u1+L4U1VoE+eqkwTQKD
uyurHJYZGic6G/yRNyptDCOAKpqEBJ7IWa8wBT7G1ZstzMXOgjRuzfcrxgX5lgmNO9k6vqgbVMzM
AVJ034mGVk7KAMDFSuYec3HvrWncTAQAIF5PP5AoouyC0QbnFY44C8HU3sS4jzaL8ybzF4zrbssq
PGonD9NPjxkxnVy6K59K7bADRwyX/0/wpuoW2FRHtEDT3VqK66RHPFdKPvuIcZvsqUqPGB6619v4
MxANoysMwc2FKH6B12UIGCviRnDxxhcS6BdMFwVqFjiuqQ4Q09f3NlmFm/jPIGWGh/TMveIS1/Px
ipEt1apQGlMbaO+zk2X9k6DyxjpAuO9SYFp4q78KAq3yxKz/wb4fCJxCDJvM+trS3LBh4hy/AjR1
VuYPcQEa2ea9xbZ89sIHQ40L6DZJXd0MthW+JZwm3B0ogAzVYUZoCMUjrvDt2UdJsMbJIwRc6+dZ
uvF+u83pLkcMjQxd/sfd09gc+ew0kMQiLU6MbVU7H1oy7UEhZVBd9SSZpirgepcBgzKvW3z0223a
2/JUJ/CbQPWBBRaXZx7KEk+KRVDs7CuGFcFnN7erEdlAnf9DR7az78NVW6HB0tWkDodaxOudcoYg
2eO8xefA32ZptCqBXnt1nd+dKi9pmj4Hwwrim8vqCPzZolGjd9ksWytyWNuhlb5kV4UnD/qT9gZv
aVmcRb+OfbEcvIRFk3Uo5x0cNdulwDBs3PT0lfXG2aRycgL97mQh/Jfkpwzrt2FKOi4v9f+vpemF
Jj70uGzCBn1j6wEwkjwm0w4MKd+gjhwqtTOYluqdYsUdYDWlad7Fr5aAQjV6n5px2ieHB7XwTdZd
7maRnETqz7aWXliy9bqzFiJQxU05eByWPKLE6vH4rKLtd/u2trUKLdYgv5ubyJHUcGTER9pBHKbm
YpAsWJHB/Y69djAxaOwD/upypuafU+LE8qVKf0DZWDkobgX4HyRLh/8daziQrClmmo9IIfjs4Fi4
F7JPKSEDaNGulJ70iab+EePYr2NKbIjoNG/rLV7Y4GnIPeg2fJMQ5ZDI0gnhRSK4tk3u+Gptu/zQ
GjNNL8jpZOP5vCAfGkS70LHllvwfZkCA4a+1l+BE0mz3LGrKtPIqAcOg7BgPYhBGWCzI/DrtnEUf
q0qkm4QHs7Y7Gw/0XoU7M4w8NXhy4rWeTuC9HlWs3LvwHZfVZ6cBz7rPNn3tINWbhrbWks6q8alo
l7n5TYraGK7Te7Xo8xA0nCCem0GQs54/FRhCNBWi1CYWIMEhOiTswYijLm9ynDDlvc0PZdGxCnx7
MQa5bN3S1gZedZfe2GV1Fj9G+XDGaOX0B6HPqMce6AZwMgDSTgERcKwN3cz2twdcG4Fmq7Tr+QAG
t5JLRVjg//ySEvEWTvvKNB3+bXhPARprlEQtlqXYKy5BSZfdi82LjQvzI7z+gUnuF5k/j3UxyCtt
ILTRfKBzHYBWsb1OOolNSm1U3qGlkdiFn9AkNSt/iu369XN5sOYhCET+zoy8f1LXpQbVfucCQiKw
Tf5pYVrnKiHa+qe2YXwgfZAu6PB3Kkn6fXcxlvXP8ANRT+Cs+xnzxHTBiFWJaELWEBlz/eg69669
Gr5AHmq0R96axOGfHDLLYXGe/Qqc34+sehVhVBYrZZowt1kg/s1DSOS/mtCcLXXI/0XrpyGnb4DK
jHbDUZ0A4fmh3ioi3sW75hUEfjy4T+jODxTElYR9EPbi3BsYY8RNQi214EeNkKsAB/5mH++fdJG7
t+kcutiOJcUsA3mpbykCLapbu5H/h9rOCbiTQIU8lYdFX2Z92RMPLTP8Y8wOJFmvAnPW4rIRAb0G
R2Tooz+QngjQWXXBT+wQkHSuSCnrnuzIKecXaJVWMX0xZeRlA7iTR7RSWR+JAg11LKbNMyxSq2YA
kexPeI0/yQrWtZTwRlG2AWzQMKK5Vay3vhM46glP9JW0fsvHPGr/rzD1L8EJqxu0rugUZRrJiIa1
efz8TrcQrmOLxJnTTyr0emGlOyIoablcakWSnhpJbL2slYk9mCHLxP+8RHO8u5WX3tmbQjCjR7jo
TNi2XhaouwCwKjtVkKrXCLh9XsonsbEoVMTHBIGozDhBryMQmQ6gp9Xf/aKkzDGOyID7aiotiVOG
EtIrhi/WWrjkcmrCGwXLShyaIVhUnKprlLYiZ6WY/yi6ls8EglPsT5lgbYGHXV2tmNIvUREDPGuZ
EWfc1KG36dNGMD+oPjcTLVQnoxerQlDK8X/oeOj9o9XNmJC5stYqD3oUaJVk9piXm1DbfNvDP68R
TzItT5r+uNahAI9x0olJqOUL1U8yI2IvUvKfB4kTbBiD+NSquGFaFrsZvdM67VMcRBj+TB9uLEN7
1y/KfQu36rcT+o+CZxq2CNt1Nywjxv5VIIqiSwFb9xjIKZgvW6T1UIO4QJy7s/i22FU2ze0HgBXI
uuUeSMT7G79Z/kZEZTI6eScUuTUFej+JQ9WjyOZ7OfmzODpPVocaTBn+Q/0peXq4xMmg076gA/3z
7PAlW+8Ov/eJda0y7r6BND4ejEJr8kc2ye2ZaLBQNUdmk/mNHNrkX5y1CU+V1cs9s+b2ZkoEmhmq
fKWf1mDM0JKcfMedUxDsu6+q3kGg6lJbt9OFA2cj+4so+OP60Z45JEcCFSu+jgUHa6daltXv/jUq
IhgsePmamSNokRpvlvA6dK6oPxJrrRx9Z1lG2MnND2PUMGbDXyEe5nZxvN2BIllA0qsG+v9KseaR
Fni424U50dpJbU5NV5EA4I0OvfAehRhPVgsFnPfs/gRluncfgYU+4x7BN1i5ghPbxh5bvMD3hs75
x7qTgBzZUZSu223ZLSQjj8txxK9USCAQ31Gj8pi3+pFV7LMAiIgzakIxX/9Q+oiOnc/wkBwIKcoe
C/pygFK7MUP321eay7KwNSwjvaYEO8d8lpWKTZaiOml66N+OxyW4aGfGg0ZedlaAM/HjaIc4deAP
6bbSH/3kcAtbfTPNmDniWdca3qZAsVVbSwXoogwL5aPghCB8tpQ9v+BmtY6Op9TrnZwfv+mX6bkG
0KSzLsJAjavFYFGRI6tHdWFBUaI/1z+84jlaD+mDpXEjjUaQGE2AFgOXdXVJb45N3XGaI/tui5Jq
FlF3Jid00UCzqe43uV5zy90ad2mW/TRD7tMlrQkIKw9WH0/Urfs3nYhGNau4N+3gJDun1PtyfH+O
SvsnomvTcDjN5nZCaRH9sgJzLyCtjs8vkvZmbvQeMhoUdNm7IDdMsqfugcu1co4CMefjwt6+u8/i
LwE2D2O1BOgYI1WtTWTnlvR/kmiaZMxFX6zBY9m23S78eLBFwAn2akqqhFsDrZsnFR+ibz6Ub82e
I/0AP/K+5AIFLq/cMSCBbPZbpGhjJFUxT2Ur21GM5z2EWjgQSI/4G1MX3GF8kiLY70a0fuFZDODH
qMiV/lXUiENqzf1UbeTMAMwYA3ucE71rCjHJBGNGLPBpStUzJodIJwQJAtWr4s79K3h876fQyB7s
MVOjDgdW/Fv+00eTVyhWL13dA+gJckUQgkiutZVvlwOM0S76wZO2yUr5Y87V28VpbspN8W9S64as
68Y4lrYD15OkhJpVV4asWqnpEglHDn6ppIG8ziN8Wt8FhwvqyFr9CkaaFSYQOU8/23dyfWh5RKww
BL4Nb/znJOIO92HFSEB3npmu5qXeA0+nA/13bBlmjzcerNi/k3LrPkE7+ozEzef6Wm8f5PRlAO1p
5gv/yQc4+d4QWle/zcgTMt9M5LJPvyxVx/bdVelZmZO+4jWDOsEPSe3llM7iF6q4HazdrYP6sSbu
qPphHxxjlTZSCVuE6JPLpVkJwRFuGw//UC/v82o0zOFzBZh3UtwEXoFferZalVfBTK2LOgBzwX7G
cKrKeUGUnS8C5y+quVVejm5oVsdEbo+38raSZdTBqBZeZC6NqU/8RO0ZdvmQjxdxw43sN5JljgxY
zPqEKsDP9Hndz6P/cBFGIFx1BFQozamoIzxYy5pzZHdFOnbKZhnz6Sf96Hncg1DZ5u6e8S+LZExo
N8DrTUoj81dW0UmKTOrN2L7/A1Sxo7He1j8Wr0zZKZU6Py212GoTnclmIj0+MRSkMD0HBvJ6UVEQ
aRHdg2YwINyBRwT6sGp4d/BD4C6ZOBdW4jbrcZqcZi6BhKj32O2shKxyxr5p/aHFENzZHE+pprH5
euyt74RFbwyJCYE57q2BU2dS0QSbbLq62f/dLTZQFY+T3lU7YLga3WlwKtDGRoZjIS+iubEdihAv
JSfzzputahkmoFxWmJRKsae0bpew61X1czHq2IOikDqQspkA4kHLkY+SQxzO72ZW9tOgHLjtFWKZ
hCz43UezL8xA8sNaJH7Gm7BSGNs5dSAWyXvfazV4q9v0WGxLRlCWmHlgySb79to49io0lfdhSYx4
yryfJT/I1IAHjBhI3s7bwzGuEnVDvqFsjImGS9/YuoZKS0SejZCgUACU4HWXa1SiBlr5VWG+CSXx
A9xeicYT1tG9dc0JltPTgaGEOZcQvqwDqX14xs81HvQG1gSAYnh650AgwxlIX40U33bpIdR+0aQc
iPclcJSja6L+E+PGcHGlSsg9HRDuV54M+yjDL9+VS3z3UkHDYTuztBd2fvSnK++GFDPiwJyP/Utf
sr0TZCLNdiC8a5w3SWhfYymdETBYUhGPhISo9KvMMK37XsL420ublBF7NTnWeyADl+RY0Vu4SS+U
Q9nvuKTtqspgjl1snsISub67xT1ltKcpJqRAJpDXdwvfE5MNzOHrYMi9NmxL+JKIIpCmmAbnkkwX
ffSOvkEGsFMlDzyW2mdntE3EpRh5G5Lc70WuycjHoIUaVM2EDxQ2GAgZZVTxjkPNAUxgm3jBWgqX
rrjKhVtq+X71KzFjpnh2WAOPsJ6cx2qnEhfdXULpEcRznjbE1XrvzOnDWjvgkuVieABwZ4khCvD7
vZcKa0JUOEFGgKocASnB1+xkTzP7nkhHZEff5j1kazcX60bJ0ttTTBr+/NMZflWkDRImwmGgLcQP
oPRP6x/w9cXzYMm0V++4G1csGClpybJNKutxklRTNiDd+wuZ3Z36Mt658KCHLV+iMxerohdRPLQO
X2LvjRpaO2z8oGU0PIov+gFkcCGMOF2OKOdkTSKbnMDZp0UyMRYJzJlBn9KfeSn+pNCFiKZKaIb9
Ix6yir1oGTl9IzP68C5RGezMvkYsaDzgHEzTLX/EH5dn7TW4B0KwYsUq3yCgkAfuFty9x/KwFv13
/kWG0zjxb9TrPVZPXze9gm4OAN6fc0Gky3NHTifE7rKnpNQLy543nbFBaWZugYSPPqAYqSRXdmyg
C4W+A1gY/JI51dc1h6cOWKrTPKX1Lter8ZV4uHpBmTaK4d9wQxp61iwdYH90RB/iamT94imbfToC
+ZDdReSi3auyTUcoZVd7IEe1qSGAWcp4FJo54mamJbrKw6IZ2Ym7x3B3QORt+sFgLRNDY3scEx0p
l0yolCXcLZuaGZI8B74eIz75AXJfVHrKAifWnR5XuBkFo0+Sa9ehI40ZeoyqessXleSOOUiHa73s
Pcm6QRuX9JQvhL0GWdU++SvcK3mxuHoRIdII0jQKMRJioyNSYAc4B9ehlucYbvDEhrQzWpYnZkg1
fPin97Ta6PEDCpXiton3ZOo6CFX8TLDlADA0Gmsnv9HtIZ9+ijZVdzMwJR4/T519MRkFYdvsZbVK
yBTiXF8t6xxz512XqzDO7uJmBAgYB1F3vw1ghcV7qaPSky8B2fa9++1UF9orXGXxQ1cc83/+ZbTY
Fq3eYCI8SvIR3mZ/f2Kvyk+TcXQugsRCpfEe2GeVvfiAjkwZfZl1JWpcB1oFSgwUUG6Obfi+H5oT
nak6rPIf8xTB8sfqWvBW/23SmtO6wKoyxqGmDEpw2ofMztHyWOBqrWlaAl0CWNcFQo5L4JZjlpbB
dDneHvGGmfS8t9EX+l0Cgyua1ttiD6s4dye7EBGB8uk4DGew64g9b0FtEAVx3dM3itM+kZOsMkhG
oWaO+p3iL3Ngwe5b7Wjjw1yLQ/XFbEpdeAagCd5uecJP23MlKf4l84B9KgKn8rivyH8rtHMXhIXF
BgbDSX7wr0yEEmVhxout7GXjvnqu8lDdoqiNly/JAk2dtQYVr5Rc2tkdmTO87qBsyxyZB3KzBL9A
ccI+ASDfFAjTRFFfjnio0mt8k/lgxQQbQ3CY1eigiyR8gMZCdaDyh9M0u7I/bBJ6nGBv/ws2neJD
bufceg/qF9VkfiiWEQ89cvX7ndBkX9JsdCbLP/wdW69cUSkP+ciDSddeB/MSV9AHA75mCZn68Z7L
gA1+5eisbIN8cFLJeq6xhAYUnBnIWJI/0NgWeNUFlx6ziFTT7mGhMfup4dcpg59VgU0MRCUKLtoI
pu+o61GhJ8nlAIukVkdPdffF3EfwcvTjP9ya5qz9SxDj8pPYy/U+T2aAD9Y5cqVlUg2ZOyvFKF5s
fdfXFJ9AOFxyXT4K0hwESBkKRw7s7wsJs2QhUSXa5VXpw96tXhrJCeNO3Xl3lAgmuFCriziNcmsV
shlEl8uXP4K24k0c7P0MmHOGVYcKSULroUQKbYiwZL5MqnpCnUCl82zpYPYIOVjVvHhKqJ3xkqHx
sTreUtq7pIN03hBnsynYWEjtiEjfVte1KBZt9XEptsAkm/FjPlBXst+nzK2Y+sAQ9c3eDY4Rgw+S
v9ZsjC81f6e73bY3JBLRKtaCVGCCW28Mu1lhw1RJqDavy7wipohq8wlQYUnTt347B4JS9kwFCJJ4
13DReyskv83k5tnDmcgsAh9Z2udEgA5d5iiKEVtIBfmMHkZKPyfaVwt2nuOUqIw6v4FcN+MYP2xj
xS4jSRYxcpcZiwNfrbGSOFRLyYbcvIXvi1eGXcBQV/EewX5z39qMf9Ob6NJWHa+MDKfBJwz4epd+
FJhUy1cZLEZEBpB35UbfIGWAaziKomeAX5dmzFiw5FNcG0pzKMVuR4N9JIe6Me1D3pUmPe81+A6G
uWEhkgEZlyO3JLDmso108IkdIdpWvU2Qu+YIHqIOz2vYnMBiorNMAJw/6re7h30liD2q7WDbU++t
sBO26Ty5vblE1zjU6nBoeU5PeEq1CNXQCJHxVJ7S9QGHwrBs0tS315+9TssrkZaOyrfRgYKtyHnN
kRPJE+RoIMUdy55KEThF6fdW99Z9cnfZQS0pHiGR58CWHXupGIGXSt6v32YPO3VHkya0q6RqDi58
9rcVIVWSrWNFOCcQvuC1hvciEmSmsd4Z4kIAMKRDa04Oq5Db4DOrk+Hpj6yTohz+oGfRbF1DFeR5
HKVw4q3ZzYbJK2tO5CKG1VkSTmLpXy/TLxE5yIGCmdHZPt0pv87aR8thRkOiesjK4UtW8Qig824T
Mc6+fGgYNbSbWU5XSDkqTXZRwTr+RTHTnu4hFH2So3Rc9CWDRu+qIbw+K3SVC8YrYhMjx3dWdCD3
3JIx8Q+SqGN9OieThI0ymuUgl2jSaXZl9fCcIEFIiNqOxLoHEQr5HDFrlALFx4YrcnPAb+CQvS0P
YVBpTbxcpQoyaH2P2xXY8jC0JUXma2kg5j3wWKgcUQBA74sWvZqOr5/OINxR1jkDd86mnfj8l2oN
EQyTI9jyqCnLe3R45ex83Ry4quRWEUnuwkQf1Ku1cS4dU9k9J2AJDZud5h0GKYrN+uF9R4vyij9G
QlM8SnQObHt3rLrWwCQ3XRAsJMegJ+vUvdTDBYwOq9GoDN37qbOW2ihOYYk6+kE++ZkcZv7QF2L7
9QFx7MoSKckVHV7dXVKXTZfT7B9euWqSQ0BDXxlfGf3slJnDDiLpPivD+23MKNQfeDS+WqTNCmzg
V2eg6Vi7q8/W9IkTwkKEJeXKUlL+JLxif82Dgi/ACRDZ8bply4UheKbIebiTuD7G3rYCbnocWC3s
lI+91Ls64qDc5PO16Sh7bOUTFMPpwjMrYh6MxbFwbd9gzKo24rQQuc25Uzk9S1FHNk90WnISCy8L
AH9LiVEvNsQT09I5wlS0H4LCuW7UU354an8vasnyfltpCoq8OvYseMKFSn50IfTMkEVnatDvLGjQ
z97m6JEitZUc9yKnnYk9/JTa4BXWL5O1BXdvqOwxJgp6ludpnpHpWmFsGCJr1H0ck072wJ+BwvmG
o6gkXYovQzXKyk+8JbHEjAsAvszxd/DrA1M2kcXXUUcK4dy6sHluXrNMfCK7wb+sXKko0EsdqdAP
xiiLNmdk1qAKe7cH79fsavZxP9Ot2s+AvaEGYygpb1rIJX4glkNqUBeFyzVOqTW1EnNn0F69QjQ0
9uh+dKPMxguY0G16i7SSP7fqZdnjw9nCPXCC+24GVdZTCkCkHbcZjsjk0Y4YQfernUetkv+1pwfr
FE9YVuxubgW7iZyTCTlsPZbSgsJ3KO5iDl2FxMC9b/LmR2xNPczV9t5DXTaKMOs9NcGPxgw+5QQt
ekFjIGGP8V5SA7TZW5NSi9ahUXHG9f5gqmKRWqSyFviIKJkjzOIwP0+0/jxySo67tSp3lbS4Cw5B
ySpHk8woLdnEyaOn2FqndUzTe3Ciy3ZVPPgfV+DWYZgjN9JM15Rq7w0CzLba9RUhLp/IVbnGu08z
PGO0rhsl7AonqPB77BTpto6J/ZsF0Nu5Vwa9LIP9J5eR4JYNdbtMnXsJEMa6+NfGCNcDqSkuvZf0
HAE605ZPPJNQ45KqcMawryTbo7qTAP9bp424tU0+A0vQ/DVKoMxGSo9rqFkasof5ep1ZTAkzPfFu
AL/w3UdBwKaWB9oGEpnMbnM0oXo97b0DZICibCXswyWUcT8rJJpYD0CyVoHxrta8G0V92SQ7TncE
U/YWWl3itEbxbyQc3yDZ/r1TLqxOKdHzeQpVgwiyE+5ma1byvZ91cWVvV7VLWx/rp/J3Zs01kqU6
lBG7Gvfsu04oBfiGFaxb15jKw2cCYc1a4PdeeUrSRN+ytpq9wUxtJcw0vT85Iadx/BbPTlPkwchL
zx6uArLesbwMZPmrg7XrYhA0DHbiu0Ja5nFc/CnR+4sm5+PE0nfqfipZFiCKzE3pppjEIWLeO+FY
T/fnTyTHw1z4rZ9+heV1RY8eKhyLXQ+p8/DUyCaFzM1AHjJkoZ3f5LHKI84M+NF06p1fmkN3eUam
Yu2/FYzAzoAQA+ARMvhhd+R0S4BqoYY7dAx6VCSx9oYX0Taan8r4R+icl30R6A8+X/seUpn+BE+E
MXlspwCMudX5vRyMFEwIF1/7PL9KXYTIqwxK9V6lEctCT5ZPYX1kI5Cl4vF2yUvwiVZ0K5ZFf0rT
kzp3WO3Wb5HhQxVue+LB1p7G17BK3pZAdLp2MYac+pNpRQ0CwSdv7jvdK8fXZFDkApnoHwSQSCOc
5L033Y6G2y3NVyHT2qjswZqnBXifIk6+IisCX/E1Ng9WmjTbFt5G/JqiHUGT2DiGDJ57tKAAE1jL
DF8rUX1IkUnM8mvc+Eb2Y3KOplCX8mtDE37Uqra4YkxWXKezTpNEYJ3nYWJxVLJ106SVe5Ne1aHL
DtS0daSdcVN5tCQ7QuudC4ocvIXMvK4kMLA8Ql/kGpmPs23J5Q272/LUnhUzSaNjekAwbdB6aEvg
g7j2f6iBMc95IfzsnIh7z1bw+tyVtVH1AVh96d3wCe14jvtbV9YrY+o3J7WUR7STu2XHHs6Yqewr
oTpXU7+tdiFAoA4JgbFBt8GKMl+OF9IBLGHx+FGPzvgZDUaZMJ4Qf8SeFycoT/nijEU1gtWCwq75
Xld9AnSiy6W9DhC1GaLck+E45Kj6GtuwTtrSbRL5p3sffTdKK9t7glLZG1rlsk4D/WscOZPizVFO
GSzI8MrcIv5u7t/+OnokiiWXNvTpBlcJZWbx/8xH7kAShfxeNXbPn7Fe9tEhvm/tRkg6qtlArhKy
5ZXyO9xcAbMjMSEhfjK/C/srOfFyxatFyl6BjeMRyJsoI8unUiLlvBJWdE60RqT5WrJDPTld50uA
+ftXAUZLFCSbFnWOPFdY6hGCRcYyNumeNlqoeDVsr6kNQL2tZuHUGqJupTXappM5EoVcRQ4cxsUw
kFVPn3Yp0vpJ4Sci05azILj9iKbNSMUaTiwQfhcaMQoIXW0jM3rMNdOXD0JkoQOccSgZvsPs+UEV
7X1hhV1wIj9Fpzd01ZJzrMLdRjmA8Sd38EXVsb/HOj9sckXP/l4LNj8z56Jm4qLFGX9ZPIhUm/or
t2Kvt5wcpGpDr57UMJNrB0Nfy6H1Qmvc8LsWOSdxeIPUujD6fSwDB1cZB/FdAlktm0POB/ZX+T3C
MDrkuQ1HkvFmfADiZH6v5hWIbhmCDMFGy3xQp/QFFUPDa6FL7x/r/HuYZa98ylbpChayy/Py46dn
6JaOSyt7IQTKRudhXjEloaWH4GOnaWvA2mLBBk9N8UuoE1/9X/LZ+e3650mrGOVeNjMY7VEedIsS
BgFTfD9Ep0woLBj6TgeIFzuuo6dlnA4NF/fsNo0fABeIWtZNL9rgHviApAP3zS3jBmvPxhtHnaxw
VdgCSMTPhiT4sT9RIc2sz1c2Tu3iii8Uk4TtPLN4HZjk/XGkbltfPpohPrb3AQwOpf2K723Kf6cD
RW0wF4/9yw1R9s4s1i4HrhhxBnwioT+oZG6SsWMCzqb7JgZWkxYhXECVzth621FrE5rPjHoXiVyW
sTUvj3SlrK+9yxUoMuPEE9EQGGgWP/FozQoks87/ZoOmyavr0YHKmAb49/7alv4kSM7MTGncB+iD
pIa8I+Gcxbb3BzxT2SqjExwhRgZArpsuAaR8ws5YKKW+TI6YFYzaTIUihbZu247mBDNOgDX77Eee
bZ2PTIdr8PvHb4K5XdMJQnnWxxcFUvHUQ0KodWU16BdD0XntDN93kkYVanMNLROfY2SkAvLqB0O+
RBvCMuR4r1vi8CPDlQH+sTPIs23hN98B67Vae87Z6LvgwOgtYiJ0XOoIE0AuL22NpsmTwlGr99HH
Ei6/MUjiO/OpcZKa7BIKRjVOT5IZ1YVkN6WCS2QLP/MpNgt9LJEsRGkkDknKnPLzXPfG1KizBAkL
i1MnHgwhB8prNI+TXYovG+tnLv1CL4r0ELE2EWcM7TtjmPRld6EifCeJCompGlZicZx7swoKaOE7
Ew7+ihuGSjE6L91g6Y7cI+IBNhvC0mrU7dsp2M5ln2f/WFqXZgeHNxH7VPgQOsTa70w6CJif798X
Zxw/KB14mlk6vcprscz3N+nXUKZnECnMejFK3J7Zs1ryWw1NWRUQjRrRYHTPT5Z261PxG94yG8gR
yIOPTW7Q+iN9cTnYgFl0Z8vhL7uCM3glm5QssT+JeW9G1uriuhmwmMmDNYhzATKhrTfIRyQQaxc6
IVQn+avphjVmaVmvhRskZv+MDFf72b4qDDHjvOmsCO4uyzlZnKNTN+bYbVvQ+aU94YnoJY8hN4fK
NrBpEFiNKgWSEnVAtg3InFvcaRISIkX43REftb4vEPE4roXQOf48Se9m6mNoL6mf5BdM/VTAYuPe
a+0uowyAf1/AO0S6A4hkspgVr30wqujWb4Pw3bs5P2isjrY+govdpnl8sOd20CmAYsXGfOirsbbC
EDyObfbxU9VjhImM8ETk6JIZ2C/EFZ2yLuJUHiB94QPQIfSLvQngICLCB2KRBUtLiK/gOJ+Yq8Al
GEjnEVN1vxvUg2Vm32Up5RjFhRYIPwzZrZApt7LXzG/ZT/ZGU+A1MlgrlO7CwLyozaUISMHji40o
nB6CeVMpi2/aymfgqf7ybeWYhDC97xgjV/agu3LrbsRD84PJSl/CdRM6tDRqChDoCvZXbx5xgXjW
D3WmqNhLLbh695EsDCXj0nlGFwiRYQN/XAF1v+GtSb48CnVlDVqTANZR87PXr8gAxDcRMyQ7aYHw
D5zpxORbj76HTsGRkIqOsVmnHQsdw0xhqTYGbOWeUreJ29tUdHqqZ9QRo4lQ0bfyFuV+CYnOuxZB
nfSeoXah9ey82d6omR5c4pSQpZxFORo6TgzNVvVWMynXU2N2ZMdcqc5qUMzvghwwlev0Hl1Cwlo2
lv/Aae9QTqSXnC/3zYQULQbH1oBxQ9qb2xJlDBK8FAVsg1MFe+Ois43K9SMxQhp1Gl09kewshs5o
j5qArqTUO8sRwrQMgHBmhAAUHmRyDFuHio4Q8hmk6lVtqUwbiBhfDC05ZREV0L3Jx3AJffQNZ3dA
2LwM7AteKu/65sRS1vexR1i7J8n0AVNYIoH3XB0fzdaugswRK2YJeH5ldGSDcfM228UwCYpiERh2
RRcjiAlEYmqENCRJFC+UJmH8Zc0DjBcrrtwoQdkO8N6ZLd2XQbi0/GsQwDEt8zIuhC+EvsimYBZP
HVB2sNncAQr4RWy8ewggs0vSK5QRC785MwuDEXYk8QhLw34IxZV36NH0Uc4xtFtVuxFXVJHlWx+p
Lc4Mt0icc3eMs2CU5NGqi8YF8tPz04UcEelW2rOKmrARqOR8eLpJYzhZyCdI+1NUV450bFKZhLMe
Uv0imcMQQonR8I8r1OmmuAPeFm48Umh1WZfvXIFw+BaeBM6esfLT9QDxnySsnnbM5XLSAvRNzO0/
Z75obLh0g3OVR7ORzU9cLjCTCyDcPeil1yvQtnbpoaEByq+O6spGHePjhQvTY/nsVrX0GC/rghjS
slow9PnS8aaoMCukb9WVoLBHMVDZusESOLkUgcAhtyT+9Yl63XydDT9erNiyqsC4AXf/asP41Not
EVCdS5xQJHLE2kztLOXgwihlXldqT9meWaCABLcFx0KKtUtQ84XzNNITuoChIT6unIWnMymiCLYO
XqRvBItJjWzrLisL4GvA1C9UcpNLDNE2MlHpzvpHJHS6E5VLmEng8ZKcscB0KNiSrZVyJ/WcPVGb
MKWgjFIjPtp5dUW+x3VulFs9+Qse/X22FxAVZcXKmtutuJ5WZLEW2wuwfgjkrqJiiZgQ0zF/EEOu
Jk0L01Q1F7WmMnWerDiLgVwGa/IMVZTmjxIcG8ZFfpkhS3GXTvsT2umMV89fGNadN1y2AykAoPMK
ENr7YiXx8S3C5nZbEuS3NyUJ7xCCRa4lxOtC5NRge4VQbtAmbM1T1FaYAIt5YaaI5YVvOKpPqCES
QEBlq0fHLztEVbQ55bjuQ1JuM0nSoU27jVpcA18p7rdjn0Hv+qaFGuVn7Dyl4l26kvmI5rOjfSLZ
7y9fq/tPYZhUSc286iI6zKZBYdAcZSA2TeRgG+h7kg4lFwPn9QtGeaNL2jkgF+/j1rRC83PWGwV9
Ugy4+s5rGnAIRsiqbUqr7PpaZKoJpxfb3WnAkOn26iUvmCaoY/hO0z2OSdt2eIe7uySnPwFGwR5z
1xMmuYG0fJcdpxVlyJehOvMXZrBx+e6suP0U1QWyO75nM7YDIihew67d7GVdfHxhJ3QJ/ceTDQr1
oyRFOTUVxiPuE+0z6jj1FJhDVVBBAysxOj1lT4ecdFsPW0stDgQv8zRGTGVj4pmR66l6P7zDWQ4m
MhygAx7mE1aP5O2Lc2Xfz0dFCjvdCzTfPhGMArxJIfRA2UfLzJFiSTmElxzjeILrH9yYjiaImacy
BupaJNdqP4h86/jMwUThANiFq81IuaUt+ZT33cqXxcH6lbtq8oT9BIm0lWwwyVO12XN/V5gpzzGH
Qgfia9NAjvBgsczq883Y0I2y8E9fNToO0wcuBgUTQ9tr75afTGFB8jBKNfJ/yWBV5yw8Z2esmFC/
Yz2xuhdryjBNEfrjBxOlhWMdGwE29YnHa530ogjL5tfxgv1e6gKgP8q2xJDOb39VRiMCD/RBHqZ+
T9AxFiE9tcn7YI5gyaByNAZociaQqjIA59yNtGziTyqo93gTRmuPMr0qVnYvgfjx07TOHdYiZjy5
jRYN8Oa3U1T0UskN3C6d/rr0n3qL1SSA1ZCksUoJKAHlWntUHSRaptOx9ihDith3YtqoP+EbgR8J
07ADERSOeYBzohlfVXb+f0MPhfULDRiRh+wvwg4ptZS82uMv2QKCzzIMy33gOkm7ZDDWcAYVHSwB
D8D94U7mW9cl9IJ/DT8+ve04Rt675jXsd37Q/myLfstlIHcdgK/OeU4LmPiSjAgEMzY5xwXGxPVN
8IeKZiHVH+5JQPZHTojetYlvAj9+LRfzfwdWsPtVrVVnd55CfwH8c9rv+tgbMGB23UJ1fUhJbG5B
wml54UHUkHzQ/FZnnm04R9KFp3Oj5Hnuth5aBpTTqfmUXgtjj8m65HCiwc9XJubQSTpACsE5e5uP
mRdY9aLDxGnPsDxR6hqwHsXP6Aoq94oVvaoLmLPn2antKy8k0vUXKj1Zz6G3YxSNYBtC/svPQVkW
homnK/hxwc94cvN3DNyfTw5dA24vpTW+K7ZyNC225mqAqiWlzf9VgvZ4a3uOJ0Y6QsItsukpTTLS
WDMWPIVzO3/rg8rmHh1PVXQYY3mHIoBEEf7cLXJrAIvurF8Sxql/U2TCfz7G3SHciw1xlz/f5fdZ
lQL9CciyC8zBngQ+IlQ7v3/FzcQaBxsgOgmPIu1kM3g8FCyQSB+4z39gKPUmCX8c9sO/begHUXJ1
C8yWU+CN6bCEn4SWNfT1Bb8MGdZWB+WZOnfwcTrtlw7wxbq58UF9AQoZm1oIPstetYV3J7WimyjH
HEZ9wYnPgWIX/YEWY5HuvDMuLqdNX87j+fdn3vIAdZts6MtYllBXU2rUfAdZ+0HCl0LthBfqiaji
2QHVOMMqibpDpRbqKglyiALRsAs0fnNzYD5/kekq6Nv++WWnSEtl0yfz4KFFwExckyruXQa9AVer
XYBbZxYdoypBZM4KDOrW0bgoID8rtENnDmwl3fZ7o9z3Dbh1VWXHrV8q4+gQU4v2WU1urGCDFAMy
V3k86K67oPy7KsQQMN2Gx+lj+A09j/PZQsE1n5Ji8WlYoFTuokwr5ignnVKx8iqs3oL0WFqNJxdk
UTz+TcK4wuXTej+31hIsIlM7NkgWz7d9BVWL8ctdeslJKULbml5ogrh94xt7oKGGbQQBRHwWBDUu
HAP3SiCaMwW8hRMuYvfK7UZC7nw8SVWdJP2PpTXAdAf1vZFGNAH3fMPGKQEwQwY/MvyjCwWbzHbz
3j1SKIZeO2kHwGFjmeyyalxdx2llgkYpOS2tO1ppfhMm+ueROkPKUY+6C89FlH/mOYpxgO6a6usP
++NS/7iG3exBxKaKNcK7JZmDoxpOzhKOQyB+cQ0ac5IIy3LZJ0js9uTh5pmSAF2WYKJgQoht4dVC
yKa3W/cbUHbbC93Ow4zu8gpF7vPtDARmzEaSkuEu6qqimozpJUv5FerU8mBXtOKqoWW/rqhhqEOi
tCvKrRsbt4uvOIxgHqv0Lt6k6rKPLDxpZk+mwEtD8Fj+L0gT+s7Wh+l2eqHwhMzRLdYtHbux8NUh
F/3vAKWFPlBFEGXrhw0t1GQGYe1nITBzNZ6ek11Geh379sQf7quKaM35qr3Yj5m6guiMz1ihy21o
zyJjtZiZ9n4sILhycvr2+XxQpxqeZ311WEU+VmeBK8/XIAvZAH2z3itKnCo1mEAsczumXGg0kF6W
e31aB1jjlcAqXopmvTKWRMjhTegignf+mYZjwaRGkj+IF8pKjZQQPyJZ0L+Ibozt2K+u4Rs8gDDU
kNjB3i2PPoQt5hYeBh8wtgpHQV0usuxzwS5dC0RFeOtnPQWwMUO79bUErr1M0MepDY8L33p2RjD8
QCWcuppB6UkyqWgxBQmGmz4XGrstWymxrJKSDhd8WVv6pjB8O/oCpBALYsu8qVZGYbWL2W56cWR5
IP1HeVZ99p302aiSB699L1tevkNLDr/kR2CzmQFh9azHWDAZE1PoBlT+jXA655Kt5tfWQDCpX9uT
zvRuq0s/SQ8y+mACcZnJgenoSIj5/+L0na/VaMTYGWjRPPCy2D7x7JxCPf5zmCQneK7Qf8b0lfWo
O20VwYIj84P9CmGJ0ZZG0zx5uHw6hqQZEBAAaqCI/lvxy4m8ewnDcN5t95gUx9HNvZcHuRDzaz+Q
rO4siXd+hbB8flY/VuqrYW/sHoFnqE12X6Kb+7XeS5Oo99Un7VgtPTn7yU85mHOhB51JdLbwMBJM
bBJhQ/sL9NBv7qujQZ57NY5Xdf4gGKMxsm48gwmzcALJ/4QdnubDfjVVI8eM7jIuSC2PgHmu+YTG
AP7fKmS8jV4+Uqu1vJsEIDpKlbgl/AfmNWX7H3v9Fj10WTN3l6GcXseqyJRxDe4s7r/IEFWQWxuT
zPMDfMco4ArhmgKfGQebtx8zGfPTx43rgROZ4MPD08Cmqss/xsog9ywx7xkwZdNKxvvc+oOE2yqP
AbosZyi0lN8speH6/JxbrBNNRjyRQmsm0roZzKSSX627h2XrqPKJYw6ZsOv3JD8uodb9DmIVGTYZ
DSAPCt4eqGE9lGKhMvNpJgFiz88Io4hL+fZ6q4sfmO+Yh9GfkSJInch+rBsJYdYZeeCHXqRiS25Y
GZpGBn6vPKRIUR/rgJB5f2JvLFB9r4szzdCL67o6VpGcr8XEdKdvBhDljpv72OFyu6Q68r7zrSaN
2aEYq4mqP6PWJNZwe1e25whyiG3NGQYWssSN1G9gywALxqv1e/D7EqEqsgMSAsAToEIrjFX43OrI
2rM/sqllDc0W9NQD/WtfxB45lXlS6oANmK8VHTj3hvQc7xx+sTZChQEEze6GrHGM8Z8eNiTyivB8
Qy8wrVh0RBH2SjZeFc2WKS6oejVfgWSIAL+Bt8zaYSRlGdIJ8xo44QZHz7hSeU3Xd5EHLIZYLn1A
XURck9dGIiptiCSRnoKv/wggPCIDX4MDGgN/MiNpHuXfu1wZEliHIt5sUUCxCtKB7kw5k9iql1DE
PJZ4RVrgpeF0/DnQOGZicC5Z1UMCAVD4H9Y1Uv9KWEMpQy8u2Jhr+vDqtW/IYmq1C7inoTN9yP9V
zbHWA9rlyNengRUsUDM/7lr/OEI/iuaUpQbc6oSKDdI90i/cgWSIWZWWtcQpgJLDzbEj9VwKvVUw
izji6da2ss7e5IyRpxbdZYSLB2zBEtAvr/iithp0Da7KRS9HB6dnnXR/DPKRU1jjZ6h2rTziYe0B
hIyThu1YYd8Y5m+FpkJ/9kBSBFM/Pif4NR6I3HJ1nOtpY2tPitJRp3C4tQ/qDXNFt514M1q70cyI
qBq3AVIcGKc3IOT7Lg8fMITpXjsmebd8nJu0ibgRhmaLfwLvWx8SH+UFfcse0LR9Qa9HqwoZQwI/
XznyqfWk8PLa1v71P6TN4i2zBBHlWPbAINl2SltiUFVl1QiteWPVRcEwVCAo0hxc/tfsqqTZqG+S
pLYm24/K4qFCTrHxqkryqLUca4BHjbGHwig2FB/MGJs/LxbkSlbxD8/gyK1uo9HR5fd0FENFeDWz
k0lahtPKrP4xLhEakg3qcQWII7hvfWdNJ0mq6V3mLZ3YN2y4B+BzHLDnfkzggXJ+VJfdI9aIzYZ2
TyH/oQsDyUPbUHixkviL7NuEVGV4EQSxIDszamy0DNhqvVWvrbbNA4E41U8LU22sS70IlRc5I53U
DuIGAP6s2S/3guDvpDgh+pnJAWhwLdTVcmIky3iUQgx+SJ8YLPRSVHMzYp2fM75nha+wsD77dNOZ
YcB44azYo6Re0xMK9k8HxsBi0bDB0rWuo8s8ISyjmA7GbXUbJE+CMRVQdNkTWQSge2mX2eoKbYcz
YPVFRLpIInGdK4US6b/VZAikYDu20inSbKLIa7aJO2s//TTWaMx1GXo4EtCTvhi8BH2lqnOveAHG
cZ910awAufgaPwb5fcEyhrU9jzVvSUXSZZ9ZR2XTZtAzpdpma++Vo6ShOyUREkE12rp9V0sAycOX
kdPvfWHoYmdyFmWTosaRUlQxjPTODDtVJJRxS8wa1vmFr3aqCWj+L7WbqLFBmg3Dekj/PQChIbWO
0L0kJKaf6K1jLQzg9VivY9G0us7h5SFNh7IrlC4uCrOZdXk8ZutbTagnCQrsonpn2CxWueYBVu0p
laW0KURg6qJ01wxsW7CbKFFsXLMqkCTmiQq0CVcSVosOLcKKy+FFkg5kzoUmrojutDPvk3sFZk8c
ikqRFE7GM/P9sfZ4+zMEp4OQsW/+QpAGOLnEqFiFOQ9IAnVSZeU1qv2Q1WO3Zks1t844evGryJeO
xJFAidghyYAA37EgzycAFOApeDubsXD4WHHL5QtWGEoS37iJoEPpSGRmfzThUUcKmCJsBdnzpl42
AUadMaZAkVLR17T45kdPMDpkmUoJJRQwFykcVVNgtuf5NhE7u+FUGEKClpxy+O40B5O3ZmYa+v8A
FXEw/9xMIdvwGNo1mHFdH5mc+IEI7isaIRxYOJUfWyp8jJ9RCgKadZ65fXtP9dOULNp5SMCiGKyN
BPRip2Q5yLwvnztfbVXVvgLgsLX6dl8rg5UNvvtLi4kMID0TRYZRcGQbm+9lGok6BKtEgXGRXl7q
KE8mlCo02YqM69eWRZWdet+UaCEv4TUrLKHupIaBccO/vgF3sZ9bl8EHxkgq9n2mUK+PTsNdO3Ng
h1d5cSmOU+7nIpZuWNyUEDnRVXKpBYZQoVkDBlS3P/I6+NQOgZCRESk3ZNuyxgKI6z5MxVqMEDUJ
JL6fJUm/Xia1rvbZTgNb68rtzZpwX9NW3wLLXHqeOIndVMFQI+UQnQAAMrBSFewOFR1CtjAb9EM6
UlK+XWn/Y59LCrSJd4Kyeo3polL2inN4NnfDMP/PT+szfeJqMZnNl5JMstPXT4RwJahrTJa5ZW1u
Hok3SKw+DVeMtDrPr4WaKSjz7BjsjAC65SBBZfUrK5XdrtfMki6Eaq6QcmedgbOIIczOpNXEO0gT
WEKcw/52kH+ZhbyR03qOAlIPUmNsX0BAZExvFkQ82DprNL0bssPGMxVc9DXvabXiUsCllDFqkzEm
VUmOzIvljbnUW/aC0U+4Kn1TVqFHPj8uEAn/cy8TzT8fa/oYLYoUIiV4hN9+xVPVMsPvyrX7Lp8i
CheAImbtZr+1Tta7Twp9sFqT+US1bRUFiSAaZEWyiBf0ilCqoDIRTyOobTdKjkSI+3iX3CbL0SKR
kF47dyAokfAw/3IIeepBz8F6ro3h6C5mNvgExuqEsn5XMzIEmmrbzb+BBr1CskLtl8yJFBmULT9z
lDSPgpIfzRqrp00kDJPDgoPYPAxkj6YBxczE4egmtdvTGsT7E8lFC/GWNypO9/aIYVWXU4kXmFZZ
wQt6yNoRgho1r+SBUzFEq2b8rJNvdi6aEmwmgXpSclGJF8H5vA1ND5HZB/IzG8V3C89pEhV2cbDG
f5TNIpG+7v1NeeURyE+zpf1WjYcTwE/Rt/9jxpb3mUoD6mWASNrDLRbS4519IiLmTuivnh/zuWZ5
ZmibDk/pkz/HHoyXsLLpxH4JMHwmDBKd3R7JSQsG2SOxPYF5ZOAtWwhWX50DR79F4CA5BziwqNMS
K8hBUHxScd+gT8mwyZEEVk7x1oaNY7Zp+SZKqDk17Nr9i4Uvw4qdOg/Ad7kxlRW1Qim3zyDyHUo4
9Y9Pyqq+2nxgDkpQf9ck+Vgt3oPvgUNq9NLBxTmYLxE8h4tshxTopn3VFMnKGAvZx9kcU3/+QoF/
xL9q/IFOBiiiSHEzXbtkt1M5UgkQAlZrwIBQ/kIog2BmF9S94ZBWJPmhSECI1a3N+63cf6lhtkyG
QDuR9qWDy56AWsgBJN4fHnWUUaaRoKmiac6TOFnEZ/l5X0z8HIwNY4CdOHJZ5IXul/tYn+aVXcq6
TTAhukBCY4D6n0beDZIxyit2N2xzqlMWlWnh37amwFzyB33A7sRn/i2OpuJNHy+QvaUxAdCsErGl
8jCg3Uo1bKZzikRJPQw5RU5iTwri4/0kgHOpJIZTyuTQEzTKA2UBkI3q0WIzUWvNHMtz9Bi2B1iw
NLXemcHUfGgqXeDCkYj5mFoSW+mmTZIk1AGv5hj+tYrv+nKbr3XUT2KUK44CipuDRp9a13kJfgSk
eXTzD7Tx/SyoGvPCpj42v5lC3MTPW8eaHM/nxp2hhozQiCj/EQIL/Y8h5xl5NQlx753s0gSgR9d7
UMcqxh32ZIjzxFmbwFtdYOd729IJq6C3e9ks2zyWub4UPL62LSaRlgeYpt0ZeDaO1IymJcvPJDDj
NrnWrPnEmjaU+kSEIQ4sMJZBx0EoC5be+SKvNcVAvTHdsHPzFmg5pAi6HwLSFmIE+nsR6FZdThAZ
AX17tuysoO08PeA91e+blTcIpoy4Bc6CgysaVovKOIr83kS2FmpmvHSx71pzU5/Z1j9/INzd2cji
rqR3ceIOLNQORMXikDrkcmwXVduD3QLMZ5k10z7HRSbNQawJachxW8MD8vt5Z2z6qNztIntBQPJu
MOLgzuvPW6q3RkFqiLUxF7NTj8QLg5YQXO4w+4NEThxTVDINnpCtdw5SRUxP6t3nc7oFl8bsZjhG
JmW9122IrbzfpIfdkZZiqMVAQjiFY5tlIOA/N8gTNpKE42fihgTVsGomBC6Y7FvH2pKDEHG/FA9r
EmkmcAGKbJ+tdql+LbQvl4OrrAvv0KNAl7EWvnHOdXilRVin9j3HjS8wQtCI+K4qJpUnIOdEJ1cF
l2FeWLLnEpUi1tj5dfj5vljijMM5eiJLXJaEz6HjHqqNWrLKMaduBSJxPi9flGsQkMA1cfkc819P
AHXvWBXQmHUph3BA0Geu+eBCySVjCCV1j3JAb3UJbE/xjG+X8Mh9ERVXFruL2hgtLiOXOuyhf9u1
0HlEijG0zBKp2MAPoXtDd9LL+ac0QHnuZH54MHZLZ6jBI5B2NHZirfaohXBxTMoqJhoOsJQMSU63
EBeLYYJlTGnIUTzUh7m5MDgpoiiUnYLxqYIBSsSsbBzuq7rSNgDY3Oq0eOrz9+uc7sdX2lbJu7Cx
yy6JxPwXQYh1ksdEsuaW/xgfwBjqlfJI1VOqR5H/qkkypf0Udn5gzvW52IyKJW1+Wn1Hzk8Tikel
2v12c4tb6F1cl4rqABYD3cIfa9ReAvhaUHyhRn3+IPnex0A+E8YZik4C6zdghcX1KB9arieFdD3h
2v/myIGpIMorf3BiU7sDWaTgx+WqAUQdSRek+9Hw8ke1kGl8Z/Zs9LVNOKb1D5Xpqy3kpqZT45gc
tR8XkxzA8Ozh3xDFS5YS5nOg+3/U0vpqsU3wj6et4mhIkZo8EnpU03b6HzzVOUtq2QbOFCwH8ruG
Fpqcvnm1SqlHz0LblTgGGfWPmVkj7mZi0wg45VWnSx4Oef2soZH0l6CKO83vSdp23szTcsd7b4bo
N50u9/ugiPDRCWlgXX7bjGL13GAxxpyOgr3uVqhe73NzLXPjPeLNbzU+2xRbF6EhDe2+ECN7idTK
Zh0xZ2gqWZk+YlRhlC5tdJYAljaogBXvNTF8k81bZOfuYgCT0O51/Ge1yzCkxIdKIEaeYqGboOM1
WCGjBYWRxUSoYWpvnbiXGG00sghsPRYMZW6Fwwfkp4Qf6nCauQiZIPdZm6vlob2VkYt7dQXmsSeM
Ly3YqrMOTEkSZQZbyRKMI2mJWyFEkirpqccxwmuzUDCqajiT+3RKzSSbF+BVRW3hcCYZL6PrZZTn
0S35xzzmPoa1bb/VQVWHqRCVubKgeHt8ZM5XOaxE1/2i6ZAUqkpRIhr9zWCOWp5/g4Ix+A54gUc5
0fK/qSYW+INWV+71KSUQsD+LI4CjreKU+8qMVYiA/X4005UTrP+xFZesL4SBvBwLgIFuZMDVAtU4
+rqdaPq+uRE0R0GA48NdJrSow2GJcia6MGPok12zv9XXgQUqElAmap6ddKyidi0vURhkRCUYsjD6
dI61d2e5i77pjCP+jiwFLa2fnnaKtM40PUtlxqY5/iaZmENLyPstPzmFxPb0znvF3tQo6I6CBkxt
kH5XM48IhOMg0EqlG2jASr8tOuJIAkcf1AUDWwCo3UBYLiUIDdq+8UMYNuwjvT58iJuhEqoDrgcI
CwPMK3kWR4NSuSptaEvLqq/naR2gsBj6F5lN+uEojwbNv17g5lO3T7GdMbNiEXCnlfSs/GU841mI
t6pIMcrC5Q5rtb26bTBeITyXcLrLBmP03FBVewWqxEkwPcp4knje0O2/LGhVfvSgx8ePMdV+qsYb
ZV+5nXT5GQwztzU5vxyNvMps/PN901rEiT7PrslF6PTX+euRVWzqFJ9nHuWAloanFaLWPmLfujYw
hl2fJU3uPZvAeBAjBL4KQ4GdBAYfDvnE+CxaHRFgWjaBWDxQT5TyrHrWAFJPHtx5G0XwpWMMPKFw
EfTBmtCCLykfr85meO+WJvIUyS/yNsWe1opuNxrvaU1zUZk65dYLvKKV6jMh7mk6mKiY/szPEFJl
3a31lofV4FlxfUFw3mdXoRs5k6kOT2qN31DIZASPEaiNz5LQVh5O8LDnSc0ZLyNyuaYwuIFIqCRN
IGNceRVZnEuNZIDux96tOqz8fzCq6Zna09Fiu7H9Dbbqng+r/1G4Bo6loyDS1aw6Szua+1Bsn1kZ
d1Yc3pzC3TXOJQ12JPkbxn1chA/YcdjViQr13Kc/iSnSNlAhE5j6EMgED+HVZhFH0770wCM5oTs7
9LSXM/czK5xMPjXYvKgv6gxLxdcdmWQit9QowYcUyM0gFu10X8K3i8KQT6Iph9Sim4lBQ4h0OsGG
YgjAxWvzbCfzxF5eNuejdRro+tEqSqWIbQ1oKOyQRPkcqIJws3hZ8o49bPQvOzgh+k4ptBoo7nC/
D4OxDtPU1C55xCbiBokzYD4qPDY9nJ2IJcsRZ5Itt65h6FgH0hHM+76qI2+ogx8X+sjr+D8QbfY3
Zb9WnNX+coE3igEzmToN7jevUneebgg2pjzgNrvV3zZX2Xzfed7my+dvcNX5dIGPR5JT4JUR+pZj
kErNxzH2Xcpk+JRF9IqGg6Dq6zyy7B4I/c7MWC8zeDMeNP0SWEhmK6jjlZRiqjPcktAiDJJwI3us
WW+fw8OHIXrCxT92ZkQtw0Y+LaFAJHcpydWxOoFWTsbXGuYxd7hmYA/yvHMlfo14FkukkR0w6pTr
rqEnQSUGwJk+P56Go6EfMjOU2E2bxyEuWPqHM0/cVlWaZzKwlWz1To7Aot7wAMVm3B+WXs0yuE3W
0L4EkD1aJakkBTgt/t+frQQpzZFDnRhEhd/MUFse5YVeYwknIKG87hERJgCxf1A3XVSA7g+BpwR3
3aLb8cB6dQnFpSgBmdu2jNgq/Y8HIG9xGbr52AffR5lBZ6ddTrBmLB0wtkxsPEJXKl0iP99xgYfy
b4ruBxSyYA3dl1xjJFOUUPgN8bLXJxhDfiWElhbVUjwkDF4n2AAg/F0wx+y/oVFVopVAXZ1Zin9S
ow7gGUN6DhIla7eIE+GII2D7Hxs8KOZMsY3ld956vS36bsmkhNIwVgnhrX1W2iqgZHwkUqP7pLuJ
MC7fawOapNuDshfPAq4ThnnTPQbJL2nEzzZHMMJacVtya2OT/TXiIJJkX28lGtxNQ0LFN727bTg/
bdXmRlrpJqXu82w6W8OqH5VIiBIotfystpJHQwJgfmJ6oDe75woRGnKXehNy/MYS2hIkuGQr7YAH
ndvZgC6Zp13u0F/0nruhIsQ0/ton4MPhJwMo7yyuM/+lyl+cIiMK0iog2Xq/v09UR7PUoL57ZL4y
n7RSgm4gKC9VuPuIIlt9iUlqq8Qg2/wfkJ7SDm+ipAQdV8/MHt9t9G971dcmZPyz0Mxr/kenNcsH
+eT0KvL44Iz5Yv1dmpOiFrxazAsoet5qcA0YK87gCgyuVz6EdKaQoeFwoxpCZifLoakJOVOm1ua2
jeQ2CPMkC6ewzO2z9NOPR4jmdQ9WOWqqQ6vNRL/42I22Ws+75NpNPcCiG6Z9oR3KavRVifzn/O/S
ywj5jbd860DHF+dzHQ5kZvBYj2f+ZtvmrXQSrQfP6/D/5zSypLO8yuTEDMLFC21ucGir4fMlAE1o
HLZVYlCsRiINoHVQ9ckosn0d7bvqq1GdCeAT6T9cMl7mHwEHjXsc9i/RBmRzeSQg/ITmu9GNEvKD
jZUfCCAb8VfDG8l1HH1WEnRKOKJA6XkcuFCd61xhHFsJQtIaOPzrqRpb5wnhVr2e2VWdQVG3nOoZ
EYD2mpoFcgcVw4neubfSBFgRq18Rh/5IMHXqbsV5zHM4JVlJy5pGG/r8NNMcPNI0RNHCET+/U6qk
8hJmrztipUv4SHyY7rm1FjslRbUUagBvWzwWkWO+1a8cBin3RIZ3LkGFZ/g8AXqjc5BBa9olZThH
eBFbeA7i6LZ3FRdPHgw0k5lCBR2sG3bPnTKSYenhakDeujBtrqcSnsrQL5FvA0irLtnseJ6mnwTP
rPmisg+Uvi4gJlAwAvXZq1FFGG9Oim7EazgR1QWRq8cDY+GVXN12rkABrDS0MBkC0ShGPBJO/qJQ
/FvARYK3zmf5hwPclEWwM2md6ZtMoolT3bquIGuZggSup7uAPXFCvRRxz5d6+abp70c9hJXPzkwD
pQm+qA7xc5B3jb4XLQQbF6CEZgO5BLiaHuZQZ/YjwBT6WVMGbW8oh53elbX8la+NwPn9AH2AOmFX
qQHfgEhd+o+4Jq3zloBxjN8lLyxlnTWCz0S18jb+Y3xy0U9s6+RDKDAVVo/7sVe3g6/5yjff2JgO
p2IJNCDdrLPh0SIMTLExS+59Mn5ou1NtnVUD4gDOccaS0RnKMq6Eu7YqNnYMTJgLnOOXYztSljqT
0y+MW3RPEW+REPhBiLcBjrMSqrlKm0R7CVuKw2Y2DPYMjzlwyJan6UU5fSLGaijpx1iAtVEoFfCL
E0ZlKhAhK9TrvqwvuU0wg00/+Me1amszrZjAizH/UIOn3LfmqYIFJ5IfAAYO+PSV1g70YImailgK
3C8cSfP8YgOd1YsY/LB742oJ4ALECFM9EAztBnmJqMgERo1QLGcSznMWRrCQn62Goez7fIdRjtY1
/H8NlPza+cRK3RShmcOCy3S/fqF8D5JSg2D8pu2a/wxAwjxroc2XQASlPVMWlnKmeJdJ+H7MXcv6
uzBQfsexjRjYgnCSi8mDUx1aP6mPXX7y9Bs2XRwAx8LoF0fAvTxZKNIWMjyLZXQM1l8/4pwOWQMe
HGmDo4wgoHkXmbCnFDc1lNAcX+BiVe9l3JKdZAk9Ts2JvbP+JE9chxUFN1xv9Rk1bzcVQOHignxI
8blPotOhKbSqs7zu/ydkxbn+6ry89Eo2jkA5w+lXnmrZl7IVT8K2R9+tnP6Oa5KVceYhiCffdR3s
kdGleSUYbPzi9PWYUN9NTCrFAUVsVhEyJOYHKuzvzUuvhshgsms0o+5LFeIKxjI0FPHxnyTDhV+r
1CzAauiXWKXoSP6woLVUOrIX4m9Y3L9cVvqRPW4zVlxYpMe1oVrdX/dyBsDW8bKzLDa8rLl0ShgC
2/sm38E28Xg7ZzfAJMiAcJkjAiU7Z0Max5Dd4a1D4nviWvbvN0ySNw+9au5edocIEKSFVHmzAZIE
tpt6wbquzsaxVP+nOHtgNPRbGcXoUMyW7VLdcKeNhjSRWSxOk09ml0+SCAu0rd2py+cMdZzg5Gi7
SC/4u38J3masIdwxoCjgg91DF3xPxA2/EGJkI/fNEvLCAzAbQpk+irLf7cckIUA02VINEN4JYZlI
LGZ9cBN4JiIyg+Zv9MDo8DMFW+eTlgWvwV/kmUxbiJihRIqnDr6F11QkTjSA/CsFqk/4jm+KSuH8
tv2mGxDy6pl0t6FQ5AcmBhw4yq8LyVyc1JivAYOLWreVxC92cs/eUVzQG0Ir0s8g8e2x6WdA9roA
mx0xsN1rmqNMzziOs+Bp/vqy9ovZI5WeBm8FtlOfdxDYQ5vY+9rjPCJdrwKfMF8jZSDSPpWWyFwj
BCcq5Rz4QPVZ22yLaUZaxT+BoZswXHvpjU75D5yJxtMW/4ncW8z1WbnHWRTvV71Nfgf0TIeq5aQg
xCEjA0NHWDRGsq2Uy/GQWwD2ZiVJxfUh+6jfJH2yYFF3e+iaisG+8zh/eesGNKWhToyCFafFVjrU
s207jWAt9ikwatbou5P5J3Kp0utTeL2ED9MzGPr21bVpowaNeAl6sd2e62fjVFEQhTsYpRXIvVrj
GNcge9Hdi6LFJVMgqgBD7FV5ZE06bGEfin7jAeR9a3YM2HUMajFv/sQMD4IVt72FcOilL+4hlNsf
U0DiIl4f9fDBNDmvCvHBlSklHg7o2/OPhnlkmTrhKRie1TJ3zGvBYHOmYypcGFW7XUTmUxiDAmaH
AuvBjzA0tBZKtHkjaGZVYIeFq/+jd/r33SGF7Gn8omLRLiZTFpuAGA7H2AbK5nEENZo9nKNFGHEJ
5QwrUejej7v0HRejjGh908gppzdZc3g8rfaUpAR2JEoizwk+q75WkfMpWRk2qLm14PXNYMOrUJil
B4x4NfL/MZ1jzejkWgzJOXSac3y8gsOY+vs7YRulHHqIx3xYED/XSdgzDRH1bHQ059AOls0p/npM
Jcc6r4QDKL/Ing9/C0AbGGRVrkbUvnl/FVprIyeMQ5B996Guz1NunaVNAFfcjUz8MJrLIqRSsXbm
kMDtzoo7ciroMZU3CFCNEs1zyT+HYNOADTICAOyzKimYZbQSJZHKih3A+jTtjB6DiIN1zqc07IUz
rV5TPFivQUHlJsNajtkGsqQ4l2ng8AjrW1QCp9GDJlJ4n469mHyybScJhm8JyfVXjEGbQzYUSdAB
c17ZdrkIWgdHgEuPs6NScrDd19WxeP6BURKuTnhkuLrynYhJstj4Z9itjNuX/B4jbmJVFPgl7yay
xNT2tFHf9/KRbKDiAofoSBqwSnmKBURG33ZIXMXwDBRSxkNVKAIis9rLo35cmO2QJmifAEIE4xpF
JTRdcFes4r6YUzbFJNGyDwF0dc+mt/wUZFm9uUmt3xX/g5NAz4NwtyHp5oBng6C8wMwA72dADjuF
nsPFz4xroUJYGF0vCyZ4MoZj7uBJ/FyJGNZ0gGYQ7Y1g6tqw4ucHvEgDoWhE50ifMnk8GNE7fgXO
cT6Pv0XWGvX9VJnI/Zb7YhKRYJvoPMQ/u7q0LBbs/metb4zGQe6HJMD7TXQLaBiJ5nR4zOLFlT8j
DSkDJp2oaZMelT6danFyWI0Br2RBblADYGvJfUY3jEE+XHASumkY8rvKxAMjaKd0w6UJufRIIS6G
j8j0H57OAi5OIsJ3e+txXp7kYATKpY8T4cckO1cZK0E3Qk95XnKqY7ikrlJTjC5KsC4C1pyAfqUO
Grvvv87loukTtoPLKzJEqwUj35UI7i7bYcZQlLR6E6gmFZpkd9W96FifOCTfLThR/55plSRvNyYp
cIOLsbSEWg4mBhpyedO1YIBEKGpqM+wlUbM0pWKgR4Xkr1EeqkQxqlWf3BUGyLsjxwHoczftBo3N
v9JBsJ2MV8kd6RIupQUWYyu9CWQn9W4yWaEHsUXkCbUp9FHh1pDoO0CWCfeZSuQLk+nBnEOpzFe9
UnNd35UKpyyVcOZD9m8UnIK1oBzPDt7GWQAOa2KIrUhqKm+kggSHkZBNTcz3C5U9+9CsBDt8heOe
SCt3FSVjrCVuPIwvDHqQm9ztdxaUhJJnNaeDIPh1J0hPah6PAqxDaGPGH66tb+wm3frkb9H4/9mK
wMFojL1+0kxDEUEGM0YAsykbZm57VOIPRx+IXPq5iIu+HzqlVU/pB/uW0AG8Ajopmu+99VEAOcNJ
ecuxegLCaaacGPEzvH2FYZiBZyXthryNvuY/hXCauDUZGYxQsPxFvJGt0GOOnZKhEextX8Q3cxzR
12yujckf+KdePooyEbVaiHXWC0+NFFQEHsuLd/xestBH7J3L4YljryNpkpAi/jg0lKLO82lGiaXc
/KHfnL2lO3JmrVLqMt8OKH9F7TP7qmyxb021i+EuVFChjUss8NrZS6Yw7GO9WJX98ROeWIFkCEVv
mNoJal+aw0FP0SEiodwdZzM+viV+BrJqOrxCV4RDkTPj75zDckBFQaQTEHarAlm1QrHcpiGAJKWP
/qRJoYh9lCzNVFNSe7oUzYx9C7a3ZfNHwjfj6cWzJ/vmxREeYgHPKmgD+F+CamEOTZT8bSwKWbx5
vMuo9DKehCVH7NDP5+BQK4n/0feqacR7G2NuMZswdD96AAKukrEz59lccFrbR/CVCF6wVz3K7AXu
kj9WH1UB6u6ACSm4Pefd0oz8UM2PGwxKVbZ3+NDHv4uszM0/EkBwkFDZP4OZO07B7eTsX45/XqlP
IEsifgE7XSvuYveJz9Y+HjQk3G+RKZf0OXd/ImY749dOtkKh17Ep75EZbcr8I670yAjdJGn48FtX
GECaRknxvYjJ7Uv3u1ZMAOmpLbu20t9eJdS0YqzdLB6qsEBd3AJT1FEdOZ0R+fYx31kV1DlNkD1V
nKvHod5a/HLReE0wHIKBocIQlgJ5jcSSqI1JZ4qC6qvIwCRb4/VNDfqmP4m/bYJcBOPNnO4Rp+u7
32G6+LxCKDW9Ac3i6CDRaLpRk+er5zyjXw5ALfjlg3rfarUYiQYjJtREjxyXgzrTa8iBFs8R9M+p
MeQuBgNplfmU0KRGwmDB4vkLVafRl+usxe2wfgD3uoww5G4qHjyP3ZhVP+7a/VHrrB6HKWtghoQd
btJex7G0K4nzmseRlhA/Vu7/5g2KP7lsljmTwdGWZ3JqRPO2UAyUXEdeYcgTbqMNzm+U8NQeqY9a
flGzVunQwwGp3Hzk/ZFHM5xKRREkdx0Kqg3lNazl8xkAasJvl7o/vovWJ5J0M8E+BLMembDc8VAV
dyyyR+aCxnjC9ic+VoM1f+Y3Ic9bbOG9l8F8DMY/UVrW1HUZEhFnsb6/kMRFSXpLcow0+kvWHMbb
mfLiXjLCYFvySC4jdzdcOZVDnok24zUWIjhZFuuSAss0as1qecfIa9QUtQD2PjGd/EA/FC66XJtY
zV8GjU0sWeNkUcg1qW4MYbRVb3I56l89AiJzXO7SkWCRWIdEjEsXsxTROyQu6NlOIyGxjH+lnUwM
Lj3si/1WWut3k+2riTO/NcXueVEH0XsMq0AkS4CXKYvaie4Tl/YxGgPn+tbEgkpo/IgqmFJpdmyW
QdnPJQtB0KcbZBwBwQYd9ne4k9mJVSQHJ88hXCGPt/UpoHdLFxFxS+Owz41VCgijfUmqbm4m4Sur
ZCymkCELJvIAXrMqKhH8IUBE2eEK5NByNM41R+9EhlQpuxB5VRs2ahJHB6oqT+gspZYE5MWjy+UF
dnW2aw4ib3g6PPFF6C4F4u9Mg/w1EttYhUo6+CXK8UN5Q6RIjYQsnYBmITuVsXKw6bB3Xr8wsock
kh6NPAscFSb7FyaiBzYRlRlj5uYpT4FCCwigDJ8A/yJG+piGt0ntSS9ajlP3POXdPXEo3bnK8qlY
GkOLZ48CoXSVfINzvbrUV8IyU+LWjrSxGuynLlAEieoKa8s5Life63ReSQs/TDSvq4rFTTt8Pz6g
T0r4LbLCnIiWQJHLXCUnxpLh9WZG2Y9nmq38SLMn00vwnqLlnSPaYbl0Mmh50j9tnQcLOMDLTOxi
eHloB7dfCYf5yokirpDVXLczI221T+7kZz7yXGRb6JjcORGpd1k60YwvI9HZtK0iMXq2hUzr+Ba7
zTsN/aO5I8ebyya1uQodqUxgQXP7i/KMeDTO+6IrAoEzAWkYv+Eub6ajgpz8gYozMXdkrxYbGtWl
1roTA+bCXmTUg+QWkVeAD50qeQ3fWxDiEjNJstGGXnGrq3YAcb+7jNH49d4D1JePXG5B9cvzDdIN
RYIWhQzVLwZHPBIT8Z2WaaKXDAqomKO8B702ByO67OuwXsrwCYRxVPyYZ7zGuJ1DcWjn1mZLpDVp
qWcM1XCfOprcNz8AzzpWtFkQvm7imWwfccEaJV2Vcl2VaJlCLJMz3MdY/CvZdAHXNJPkE+wEX7Q8
Wxi4o2gax0zDGFqAUKQYs49b1K9RqHkJcSmpqBAWeN8NBuFSC9HUoUa0nNNc1nH0jZCUoq2YpSHD
6jOpMDOj+ATedcHjd/hEYcbLh8vjYpwDaa8oktVY/LHS2Hs0oatogqFpvSbgWculWuJh/ETtfnp2
5tkzOLFYCmqJqX/lmCF8owOEZHe5IYt6m20Z3NBpXWf4RhUngntexfy+Iu72d57U5OVMI0BqRwNS
SCr0Ek+9y82aucT70hOxJuqzkupakSZTNiRPrSpYp/36+HqJ9YzixS03Cgd47qHpOKgNNp96YvtJ
HQC/rymcPnKVdaiwZ3iswIc7RwJpwBn6fvZMMSUMklhNj/B7hdkMOV7sJZDqntBACvEO5wIT7wyE
5UXwaUYQrOSQZ4I1zhaweo4N5MZFjqmSBpLZa617BRYeU3BA5Ny5EQF4san4x9tXxpDhz6hdlB+k
yL+MBFzdmsLh3QqxdEjUOfRO5Nam7Txgn7o7O1glB3FhIpEcS7iFaDHQwXZvFruFWIQjvgxUp3FX
I+QQ+Ahurxo8+3MAKggGf0OA7Zk6LChS+MY8O4CmCyhy0ohrRtDWr5344fx+pru7KWPq6p3cTSqn
TJL45mYVinpGmOd4C6rKz4IDdG2dupRsrY6GI2Z6mN4PGSDF2RR08sGJKnAJJ/Hb1NuZvirrEvIo
ibhN7hThE76cFEfVWXpHPchsHZQrBvFs9Jhxw8Ye0B/V7wSsY+yfg8riL0AUUXSoLgRePeq3oNMZ
SAsGcJlL7kc5zD2bcmUOlmzopTzOzI1uPBUnCTiPVic9I7nAguxlXYd0PMFUAIZ1hMGAtfnvadcE
RUJQyqrU5qF4PKKCF3GUFp6sF1bvg4/UPgbO2ulh8YPHCTVbF7rbsI4kdKx6t2nedmzxC/gkm+QM
6dhZJTZ4d4o4fzTo7hIrsvcU/2WxvaCYSGHlucb/0/XSdjkIf2Sb3pXeX1BBXtcWM9Ni9C9OyEw+
AHEi20v2IehkEQhK+7hHKYdnU7das2su01tFEkHh97tywqAMJKuZBL6VTg02O+i520ps/FcE5+yM
sq4w2odmEjCDJILWwZLb5w4OTdl8EHd4jFMDbCVz7muSn1a+KwVBpt/N8VDkQmfqpql0eRXrbb97
eDut8/dRUxWjmXID0IepcLxsFX4mujtPQjctJjw5mHTKOxBCd9xhMC9UJN4GmNUqfe1r1hfLu4d3
udCGhDZvQOmRyo6ftC5kGvpvL0NohLNAHLRZcsVN9rcbE68enbBBbm0LlhHb1ERN/3GjhwUm89We
ZSMSenWp0axWcrNd2fevv/1c6HkcXqUIOj2CO5JqX0bolMzRU++CqROmWdqX6kezd2MH91t1r6iF
WZ1483Akp/7yNoCY8iHx1GQI9WpOEg5VsjreV6sr1V5HGBfkrjFiIb2zRP5TyD4QgM/MWZk+zAZF
PL8dLtwWVDddRtzY+wsKB4yr+2G+K2dNeLtUZLCLXofsdfLkaU498U+W6puldtrDPHbtLStBuXPn
0ApFEjxJxz4xvJLfDtiXz01shakvDWjlopDPMvmsJmUAswt5vHtDS8y9lgjs8H7pg3GJFHbqB0mw
ErcVE4CUfqdRSP4MiAWWzcsr8wY37m0zoDvy7LNKCGo2v/NJM1t6gJE6fgytONaID34vFqWCNk1S
FjoLVR7iNoBRuOSqyVBbr+ndlwHOwu7+NO1hLsU58lk83p1UGPSrotlS6cxIA6nz00LHdGl6jDpz
FFtJHQnxzZTI5zJq98rkxpN/MNG6FFd6WzW2F3GYABmjmmwE+kAit1Ul7VXTe4qKun+jqUx52qJU
M5foSmGrVHE4ZxdSNGH+mqG6/nYhahrHiozu141AEBNbsqw5P/uFLMR3IAFpDglCOHyqeUoZg/J+
cmrKZkr2tPAmJdPdZwLoJ+Zg4uEk0fSVm8AEcEB4HS0MPVJPhPPqaE5JUElRRbyyXqNAUYWB7DYs
JF2mbntYSKW4b/RXfWQ7bfJOUdc1F63BvM2XAW3kgWAqKmlxFqn8ntqn3O+cQMp1LVTESrIlWXQh
msNJtKs38oiC4DSoFJVgE4l+8zOSWysoOtSFWCjaZia4TnlVeq6wG8F02VwiAk9+xH9jF7rZeT2c
FyjWem6N+qzKGY5Pi6tuHwIZYESSBR79hKhAYaH9z+W4x8RJMKyOdss79/yinoodWc1vSxFsbhMc
bVFRPyD2PzVGtnH+7Uq3tDh/ifPE5NtQTY8in3evaCUZiEGPNtD117CoS6Yp7/pqxe6cj913SfN+
WIQ3U3SXlTNXwPpSGXp3Fzq1YIa5Aq8wxxSz0wFeQHvUB44GQoAiDRo4yt3qJSoB60fVDCctgKZp
uuMWaXy3y/KMmkDvne/XEqpA9edcsM+RVOlbTmjy5FbEgxxfXFvjXtaxCj+zfZyXXLcxD/i1s3Xg
zrjWjyw+2oRlQMcf2ipP0EvehsJvB7XGrNiWQl9ou5z34aJQ+neLiakZQWs0ng9oGqkYKs0/6Cmo
IuPeWvNOrmk0bra1xHKxhICuRZ1E/iaWko0NVDYbWsm+oemEqbc4xYa8BxbrxbZjkucozm30nKpp
+yeOShSWM3+4r7Lg2Z+DSaVrwZO0menAfM5pIzf9INOu9nJ+aEGCcoQw+3bizU3dEJi8Em8tx88s
dxs45GmFeOzXgZBUQsyiWsrqzL6lU4nks5xT9xVMI1bbXZ4E69nOJ068n2+2rwx0IPLF2y3KyXwH
LcJ9igYPbrS/etNPjOvu7oexNhr21rB1kCLP/Yp30fAA7WR+oyfQtTGBGiBnI4fQTtyGPa7HxCCa
uq0JnSqNbZt/V6NszDTPKjGiW3t1XWhVFkIY1Ate/M+nX7BxHAVpDmMnhhy1DTr5E4bwYMslnDzF
o+RyUjFMnneclAAP7NLp4zFEVArzDiUCjJPvntViLvdsj02QflY+Tp+kIRHTc/Q5EirswKmCnYOO
whfnd1yqmXSP1HZZjK4BlGlzBj16gf97rTp8S5jwy6xJ8cQs1ttgVbipp80wtCkgnnh9ddnsv5M+
DKcqWgg9HSTRqrF+tn2HguwJNaSiomrbn6gI49n4mfTmeLbpPHZtlbEiJZMGFqHxvh5QJYbck70E
9iis0fdPcPlQL+ilId35gyYhF9J9cEL2nNQE7au81icszIsMaig40lL7o3fPHMMLd2AcCkM9WulA
vQOeuqf5ACi+DU+tTTrOo2vVUzP0lh2aPi6pcze9VQrDdKdcGgSQXfT5a79XqoXW+UfxokHZgu6B
PBhEgUrpMO0nK6IHyn2YY4H1YPjXnGPC+OnDUwul6WIpeGitQu+6PNgKyPBao9eq1FLPkNxKEU+X
lB79dkOgvg5fIP1F5LzlK62HJQIiSP2RZvi1QaMyCICp4Gmiug1a+yfv4BEjFNwQkFB0QYDAqfw7
dPvZ4hZcrXJX5xKY4NnK2o3rHHS4Up0dS3SR596JHYD+sKARSHj8Hf+AXzrITMbtEL2Z4d8neqRW
dp6QFg9cdmwhkXxDvdA5pQGqlS+Ije+LTlOfs5xulcKSBa6waZ3A6zf/w6tmXPe7d1Gp4JjefvyV
OIES6zK814DMHiQujUZ5BdWyOugRS7725FpYj78d4lsEZYaurNuYfCwlyWo7WZBdoZtaSfuIIpaS
QZO31S3GJ+1/UxZKj+tT8zD83kiUHJpTOFb42xsqXUMXGJb8hqtn+eqOJFwU7mSnpM25jGGPJwzK
PzvVC/i3NDwhLe2fRN/5Clq6ZZatsbuStm+8306wkh+nrS887E7cLDYMU83dg2F3jLAuMzmrDGYd
FNKZwF1V5QH5VbMy0D93yGCQ6bm2P/RQrW8jjGYmCRxdOBOsJ5hMcsq2XCIBYRgERitKi3Sx6mxC
d3K68M9b+CeQ76v0QOZZODkZ0muxXOSQpbBIkMPQHkct31wWSj5+hD7ZG1wRtgdM2akYMA5V8xFi
qR+KQ8zsMujCVqbJkY70w1kXGFIoC+oBfMxb5XPUTL/Kdxp+i/YKqtxjf927VvFr2oEpzRcl3IoT
UIbI807T/k4kFy7x9mmk60nAFqZ4avwIx+D/vw+hLbrqJajJ12raByrPTOzETO0De9XdaJT1aAOD
ztyejP39X0FMghlVKG3rYu2Hxs/QqvUVBMflMBrrfJe6fooHKmEQiGN9VEPUQE0taavnnMlvQ2Zs
5+7T7ZxPEEkxpjtT/cfyKcX1to/7HBDlyCi+kErEfjyIRSMrdxcKb6FlQdosIAN1XDU2jj+AxtS4
uVreL5zNdbHFfWtE+ORe+U32x6k03rAn0IIXDnr03z2xfKDf6SL24GUAgjVV4gIgBNyFJF5RaOLK
O6IT16/olQmSVL8cTYl/Y7ZJLc6OjaL8e5mG5obZX5Lb3iSSEf35/S5ZPFuPDyfszjIFBBObJdN5
VDCtIdKD4JLDJ8dJB3a++My5kHhGZgnz3mbbVo6x6koLoKb6j8qXxNL5b/Wx/4k8+Xykm/cFX9IC
/gasEw831tct5ysOFfCGk4ggGHvlgoRkYlksOcfweqhlOC6/4JbNP5xalRcnx4I5IEPeQ9KqRigJ
FzzmDPn7i066hC6pHKuCxMkCY0+JahKFFpyElUeUDPwH4CZ5ATmlvhAuvQL/wzyOGQzqrhLxPFaA
x+rgJCz4yYtr9eEmgqT0Yp7PXfn2dTrDO9x2PklM9KDwUCRZxPmwBtQ6B8CxT/6KALOl/H5iuSro
bX3HdhdU8Pm7HJ2aTKs8Gd20SKrTLBOI/GbSqcUmp/4RMAi3mOwKbiM7ziA1jEQst/BVInnXA73e
lE6JTXKavpWK3+HniFK5NS/G6JtPym7kOwwzyOYXYTc9fa2ae1dZhahsZpZQUdUgcIYIcKe/mmmP
duHEEl7AaB9/mshVbEg9XG2c288WIhMtuolTD2Kg++F89tCcjaXHc5dUk2Ofd8KMj5ti3hziZuL1
lUZgi+VPx6TdZ2I0K8SeczKu6DmxmRb+O0yaM4X9cnDpRtfvYEUNN5NuzVKpEb+uhKPxtbGExx6S
KTsm+HG2uEss5oVHYTnEMeLjWj236tldyFnWk+XMfKDci5XrBSPS0kU1PSjixPwwMNZRgbjB93aW
jq15Mpd2TEf5iRMpZOKE1iCU68schRYwqf2idFOLYA0QyknVy+hNRG/WRw8MwYetT0WZG3bJmgGR
5UXJTRjHR6UT3tAKylVBUbtn5EwzsyX/Ng6vQsdOK2mp8eOC+AS0kAoqNr7LXzco7BIwHbnZvdGF
fRm+c5WqmpWQyPdLRRuH3X+WV5yc40XdVKZuA+coyTp2Jl91MaAOvewRih3eJZJMkdGtLREBxLSp
ZxQ/q9s87NNmub6XBYtdwS9DqzoEfjTa50CPnxzhJNuw0t0OjoV2V0aUNxVKirT8pcubFb9rGF7P
wOqQecSAgn0EtT+hwJz0/1OMm5D54ox86m7tISh8dpyglqTNEn6zx4nW8N08XXy7ErR9OTFNqvD0
lpdsf6ZaW34uCpiPN53iG4R+eTL7pEneoBCoav0XP1S5gicwYq0BapY1bV8ezNHk5MnICxgSqpQU
Oe/6W+u/MqiKSsrjSo3neSc89oCLMT4nFxeJ9TL2LVpiBPY7Ua9vcAT3Y7PaYP6XW9WFhKv3nXK0
3VEHLnQ/oA9WAHK7rG8FICot45EUG3tx31A53YCHgTroGpjbBV5tDki6Kl4pp2pABOUenXqg4mJw
JRq5nuaZqx1OzYvWKsnJIfo175vBC89Uw+3FLg3dsEHfLBX5FyU2VfTXJYe7Ft0aV56FzHJH0kFV
L7RmlBPt2dyGw14hV5PBfYWPXqsMKgdA7c/ZxXwplkvY4jqBk9SF1Yib6Nj0HT7yymUk2bCibeb0
QVKNERamNEeBfc9241YS61z/H45QaGIwCYWenxRNa2jPLVDjxSKy2JQNPbHqGuDADKneHHrKVIb4
nljhSqDSW/6x8huIUv6LffPsEncPQp5oDV3UvE+B73gTLmzv8FKTCHQV/SPaelZtQ5CWM4n7tGI3
9OFoExlQO9VN3bE2b1hraoAAXmeFBCTa8p/4Ly1/bkAiE/JTkY54aZCHS/WfBi2CREnk8EU1hiN0
+51pImZ1wHpQO2w5zSKgIgOZEmcvwGoUfaOuzlgW6HkcknUbCu16tl1V0xZLhXuVD3iJ3w4g+okH
V3kuEAlx3cfzYOOBHG40M0PECP34OldRKI298Zk7B23o0roavWf4PJqsexYLVqEuCBYC8TmryZuR
Pe5h+41JZ3B73N3hZ9ExZ2DNvqGMKpC7jnUASoLKvQ7BnuPVa/o69uVJOcVPqY586j1gyCjQNpvp
nFz89IG/IjOOXy6VD4ikXVGEdMa175VFnELK7MyDH80xEqshaWyopeUAEM56T+//zkIKlHvwQSd/
ldj8lzFvP3xy2JrntFbEesLRfbc+LFL/2wQXmzbOAvbhMoW59CLxf60eVgv4M/EKKwkxXuAFsUqt
n4+Nq6J3dsRY81IZWeHbVEJe9ymOifovBDuzhPgftVGH7D2fM6q5RM1/671Z8WPg22dOtVoUfm7p
pK4vaOxvFzuabYNJbffjI6HqN3GTjF5r2FFhDtYLmahutyYVepch5/Q5azyZF9PmVPOp7Pu1ABhc
4zlb2mVAL7Y9n2DFvu8xXk1rwAf9Y3dgufVaKQta5I+XLotU+06FRZmt4UXyB6pUYHdEOOzrsnnI
jrTjbtGYJMvhNIGOFgwte4tOW52K6hnB0QWoOc7Fg47KrMSnzD59x/88aiV9Q+/GxmZo7rCObf4I
d5hiOSRaObeN05WkGQ6KC9Olf6AlKV2+qX0pDMp7XhEGtDJukYJMFFjDzBCBUKdwUubIU4ykKKbJ
yXaCvrwVQur+Cv6vFub7ibMdv+/vjkLqmIdQ/oW55Xy3TC/UwdCxINmxvFxteO0N5NeU98RT2vqO
sCsp9G3n7M/fbzsDjmOCILFCiXhOKDaByMtAK8+BEcL1zVDhdIjNNlwGxreht+UEN/IKvK0lOGdK
IDKJxOhXzzCTO54pLXJBHLdWSe3ipYZCi/SyhtUaw1FXewny1eS9SnMxtB2F985FbJvzXhSQA798
/PVNeDEv4BNPenzj/UYSZbweqkJC9N9BAqvexDRw4IdMZPJeiyaVfCXBOWLI+n+jEdDP7fB7B1xG
UXsbBuNbQwIaWT2hMzTqac3Gs6ayINCKb6BtIsg++6wQmpQyC1CES/Ng+plpEgm4urJAvq/vuMkD
Pt097ELuRWFtx9v6FJ5BjWSgs7yL0aK1OLbaMislbqcyL01sakXrb30WuN0Qb97eZrP1uyJy9RGi
q7RSQi2gA9oTdZ0R9PZ0qdd9AJgsxduo5zl5OgQdTh/nfTm0dw8CPESGzBpMd2ANHcvLLZOROLq+
l5vt2hj8+HdHXUPorhuWbg0FrStApy/QB9nQOAL+9PJqxHoqrSAUnKDuBDh7EZXiw7aJQvxcIeWb
nWScmH7OQ13z7q2sDxPFVHylFGEBTzKtuIyZz62JbO2wTBVa3FfiMZBPH6kNyxMiFB6myf+aaJZY
NaiOhcqbUgzywup0H2t7iHk3Gz+qHCgHNkk5ZGqjOqUzgXZFVSLFVlg1pwf1R8/sy0HOTmbIEjBJ
j9Rf4lh919tUlNhWjQeB8ieKGqCkA2bTDEocwWOMOEjp+xbXCWCggwL+KElFE2/afueQTyjzYPwb
W0/6RSceThfI/+htXf9UdPQXwo5uE5jwNj5AfoI6WgBuYMlJ1arPaY/WvUtKCercqh7nh4f0XHRy
wvQtzxqoFwo2KQL9oPAsC24ZZfrp5s9N7cxVUvC/lwh2oNAGo7j4EVKY6SQ/S0jduskMAD8iutu5
vfiuZiGbh0m3pQGyIP+iSW0nuD/l3PP6yeup2n+4ZkNd6fGKwEkgo/ifgIL+pCfRDWkNZY87PNNl
Lxp01HT24tdA/kETCO8jNgxmuFbV9zIS/Owi7Vg1Zq7fIbxzpmvkWr7kbqnYHzIhOYca/0FeRw62
CsoO2OELZSDexHwmVUwHxl7YvUaWmKJyrbX+TA2lSiAq63p4teOeT31CKWNQN6AIHxMvOXFMXtyE
V4VvIl/8zxaMvOMlpL+XHCMs2Dm35vJLLCkX/LEEz3l7XbI+eDXGnrU95kL622xVrC9+ITkSOAZG
fJizYceKtNuIuFpYcmmxj5yQTJOmgQVFX5ppJEGnAaGSZvEMY/Ddd3sxuHvFSOGg0mZMde8oeK0O
AuOuCX5YmErZ18VgXYAjC4qu/a4KejBHF+2Kx6/EVrw6pEgTPQOF/TUkyz8PselZuJE/2Y/IuEhU
ndr+732t5RlEngVlE2O+dhZPdnPMBwH2x6oBQHD9CGNeAQzgvVBAXBMm/bZcnO68Q3MpFOiT506v
rUD3O6eCqyb+wxt3MwchUA235hTgIuVyhEM6f5hHWGxLdJDmxMyZGiMTbG44xoK1J4fyrwgiAcpW
/mAsMRRAL8fHld/+Gpyt8XVuKK294hV6oivyu//RRBvqOjze7V69can314zBNUMd7QyDlcfHXXNz
LkWw9W1BYCzzFf00SDQEb7ztNUiaKLlrBaKZWU8fRCwI57ctxgHjB98St59wCKLwR0ZUUMcH5vkT
GWohSnrvIl/AP4HeuiRrDuxWK+0kNcNbzCdX1xYfm/2/A0x3h73J1wI/PmE17mY5cP6nzSEXOGPL
I/s88n15gMJD13zSY3pXxxs6YyvNmRo4FLTVsSG+qvrIZIey4i6QhpQVOVcHO96RhEWQDRnjK1pJ
AbeLBlaWpTX+BLjb6e5FYsI3sPaXm9sjQVO85fW2/8wqyyLQY4kiSvSEuNmZLc45BAErf1jUBjjl
2Onwjs/bDxeELd6PF+M/kenLXyXJ8fAIqGqmA2n949LzMTyLL8+RJ+6ED252UF90eQ1xHbK4i39b
PozBRuLMjM1Id2Px59k5CzxsJMb59l1GBRiFxp2ArF3j4NidFERPIVTtRMCu0bZH6yms+oBNOkxi
ZKwS0TNIE/ksx3hkbgT8a6rYvD8dqp8stWIAEhKaT3wwKWIgMRefYrBssc8Sz7zL2TGi3atvRZ2e
O4PHcHVfoZ4bgMniIAaTkWl4oR7zCb85yaAHA1eKIzkxRkY3dSOKsFKBZCTwnPo3+5Stx96z4C3g
wEamGhLux88ExOJ1mzWvD9MKlmt+YEUB9yUiLqs4jcYguS2FhoNWsmRODjkpC3mQ7ldOND1nmOig
DYzKl2COTLKlzFJyfdVBt5ajvpj1MyFbzx+EQyLFiICRgOHzIlb/S92+Hxt0Cs+92kzsKdsqjgNZ
Kx1qeVN4mIr5ZgfeBl+5Jp8A7Vs/Sl4l0La7nnC+uAfQayK+EUHllkYi55UD4bK+3BXD8hHTvoPO
av8TIlGBzPmrnJLKgCXeerhF4jLdrleMvgJwEXEtCBtxAiheL2EAaStP9X1f6LE17f5mFkd1NR2d
anEvxgWHQRxMMdJ1QpxtEPqOfFWq4mTHFl1kSsr8o+lmj8xotmXL+7aupY1z3YVbjtBOrg27lCiL
VsdcKhL8KMuuoD2MdWidHecHsIENAwXG8WRXiHhDOspCPvJYXyKGO56tyJFGYrzR4wbZzC8R4mbD
bSXicq+nOgUIB1hqmYRqzIiS/N75JDC7Ayp3gG0ccSkyZ+lQBiFqoeiH9OeEsKUbj48PD7bw26o6
jrZqYsHY8BpPalGAKJdB0igZglWblzf6fzubqdB6xWKPa9m5bE9iY4Jnwi8skRPUUzisDCHMse+z
y2FRx9Np+ueIE9Zq6sKzvKGI4uNJiwoA7+m5xs81dvj5mV3GqUTBjrF4pI6TN/36Bg/pnpva8Xb1
5IJkx5pynoT6sndUihkpIPTkcweVL8ifYINv7+jkv49dpW1aTWdfNfm12hsMD9l7L+IDhKLC/vAy
T36mWSu0htGR0A+9Gqgirgo/acFOqqBzE8xnHTmi4ec5NJRFeqCnFxGQHZAdH5xJ07d+CCRr77WC
b7exm5fIImg3wFHlXCK7cin5mENd60SQebpRzTVNIl/hytOKeGBpYed5dKebadUyLhCp6AjSVkc7
VxMFe5/KLmOdofTOMIDOKYj7gqWWvIgpOGrdNXyJqU1T3gJop3uKfP0jcTETMagvSUVAehQDsSDF
kh3JiNFFdfBpJ87vjlzGMTt/5zfmXH3122eiaM1G6l+XxQs6pH906gMlQgmhh6lQiVr3YVy/KnH2
8XLOf4O/lJAeAZBtUE8sBPJbrnWB5+iQ6H4qgFN0aDhjoe7Gpe3VgglUxieFV+DYxFvmE6qOj61I
n5JP2Q0zD+SEOKTaUa/eBHkKoKHXevF9hrorrlNnaD3tO7cp0fJRozchW3TM1n1GfQyoIfNZrxBr
ERBliqCG+Rnk78ZSWo/ScM8SWg35G5cpzPzeVkSOyi3qogqqhMlpGROtMVjWEISxxrXsXT8bb11S
gQa0Y0vi3LqWu1k/y8Zr1aK1HSKautp8XVcUvQqSGhPAGO8HVNQ8VyTgETyhbNZADT24WdKN4hIP
PkUa+1gyVCfUDG9Hx8hoNH0nfi5v5IJi+1W828sBHBWcibM6gxAthEXp1yO9cbRzpuSg10ZxvPq2
9W61o89DGtjcYfHV4EWe+0PQqAE+dILf0E88HdWOIpLs7TD0S9sxMab2/fFySj8u6lOCgfdcuqdP
SqUbBhiu9oe1d+ACoOT9Ry3yOHnJJ6405db5TAMy9SWx9HE3Tc7eejGMDgbpu3Rp0MpXTIJlHXjB
7vB55l5SB8gvMFkRcnc/YQ0SrzmPgtGn5Qbt1D9IX6ZwFCAvRhP/B5yZpmAn3IWImTgmM8PkkrQm
4udIeg/R+iBl8jo5chwV7VGBuZ67zWiKtEkKTZFh1De7rOGGCSnqcs1Zt+dHRZcuUVJ+Y3SBHeqm
eILTYhwHRxdk6f2IiBxxft6dEe0cGNJqqpXFm2dhx7sv4EmYoh3EJ0GOwXgsZDZtCsoDk7DRApft
bS4QRPJV3/xELDtAvPxG0XDWy9TUywiXriypTfBF8Z0c8wyMwsgsAJEgboyPBgQ8WyCR9xDm+Is8
LFmzQzfyy+7glYd7OoWFJSVfiVSUiBlAKPNKxglLvHIuPN5BdujQ6i3odBJWAd7TSn60kJB0F90G
XHuMb9+o/NUMaiwk+KMXNE0/OaUqaQ1KwqzigYa7N7ki7+lYOEU1eg3D25venCF4IKPuhI0rVsmN
aQr01US9l9GoApPv+IZY2w/OHab5yVYqyu/Il8AaJ7EME55jJjHVjVaEJYvnzMcRJ4WkL5qwOIzA
t9rHwIQ0ogSbFpGY6mXYIFgvTVfIP1xVJ/OsO8AC4kr9jc/Mrqkezasb/BHkPvg7ddYTGU4bCiiX
0HFzsDLpv2obljE27CyT7uPno5Ep6dEwl0n6zIp9tjcaENzWtm3Rz7EpI6qNqJwDlU8SVs/Goylb
URgtpE5Lb/mwv9mZr1gSGGTlLZq7yNJdK0uPymjtsJ2HGyD03jmzdwJVcW60QrzOAfqZtntx3osp
Ln0qtp043qOUh7UboCOxOYYgkppgY2N3LxlsUTYVqp6lvU/5zp+jiCA5hxl38jYXAjG8X1+AC96M
r5SDDOhDvk64zT6e0Hdkj1n2IqBKa+k59vqxAbyaN+IAt+JsZ/bscmGqopNCmwxJr8Z+f8EipiGl
nzC8Uprl7xOtwfw4GZa3LZ1TSeQI/AblidkwoD3wCn8VVjYd+agXnmXF5vyTqgkd9DlQisQ+beWR
GZvlaulahuNDZs72PjysNTlQrHMlZxlwDYbejlWcP4ptSdeE3QKkxSrv1ZMOBQhObcXKq80Q/7eE
HQ+7PbGvMbRAG7sotF4H6psq908F+e1SpAIX2s943XPUAKfrTzwxaaajY1q3vUPlobhYRPllqXbw
ioAdqC8sColt1jwhitR+LB1bymKGs2ZLB9CzaqckqQpa8M7V2bYMYQgQeRrC2SnkaYXTAGru+rU/
EiO43L6giJzAwTL7gpy6hxZ7O/Kqa9R09E0wid6juqLexA4CiifU99XQ4t4jMRrJdaJIfgwwT4kV
5DI2cOBWTWLMwAl7noIeib0V572pjlbTZKGhdKvKF+mcnSDgd/sXR+hdaluugiqKoCOOISK4cr2+
1YLPYXQHc8q5lmyfnn3eHyehGgckif5VBGP/I+Y6sQA6KlmtccV3vj8FQvMLaBWeHSk5fesw+4PQ
+aQPQAHlFeTwge9mjgO6Tk+RolQPTsYUAEQwnKwIu/UhhR1PnOtUXytS1Oek+X+WerIa+1w1dawr
9pexHngibPJwvCvh5M651uXBMmIg4UhIG2XPYALIIQm7PWZOdvE674YxSHAQ05aI5f4c7IqlGpWx
9UIiLO+1SKq4U9juPb+3xnXjw2EmR+8hmiWgHLabwf72JGnufU6ckkWiTwYujfrmpnFZ2MzJZkh+
F5SsEFYzTY1CFVZ5on2pgvaRHfIxYOocVTxT2J/c94b5oKaN+Gxp58M7377TFW9N4YrZU5Q1jhUq
O+cssB4HZUIsRj+0gV5TFOkAmDbk5rft/UR5amTEzyiukNaAo2wYD/kb3FZroKGGjDdGUJEccXGX
avakUOiJZvocHUVWv/2xEpdF1r9fDU1+HqmuuaD7gVtlEXmRdHj/8/+mMtUBpBjlmPCvLAxGaLr6
5srugH20stOzzLJ5Cb+SUozqyCOsDuHhYctlNSTXyOQuag+dTzwNEN9ICtlYDOdGzTmjtdeVc0LH
lo57d2Ro8+RvxBaLGSsBAqxCBFyC93U+seN/OC03qb8mSSGMWaENuUdG9DHWnpG0iy233B0ZUfwi
wX2Lfa4ud20Hrgpi97OuHWWqgyLmlI3zSfc7iKzepqfvZxkv8GiqJn5/eFZQYN5q1a5PlRkE+dgi
EIXfxlTmxcWO8LtwGKhrrVb9GpiQoV5PA2Xzxj0E+yWptMACqFIOmuueKPBDjDlnuJxzwm7tQuBS
49dk2E2hG7ETLSz9n8s+I/fC2TsyHCeo0FZRREmK+rSjeQaQxNhKY/rEM9bR4Y0Nmqgt1SrL8jrT
ImRKyXhUePO3iqgX0Me6ft614ASUMNcd5ydzxYb+GCAfAcaP0Cp6/25C7XQ1mZQQ5XkZbz6QMC7f
LpGxAqmoZaBj56JE/ACTZZOkMDzGRq4ycLmk69toaY8xW0hPYKBe2+ObLKX3dZoG3yn3pg9r5Mm1
LPR8R5rm++cGIde8+/+chBbYpidRV79R3aeekICSvmMY86kzDPeJaNoSo/iuK4QFdNGCSH9R+0Wv
ZDmhn5ESIN+x01dtj5YQF7PprnusDiyriBrzwkg2Qz52BsZzP166aLkfOGCgv19DPfOp/bGU8ts0
BOcAG72ioMUaeu4K9UOPBvKNfUh85zPRDYjz+exWd7nVdPfQ+AxACDdpVSc6GV0eL9Xagajp0U7Y
/7a5Ach2vJrFN50KM+oPMJOvPp0Z9U7jBxc0QyRmSdTMAdqjDS5DeNHi1F/edLIBQz0Dofb0HMKa
oJ1fQ3KfOW/JHwaljqiTi8zWgd9xXUYOdCL7M0XYL7OdMawHApUhOgSz1ucXEp/lRNwzc5ooTdM2
6KkC4JM1iGlCL4n36m/ErV/fCUEdBX3lhcVZc4ZEWbDkb9HwG02BrmFw5MM7suo8H7+qDYQ6BLqR
66ntmyHRFRTuMLjh6I9yvenllpjkbRy6BXxPCqPWftrvWKmQnfogwtcs+1DVxkB6gglVJO9rA2uh
WLT5WMGlfImf/yU6ZpVniZwpJxV5iZ/F58E/N5g1zup7rJnj4b8TDaEzYEfVF3KuY9r2QuFAMLM1
mXv0RHtHOnRq1jkJSHe0oAkDOY2UN76PGW2Sv3+g6t9H50pI5Q89wvCwW8B8urmKjcOAE+Rkjnae
qVxeyxSVW+b2qYohPrBzoX9IaZwhQGVuwo4KaqwJcZPhui+obrHnVuvNE1hcbowKKQeQcnB6dnC6
RbHTwTi9wpW9p0/HUnCu1VUxsbMCBJPTFvbYdO2pK2iksOeKyhMtinPB0jPdSd9CuU38l9vBfZlh
yibGcSwO0NapCat2+9DJiaBzWFlVNPvjSrhbG5mDdNdKgZiZIDVwJ0yB6gVvz+9CJWIwlp44xPDI
OZXRPpce9zA4uTSWW7Ob5f9fqlfJfvNRCNm2fI0wJpS35tTZ8h/9S3TAFnP1FH42GAvRgbKkaN2A
WrWhj2KdlTEIpOMvkfaBgQExEUGOXFwpFDInAJRPRtbpK8YW+BH8JZYq07NiO7wMSJGvi7PAZRfa
tR7seeZ5a+WH1u7ddj7aR01HlUGRQfs2pA9+dnNszOpWWcQI3TNoQP6azepUp6Xo5AqHYgkiG0d6
6MurSUzdlrpa84oLsTqv/ZmseUoMKxGZmn400EvuD036Uf+V4Xcu2WgxQWw6HkGUe3EO5a7GK/Dl
7dSbuA7O2fXjSzU5gByNi2P/Oyci7n2QJDzD+yHL5/5lBdpNPWRtc+qU4gIF64gf/dDVQ0FjI+qf
ku+wejlEnNjdHaQfd4plpwT9i0UslYXiEXoNYOvhAnIEGoTGYDUz54UAMPWQ5zeRLF860y5Xf82e
7/WMXptuOuPlDyWP7oFxyulEaTRlP1hSXhvaSBbmC7dCpLNI/xXuIUJE5hx1Grsv3AP/LK9UqOB5
RchbURD2a9Tmg8loDcl2M2c5/JULeHqYqXHzmMwnevyFnrlm6cdVwC4FWKoxh+Lf+pb7kuPkd27z
pFOV8bnmeQB4ho37nQnB/eDUfDofGrFg4QKFTudGwJOfiGRmYBiH62ofjWJZR+j2TmCRoNvDcWmQ
TbN5uHXJRF6/2exZQHuqEBN6S4rh5EhtbC6XjhfBNDz3oOS+lgU3hlkmnV9guFlaJ3mf4xRf5200
0GXygGmJsQKXbKfuLaO/9nqe5gzJykZ0Y9LUDMKi9IWvEdOAdJa2UHQJpH1fN2bz0xEiAp+wApW1
8jldTorNaJ31jBvxg5RWlxifrKhhAKGz2Bo09u4iEjweR6a4gRr31SItdrgltThodIKFjA0fbGuZ
9wbXQpeOIDWi1WErrAlKk0vBssBlAkxK2aJQ7ONl6BQ6BnzpZ0wpbEnWnaaykB6NkwtxjlOS1HLz
7cmhsaNX/yXkbNwu8lKOjskGJBus3SLiXhLnxqq01MRZLt2KTbPpwdcFVVN9eLtm1eM2AfzhiAEp
3JoDlML4284VJb1h25VCSMer1iSDld2zV4MxWcKbkGU1hOH3qnftMrrkP4APUTSgtYGI7yMQ2eiz
WLYvUPvz9CZARD4iJSAPRhJRxoZgN1WoZrRvXAWrx57zUrIp/2JAASYqZiSXyWVfT/n+amfNPWoe
5moirsg/FLFI4G3mH2QowJHGpPeZxMoYeq3XJJinayCSy9Z72y0bE164VobUrmqxwsgXL2lz/6Kd
FaEoM1GQ2jmDE2qoAWD32yETA/ToNKuV0nbAhnHX9l5Q1uZzMlqUiPfDgEWvPzLOn5LWthSycoVD
JBMX5n7csG0nmusvl8gTCEwJeMq1u2teb09E2XAJUTu756TPbUGI40419Doppo8UKL8kp/jG8xYf
a8fN4yDKTi6FKMtNrDwG3+eENx3nRkznDArX6hbmMZnZA6VXPaOKicgQsUSHx/b9He9+hCOsixmE
KYIiWFJpi7saJ/pLEiA55IZLnY78QDCINYfkYcKNqAxOq5dsS5Ox5Fao1Q8tmDCeQh8xMKprToqF
95uehLQRSbli72Vko9xI3uhZnl8eZ06BS17RMBqOZpIky4t/GUgps3AA4iBGrEVIOXHkcMo0GwkX
1+H8lVT+0sxy3sou0MjhbN7/LnaOjPA6OtQjD+s2n/8x0+FJ0sFBx+UztuHljqt0vfJoA53uwCaz
zPDUhjNUav9A+HgNmUEvXjyXKu9ZAXWO9x8bR5RpU6BWArpLtF4rA1xMUi2bGy6b4+mpn6Y79vWo
8/z6Y2FxXRc+wN/vxgmUAvWdbmm0UO0hnQn3OikHGY8yvi2ovhsx6uA9dZeeKJuQ/TnF1WGxMBje
FmfTwB7me6Glz1C+IHuwfNIP8th5xv3VBm9VYupajczaartl8+JBY5lAzyoiAnp1if2zlJqXWJ+J
UjBFRLkmAhQ3FpbP4Dgfg0s5F2rLgBU6X/T5qEmgbJ7BMCcs16C+m/m/Xgp2XN0QJtDt8TvvZ6FK
E/CH4qxWC/9LLJEk2FmCJSGAfwnleOjNs5nsRZN0TeJRl9oWmIWk0FW2VImjC+yXolCxONE9ZNYv
8OuhCIl5r0pVnxcExCAu7w7QhOIayHAammYzCmhB3qJz2z+1tXAVlnPyhQ26txREgBtfHurUnxz3
vEG4ZiLdlJim2bg4fi7BxBvM4Vnl5lkPCLxAdFlTBv/ssQ916jqUIJNTiCRvUjL7xFn+a4CcsVXG
Q0YxWDrXhKGK+9orfV3V6yMcgu1WhzfaMqXaM7qf6ztpUlw7Onh78PlI42bGdsyqGo1EoEeNI5zS
T+l88BTxTNv9rNBJUljtvMGGZ0XMVdpdUW28Ink/o8xrLET+E8lZxNvRBydm35fg92aX6azXjGMk
ZTkLWRBYGk/opLImohpjnxqagimirfyx5+JLGFZ/BpwRU1x/hjoNnlkEbs1+VcqHxmqdV8r6wU4p
MHP/tzZz0vrupboZZ4kWnW0CqSJW5j1xMajcWGMr3fwKh0/ajjo41XmNRN5B6vDhBXPQ6zueVBhc
jUS9IUxAPz64bbeIPat8XSv9fFnCxW3Dy6tLj5XClJ0TJqDVnG7xY30Hk0whXLZ40XXUwtVuz946
Dtb5dlZmo2jSdmgNGVUCInfZLOM6kNPGkxtXRnkhs1oxqCO+stlQ0ogQQZLRihbkshHScATjfJl6
g6DeBPoklwa3EaWrxlrht0BlzQsgaXLETZlTd99Pycg+cFUsy0lvsU7QkraARLwp/zTxUiJHdlP2
Dq7M/L6LbkF+eNAbLbZlF/+N4mTkw56wCTLNC5T01Nh4JCsC8MEATYtsoNt4k/1iZQ9cCFCLYSFe
TyZEfa3bq8kyGEbn2yzCTAQrLLvDoZPNn5VBEDIsN3bQWcZst7LF8qeKd6w7S0QfUz11Qbqvsy0G
fSbDKWRuYfYg9I05dRtPPTOIGK7QkOxNLB3LUal1t3wTFAvcTN0Fzl8mgNj1500eJmkk2UtaziMi
WYdW0DO24zzYB2dUXA9yBt98bHY+RmYBz5ePIocfNT5xdNamQHTQCM6LL26CGZz+qitERtSlC8Iz
2W5ZmbM+838rmxd91/wBSaOfBmPMbGibZw0pVszN+km28yN4pW9aXJ4QdGJaIUgzhl4YeWaz+JE9
2rVwvFLsLmFr4rRVEU1xxkMjbj5JNXbJ/x/yQm0XNnf8rqntKbV8ElauvCeXtyBkTPPlGnnl1LBh
ZOiSMJcEik7aKnwmPsf6DNTd9w86w5yZcawTA4vtLDWlfEjrFUKlSaehLyHhyMS8PoZO2uITSYXC
oONnuNGh65a2GXBSAuGiBbmp1XANfyR0DPcf6ZuKKSeO400h6nnwvy8Jq2xKe/IY8iv553W6VBQO
3K9yZKYItWTIwp3i9/Kq4qW8f3Wsz7r0MwuTuKtOklD07eLNlWGTaT2sxiOtsRm8mcfZpuIXyVP7
0t3lgp+konw6UWRYRTP6+4qHDgFOjFwz2q7ZZX5FsB8QlWknGnY7Y5wMlVK5FO/jqS/FKLpVX2gx
cHXyCKqJNXMnqS/jzSLHRz4uci466yo2lcJztbxOYm5G56b69yNhdzTcNEOMnexwm20czeSos2Hf
2kTaWhc7Usz1wJtQSj57tZFen8y7xauNg4Y7MqzYrBOXhzWQATqis/hRXkFIZtfqpURrmw7bLBZD
k23j2WeoqoOMshjudLPUhGVyXANwevH26pKghdb/50UL+QTEZAGvSev7m7lkeGb0wcQPrV/V6xco
0+g3C0w6nsmF7iO3OuQGJgg4/9s3TDXR6xr+8578s/bxGNyxYNF8MzaxLQjC7P4fLiITNVcfhpAs
tuqLYQ8R2vsM+5Jp2UnkyGSstMXAz063ux8FFcysrQ+2iqv07Mw9GvKD+UULTTKCqFsXzcS1m4Wp
kI2kvp/GIwgQ69URdy6qfkQiA7/roKgJ/XTpkxtWgVdDDPSB6T50rveST1WksvDPhUkx/V630GNF
6ynjzV8W1RcsQEymuk0Xll61oS5y9g4xCuPYLMqFbYgo6adtlSkjGCxEZg102dbmh5w6VzflEc/w
0iDjR9B6xAy5LSjFbLlgyORU93dlAyymzGY0TC8w0Q5WkKwhLTyy5C5qu0iahZRkRBFPOL0F7P0o
4Z1BmCjkm6vrlkP+Uwxy2dJwWdWE7fleX/ByxTu8NwWAhxhOstsofPSR6LfZYDqJ49FQg37UBh+5
sfOds+ucxHxRAPUK9zJjX+gCx+zngCx8aCcXoLee7FHvkIZkCvLwTKUyJIwyJtiKLY0UslJhXDdH
oVC+tRnBDz6Aq7OpDph1avYXi272L5X4iYJrkuels08VVB2lXpXaWsZgE0YIP0bfz/3hizsb/RRp
sPk53kVyI5eKCikzGBjfhhXl+UD0bm97q0VamaW/TZy31bFjVzzfO5TXUYWT4feO0nsNbZpC3auK
j+IU8CxoU3zh4fdUblyZraXn/5FKNhjIFO4Xxcj9KYGL5lduVyt9tK2CK/lpRGoqv42BmYEP8BpI
SFtoEheB8YCPwIy8vUMhp9OjaX9XMBbqBnyB0nGWf6o+xuscywDt0wbKPkskSIdXr9lb9CGo4VSG
y6wL9GYPK0Hx5MbPl9m2p0UlwRrpqu9hQ4AUm5KKQfMxxse/tEY4EqgqaG1OcgBqEpEhdkJeDLUW
V1t+ksxS3Ur1U55oL7YRv48FNOxIKfn7s0vhEScWcHqT9fmbkQZF7rnA5ik6BVUhwOdKWUDC65Ut
fJNDfCsJDKwvoLDqEy+MdVIjmZsCFSrwglakjIvFk7zBawOI5djPl5eJDCYKYEQxWvmnnkvgR3ZQ
/N9YGcNw5AhXzeFt/eEhK9dSZvKIH0EmuJTeuLNFISJwguDiSlkJqm+yUw24ETjsmbsIKB2VsoCH
zwIF0XYQqq2ZxfP4NJbq82BXBiOAyMqVIWD0dmU6B/JpUhduXxqEN1S7qT/acsci5j8F5FSJWsLw
0D4/htGy4puRaPBhQxYdZq2maxzcDwDykR0A8jHZoMXhAjEW0bVdeZm+zZ44/5Hl0S2gvkIR2yaq
U97SmDk5h94hGbJ2dAEh6ArTxJFgvCZI4KJFaRNZx4NTsjCdTgglKQwoy3I5pBQMMUWp2xxZrszb
t/Q7FtUvcmJrmo1rrnTC1hYe7CtfflkwdP9dYW2KeGiPZRtaK590JGuO2CajBy8ztqewqPnyOQ2b
s79eDKKVo0BINjFzu8D9k2jQUvmOhe9PCtZ3egrLI2teWLQyW0Iz0wSsj6lnbtgStrJHFj3ESeep
P2YmqCikPvjF4lKBUtMZOpvm2I3B09aDXF8WXOHZYr0l6WWDWd5KE7XQsQIRLa0c+tW5ZySG4z5v
3lOlsTM2Yk2Wm+iPtMTLTI20XXRS2164KhsaX017SkAnCTER8OvtGf0Dj/MJ/fSSbStMzMPDS6oe
r5U5YkWncIqgCGcOryI6ql8ZHc6eSo/btuFEalOKGU5eZpaGseq6sbYi7AdaMustm4zTKkvQHIz3
MbixcIT4D21tqCBq7/+p33OXt3ZRbO9Ts+eYkUj0ELGuKvc7REGh2z8Hisdm/Gql9zJjFtDgumn+
B+0gTDAfW5YPUNhSkYHF+4UcZKeDDpXm4YqDPTFRxund1skvB8aaVwRLJvvRl3Ie5krPYaomskaC
D9FSomgr9ZGVa9jWSXr9y/0GVmsitkreTNZA+O59+y1aYXgOPuOiH1C5RxCkM+em9Q8p4SN/ABD0
cOPOmOfE1QHajFhQKfUbNbvhMY0xkPoDzWWT45MCd6AFQA1n9hruPTkTqY5RfhaDKonEDGZM5lHN
La257UbRZWyRYeTU/ZRGO8lg21Yac9PWsTo7ePmh1opwuJYIK1JtLXjBIJzlizYJ7sJ32xfqKUtM
g/1gCd5PO3n5RfFm9Ivx9OYHhdiX4OYP8cCOUy+3+83S99VczEKJbrRtdORYG9sy+CLvOnD2fCo0
JSpB/MnIJUkLqWa1kiuPBBUmeAIDjdbCp1bKBVQaXtv6ZPueD2pYzR3VTb8aJb0h4Ll7VMwylRW+
Og2XqYWACfws1K+PRowMl2Ira8aSmI0+Dy5RKgIZjUZrh6jRK0kJyDf/qur9/TNx8jJWJQV4RR7C
GtjnglJbTQVKJ6k2R0Yq/6rMkQIAQYx5uYdmJxqza9OI+bY7soUfB5qBGXQNuevutxvCVaRSg1IO
zimFHvVsi0XJJ1Y4DwPJguRgXtetfugvxeOX7FLAnAdWAPxSbs6wvZlXi6kvzxG7hGqBahMrURmL
tWI90oJv1JIbK2ytOznX4jJ0sU/Bs6QgdQ7B3u0pa5kELEXNTBouvSVtG3Kqmusr+p2HjqBjYFav
Iv8dig02RideyRvnRCiav9hcHLi/cR4Nr/2Uxblklleh1S2Rq4pCVrEdzwsg6EMzhJGyyH3HtL3Q
79aKq3bI2LoQC404owtiaLmte0MYZwblsBxGH0J58cuKJ8Ikhh5bI++oSmNc1fnX6Wb7D5dB+xiO
/SlpmjEfXXkoAmkYvw8vjcPCSIsn+Ra/0CTqEZShkATKqMLAdoSwy7VZ0mjDjJfdg7VsyjbKEHtS
AT+bdstj+jLwoHPZl+20W5OdLZDknq3+twuyd0iZlR7BhIrNtzPFpafQWDObrR0sO/edm9unQUxO
AAQoy/ibPGqcp70321RSRmhc1yNom3QJ3TaVqh5XCQ7vK9Iq4N3JLc1TUUAMRx9cMJb8N0LX0BBJ
s1BKXRY2b7WCyDbdas7OBkY92/cKa1R/5DfVSfe5bU2QiLF0mPmqc0Vf2ewI55rlLJZvEQMOEKWp
+jme834THeXJAfPjcteSbEMe/wm/k/cVK7vNnGIPQK/Oyat/udpiP+jedemWgAgX+GCyqTVlX3lY
yQyBLdeYAfdZvu///NkxtYKsRx7v9ShMNUfvTvy53/WqnEVrg6ieIEAZAR1+LyhmXSk+BhwcYHD+
au+GZ1rAl8lH/OJ0JefcoCoXsWEkip+nXixmu75UjbKOj7sTiRh2L5kF10l5m1msAPen6v4Deeki
U1kaEFv4ZuYDoz7yUJxdPXKwMzLnoukbRb5VijH8lobBXfdH27Zz+eFiErPOAk+48sSZzpkYtHTE
YogagH3vzzF3G5uI5jXQQ53giwwSsDN1nZsZ99TWwTa4l1Uo6LjVy6y20eZib2PEZyoVcGJBlR8n
/053zU/PkGWtLDXEAoUoV4FMrW3jSmFq83yd9+IQS22CL1sVvPtem1oh44AfU/e9jBz+GHE7IBWl
C7Eh9T4cvs3gMlBTcBUvQSZjw8k0mjIh5/WBhnx51p7SwvWr3dEe74kKJ8xA8YBTaNliWjo8xCUy
X6lUAOzQS9kEj45dfXoXexpBzIVHYkWi6j2++4YVg9sGmT9c3lngkymxAfdN8DwVnAlvpWRD6zTE
1CNMeMDtGHaiFfsGwVjLMOk9BZT+yuKCAuLpDWQJgK/3+lPVG4s05wgl72/v6R6wXOvhtAXtkZEr
g4P2ha+ZB32yRvqdjBi571ZXCmcgCf3BCRuJSAyYtpAygqkX/tX0KhR3VwF6050Rtz35rKwxauww
/BBeq+vKOU+6Y+H6MqM6KvnaZe1nY007jKIgx5tXiFEQ/QCh/kihlzDk7CxwwjW1E14iq9ZvQaPp
cUdGgICIGDxmU+S/UAx4EZpri02Q3MTxxKSQg3d5SRMhMQU4TiH2zKc0g+1uukM+YsfhuICX0aGO
fpGUEbOZhM2XwLFrdMWQkrQdmt8zfq0Ff3c4g6nRHsJ1wcFUGCTdmblCI6BSFBMDqGPnyNl6PO/v
SdbTLGONllaQzJa8uGBdPcweZFczxKGKOisULqyV8lNAmAV6IOqM78CYUK8FSfpp5LbYeuLGs+Ou
jp6UwARGddyLe6pccouw+caf+HVGvsMHZYplB9a4H0MW64BP5fJNLMSO81D3WKpa1o/JGpuaS0fd
Q8jqaCPLlkKdEBwY40Sy9UJjuVDStH+ftsChXA7CT+gqOEGxY9+mbcXAf9BGUPWnWKmL0/Pv9Uno
NVcyqW8fHbrB0WyZljcmr9B85vAcdtDBLocfF8S1A0IHo2BCp5X6Or5xeSZgRf/pthYILQor2GZJ
KF18nEEpVWL2RnOA+TzWw9lOyEZoQKdO2T6y8arbfiAi/X2Drd6/1HbTBnz4m1r3w4HX5ZiJgVXQ
1VUw1/xVOjzQ3ie3cpAz2XwdjMa0tLR0Y8xEfOONHDwCt/AOjo6ke8O4o/kettpSWs2NF1LydvcF
9RPVkGWwmO6wWJoKsFYxOEMU+WuPfa4JigdsmEyGg9V5/wmpgMVo96qdmqshPMLgSxYzT62iFrdv
k/RjBgVmWJ51Bh3P0PrMSEFE1hYXsfq+iOJ1MKXR7j3R/aE/1DIlNvNLxDOG6ovtkWCGFMc6brcD
MckZBXC7oq35RJkr3BxLRP9Rcn3YephnIcyt5Df5I8HgNsmkKAPwPuVz7wfXTHGClQ768Y9/17UX
lNYMoHoQ9BErowDk0mwPNjrQb2pbA2Q6X2cVR2ik/1WXfR+YNqVXhwPgICQ26mZdPDTjFaXeLBT8
p+TLWdfvkSO7dgPN/Gt46YnarZpyJFpyNmXKxa2d9hBB7wFzeIQhChQnMpHcZ/6y0aLgyFcOnUoI
rPNbYd+vQ+RATuSbX2opDrNf8lq5Sx09VeOO8E9TWZ7D1W7SqKXIA1O/nUvRh0d0KZ3WJNmCXGK4
G5zKyRbQmAvPIWxnSBL4yVIwXZXvsAxrdTJ1AOp5iUNa1bZR19P2egQWScLKVYTklnja0auLhAgC
bxVzFTqJHJrTXPWKmk8BVehzN9sgZMlUkher7dFC6Pgl3t13VLLISHVdfiqKBsFUpQF8qJfdgfkV
0WrLkI0tn5dv24Hhpg3nCKLc36eN1p6BlFerCgFhg68dyVVDlLnLTPkFRUA+CAZpyB+dIzPs8aqJ
JKnp70CbW90akdEJrjkyv17c0221PAV1B4UK84OjvdcZQ98Eh0H1/HjgyrUmj30/p6iBTjmBjXdX
aNo37jJ0SvS3tWDkfsUtpTXnQaUSFuv0XES03YzJ+Fsk6RYoQC+gMf4szKe8bi7EleQDryz0uj94
frxd5xa7IUkcsnMLm1UIWKmjgDJXeb1E0e2ftECev+Dv+KFPpWwVoooxoC7xzF9HKUDKEhW2Jsk1
moZO0zOmCFFgU2Ldwp+1jfemxA38uWJH4JmJoxshFyup86aoHuSug9zbmTHQEthG9I1SGPoiYB3i
NNETalZ2YPPccZz7oT9KC0N3dmrjKLKADzSAQlnfOWBtQBu/fHi7K8Q0gbrMDQ9c2GVj84Lr/kLu
aYraKL8HG/ArHCnbUVzbGJzcFIA0zO2+pgGOWdyrDjoBO9ObkE80CLPCbaYyYGxNM8lG/snWsVBC
JY6UZ6ycCJ1WaFVF/ykuRsD7DQv9Gzl6ZnYT06TSfbFdxN6fUbB1Q65pwx7Mf4P5Y5lPiajhlStu
jD09TPpV29CyQWrjNGhATCxL6pY0JL7amS1B/ptBUdubbTI+kZTDdxj3rk0FYJnBjdJzkkj1X/iX
3jRIFPWR8TgW6CL8Zh91jGzddlP9kaeo9gzlTOYjqH9UDsE88gsUTWk5+bVQa60om4nElEldlnHS
DdKTtG1LTm0p3YMjDvWBAMjB5ej01KxE++4csxYYYBSfD0R4kFjVQDWou3y4O5et9Rz8MFkg0zKz
G5ftjW7+rc8wnQ3d32fjgJKF8aOFFNsL8kCWC8R1gqxKjHFl0YdEwYkbweAxqak+z6vA0F41SZyM
kInha+M6Cl8jxoikeOsmzs3I4Vug9w13VlHN+HUvcX+ncWjHk0Sy5ESGAhWpJULX5rRcEha/2Cwr
wZFPllVVCo/J5XjxRoyftpkHx8oiGtv9rBTJxm3D9dkfXd1KEqoYkUvRz+/bW5k4d5Wa3zzpylJu
r1Ygs9MdmIWbespDbptdb98Gz3wDphQSZkBWdN+EwI/4JOP/xr1/3hcuVYs8Gk/jV9kx3Y7xzE+D
hZp1C4c/9yBY/SyKxyB6kfvLRtop39H+KSiLLh+Ki/5JPxzc0G9QzsRD4Yzlp9Bf8/5K9xT2Rd9l
ZemX9J1lPd+2F//FZeVF2ehItOmhhBDQVTKpXBH91Lb3XFsxbX0Eq56Ha5MFjuF7jgLPzkH/Lgif
eCIt69DW9LlfMySyqVYTBk35nPo/0G1+xF5JvN8nWnWTrCn0ZltQRpq5PiE3mXwlTnvgy/UE5qxC
g04huDihv91iks5nP51qrOTkQyYN1Ej92UUj0oRP0q2TMsZGJzgn4uEE1x4AZXbUilXTKO7xLpjP
nPnm7dxVsfNVL0rxiGqETFtVowgAWswWxFrpd3Wbjr4rwqxjN74aDHpxJ/wZD9Bdxs/ASEBCDV9Z
0smzhSfGnXgF7LFHVgDzr6YkZ3kg2L3m46k24AYV+KoDYOubIbsUpzVG9zbqKlcJMc9F+QI3jE2P
oe/i1xXELh35BAUZLAyduS7afKSuHQkOuhCmVjNYjB7o41kM+xrT3hEoQWSJXuXHd1zaklkqt/s6
TvfaK/MHCBm/TJToFXpe52m1WGA67WY1GC0yo/H4TXQ5tOb6/jjR5/k70CTz9celb781rX4kZyJ2
0MCooS9pLk5O4y8h3vyo2ndGiJvpGak+Chi7oFxN1Zmr9D/3MeAUUzX5ymHi1e2jeVy+QURhUoWs
jjXfzrWEuh82bXPCPeX3+mD8p0nbdKV/8e++ojNP/GUbLGMyEkCoOUoT28TVVTCZcQM9Ck0CT2Kp
SncK3dt63bjaQyfylNAYDNJl1wCMcvYRgF68+4w7LTQFquvffZ4/7BNTY5YQ0jUjK7d73bEe9xli
3QQn4RjSyO1sY/4F+xDPGXkR++epj0ahcYRDoeukc7kTNZkzlcFWSpMjvv1OMLCuMYSr95Epv07I
S6kmXrkrsnWquuNg2mkCAyzhyMUOQ+u+DZmXVrmCi8ptsdYldQ+18J1IYNGLx2FCbsN7Ft37D7e+
JFWZL62uOurndKeXRncrzWy1JpYOWDBgSfrUoAVheaBY60rX9/3eiE7rkexRMdTjZdJ0kmGuU8dv
ZJ9WIOrX6JE7cw2nsKUvDwfpq5rog6fM625g4WMtcXOxPV1LFnxc5TlnCtqbzu7gDhBOHKHbP94U
FJ6XeXdOPyRS3QApJshO6asUjXOG82PNlEciSuH6MgfDiHq0KrpZlvyIjtqyYRp2VUKtrV9oIvPB
zaiZlZqnjEprMygZ1Dapgo5jSy+q3W/JOABd+XWPBayNsDahUMVsLH4xB4+AsD48yUtkJmY9iwfJ
G8/b41VXObZxWYYd93KgVqthm+kUuPoSxjV+NwDrFFDvB85xHofjXc5kckqUI0PKkv1/CPHi0+Md
zWMNIbZergHvu+83W7oq0p0QtFZu38MDXjWo0DRV0JpOG28X3iXe5Ftj7/DPyhkCrZ7s284f+7ql
uA3kQvLx1vfUPQ8+UJyYEqlZqPXHDcu8MqjnjnkI0xm0168qipjfHDjbnEZMsruxTwSLhFmvEEMn
XjUkSU99iJKn5P9XuGM3scmCE7TZ2tMpGP20uoDy0YrZQcKEjKhrwaynqlb9eWdtkvSTuM8WhWOc
6wgDLQUxpr2AQpR0gOO/Q4T2qKCDsH3vNeo2lHqJqB/Z5FBeGblIX06gBPw0rX5cqTl7w1dXpDvs
T5SGJl/ps1SkeqjZ3J5U2gXQ78/5IFYaominbTe1ssWQqAhLbQyaSZ1WXamHg81ruJl10gNoKCwz
fGLtawfsqkUqFO3oVh/NbpHGways06dBBh/G5PJxRFcn6qlHMcs4PYjU+45rZhv7tuH0Kj8Z2/XD
mBUM2STeQgTcn/4EfUUldBdcKyXoih+f57wRae06g7UerfdmU6ArjRuD8ozM5zltTV5gnUUd73TE
VCX5MpRofL9rZoOwUoglGNsyBVZVEdXcYJOSz0pZ0nS4HchUtVul8reME3Zr/hR8uRRKOhSlhHnw
OeR5aL6/QErCESQSUhndP1sMXz2bT299Yfsw0qvWlaw76EuoP80vJFR9rKRVsgA73WAy6iyI+iW+
6/NaddmzJJVvN2cX/CxCzdaR/gA51wl16p0yZAutovolXkjbgY5+9o2em5rfIriNP1g96qoQ2b3m
6IDmVdWIvKhHENTLw5tYrLKBREcdd08mOurQs03RtbBQLvFDUbGWqPaqTk175aA5yBI3QXZzSRer
h0lgyr0he/TP/7e5KnjUa80OUWYrRp5GVrvYmI1cAq/T/dQq5dUzFMZraMnnSElWnDdfRAMm5O9U
3P2dsh0B1bmbXapwPOJ+zGoFvanb/SiVAH/yz7p7akiB+9qCiTWc6ecr9hy/l8x4YNdpjn3Ose0N
Cljk/rgh9VqzU50Bz/2Q8BCh+PayILon3uN2yZNN+OIAGFQNSiiNNvIjs+BYY3ve7JFq2m/QVNUp
j9Ocgcq7Whg7r4xgT+tQa0wcrJg4wVOtL2gzxmQ/XRPAZqZYAv1BE9pncYaNhXjwPvi0ESnfWRKS
Z+d1sh98j0FVz986kIwY59TmJg/g+nIlQ/1cOW8qnA6agzwGePdCvMoi0pVsa15UIBXAg/ExNJ1e
fh+uruuFDHqm3oI6toJ1ie6a0ae4McqS9o5MYL1eNyrMGoeFj9XnyVbDXk5H+1CUyIk7wDGzeIQw
Frq5hAs/7b+jaxRgHkc6fkHQ4HUCFqq5fSHK0w/u7L4HTHzZewrB66/0rGvtkcmtHffyiLYQPTOY
g4kDf+hI2VYuLf3COgi4/FVQHyRd/e1O6tLmmzuMDmdVzDiiMLvPiba+5i2ZB16RKTwbIYUzQbXy
GyUwWMpgUFHg5kRoNgb7SRgZHEc2o3aXvQcy3hV36oMvq0t5lYIVZEATDu3v2dXa/i8ZjDrAxecZ
xdLyEscV9ChTRd2mBur2Sww2dorG+sk5OwrnaiFQaxTkrXbCkqgnQwAhQovsCl+Zq0RuzaUnoMDA
EHhqJd56aaZKkPxpgZKr5Pzscxq7nINNHLTVj2V72Pe01qnd3lw5+5mexvyTC1LPiEj2cNvc8eAw
QxfSffWl7e++8SIalNqCsaUjEwWglHW3Hx8Hf6vWHe/SPPkHoLCASh4/XjhgQzYuIHl0g6h/noeB
NmyUghfYycD337dzQbsRE5B/zNkd+d2aQFRKIMEGM7ZB5nbUEyoDdNI22KCfrAl/PCRzjNetuTBU
S8J1MIioTpgfeXbS5nfVhiqYiESLBJBIZzqrchjxV+2P5ogg/jt4QYZQp5yT+kDCTv26wvhxCc8T
Mvx7DGy4L7zLcF5ll0WLqppdNKKnCva9lImzUq9IxukCDoTGAfX2yhhYCgE+QWF/rCKiCN6syx/8
IvIyMj1tPGkLqv4mmkwgN3tKuyinB/U76aHubldoB5RqBGsmovFyWjq5rOyigguH7A/FYOUxSCIP
GfiVAg9gXyWITzz3ohTSH3M39M1C40LggMzv8w02fwmPcyxOO8DQFFJyTFQ8MaU1Y9y06gPUxcVd
nw4ogxLcMLeYZJsiI98oFTtJK2it0S4fD32QeHs8nFEbxnpuMlgUWeUdFSsZP2k3Zu5FEIO/kxki
UiZQ/JMKU9qNsvYnx8YDKuOM0/O2BKkzCpeChJtLlsAx9khpXjrvhM3oiAu4kxhcGMCxBEnQZ9I/
u1Jmo4CbDejQoV3g0Y0zhal+nKe2u6Y2sUB61qguiGUZ/ZJqCtrwVXA5bwMXb+DYo17MiKtBYlIj
qfgos9ZSdJoZoPOm8WKorcqttQLwH5gWtS+ci2A4ym2hsDgoUC3Ia6R+gQoJ2kg87vS+8bu2+4FL
D4npKJ5o1X0uEe93CMAFuQzXeyl1MbpirgGcDFBHK4Jli91Rci4I45Rg0XfURceB1ixDdS403Or1
wNLc7OXdemN+PjAqThMzHrdk7+bf70zDzEH9KhXuIugsvOrxtwKRj8+//MfABywqEklqhKq/BBQH
r3L9gMrajxsDjnQLEogkwz0XKozULd3nq9OrC90Ksu+dl/VZWh7s1rIxQM93VenDN7k1hM2l+Otd
UWVBbpdJGYyWcxIGnhHPvZgk9UQCgjNPt5nYaQG9a8JyRejzeCcQGMWvyQsX6Szk4NjJDRfR+2w0
zLe5jfpDzGGi5Wv0bFch3SFsGTCCKQoxke/U4lh6uylFirta/5IeoFb50HJyKlsqN54sF08sVHSm
R/BayHgXF5rJAOIDD6ayW/ZHVf9sczPaQkkLbgxFIrw4ZgnGqnTxHQuzmfUWNDBSSZ1HKmzu1GmH
/8ny2f/WdXbCn/v8l5IjC0zbTru5rzIiXSKpntsyjYhP2K9IpPcg/pjNww0yIV5Ksirb3f1icinA
ne2GUXfC7R0poBJ6kdw5P4EqtgSNmGp1QidmLMA741hHdG8WxXq9LS3RFyoljiS/dg7ruTF3gEF4
0BTia8NtGX2vPqQWzKiPap2DL1j7nIiG0yXrOafbw17WYvnplnuu7qu8uKtAMxXw/2dkpeQ08iyu
rWftOm4xZ8WtTMg+k/wGkpl9bBssDCENiK7vMMNR/0fGFH8vLZonUG5+Wg/Qq4BP1Zb6OvrRz1eE
yCkfLqM16AHe7L64KxvDICVLxeGqHfJQ8A3wTdDKIdWLWJ2CTL3eUya1Ihw1hGlu559m+N2u4CKb
f70lgROrLkayQYSHZm1DeePJApC8vk4nMZsPQ6qaB8pIrJ3QQVQeXRraFtfX+fKRbvjnO09MqSY8
U27wYNOoI4JY5BT/WD6pR4E2cI/HIKSaWMtxWA14xsLvElMzdZmx11/QlvfMYtDqOTmdWgDQvqL4
0y14y3azrIBl1sSAvN1REgACNjshP0l2MQ5B+0C7KUn7TxAACUsmJQw18NPtBaZviiF7381CMJjC
QCan58//TQGp1T0BT/Zhmr8Kdy1Q1Aw/WttlPHTcWXyxxSMNOmiE9p49Gt44mxF8FFYYgSEzlRe0
oy/EdI1LaFhfLzWTbUKwtjT4IQUN9/0DEZqgqDzc605RrgSNSWZxJwsI6yulkhFc3sU3pZBagU+9
C6G9es80kEwvx+Sn+9/dTJJgVh81D1UhbS2ulaKfFaN5d7CSJOxCPaG9Cgv0hK4RpgcxMt1DtXiD
0Rb1Fv5+RocBFvwB/8isC7yevtgzLgjWKOXx2p4YawXQh29F6mfyFcv1sD4qNLwpJ5YKf+vegYH3
0JHXzGMqjyudLsXh0WocOuZz3rPHPZwWZbLMGfCSWYhK1WZMZyU7fK1QFKMpLDmRaxpk5YzrtWFH
P7eBfrGr2VqOa4rAI+LE5hGkZtUFiwIDCv5wfX4GPk8WYzjQ99PD2ILAjoFU5RX5hrB01OSnO2bs
bhEwAgqoC1iLs3fIv0doFHjRWsGh+//NszvtnMNTdghjAHcJedgBElW5/PwjcaRl2egUBdBOOhmo
K/nm33AxFQUnKJbw0s7LErmd32QuQmDaZhpVKq6DhZ+a2dqZXA6E1d/0JpsH+8aT6Ym4Lm3colOJ
wjeTIgAzJ7/yzlYvGyq6jB7Om4pI9iuINHaCFuRuibL3qAGtTXD7BimSNSqTVSNvuH8gdOrmYoPu
kEoqEukyNjBe/HLTFYVxSUHNIkMj5+5EDPB/UGPzW9divPhpY9ZQYn03eqlX7vKhi7xEoysYVb/Z
PS/1a38CaZXyS+wlg2eLtFTW59GW+ANSP8nDDvMUBNCcq0RrufdyX8615sxZsnGCKkPennjGMmk8
WJfuCVa6DcvdnXYTHQuF2UHAWFxrQGrgFVcGT/HsnLTQ5/CRcwL8NOdr+Eto6rrn+YUE4VxFQyqb
v8DSCB0i0k2ia6LhJFGvPrYirh5UGcNwD8B6mILgQUmzDZ5UDkf0CmWgpXqRxMeGjKkecsF594Ni
EuIHPJZmgc8jpx/YZf/SF1hVyc0w86HETADCNaugaoqkWEsnS6NA2mH4a9RwJIEELa228ACpzXY6
hqo7Y20Hod73BZhJJazlIJ2+/NjmVJFs35UfwWzIl7id2HL4yyBIikH30Hu2C+4ypMXqdcF5dgyh
kgJx1zXZoUdSzQ1d5DAPWm3h2C5Vh4aXcKcK3qen4fqrv3EC0NuPVbeFP+0cRkMgHx6SbOwEbhon
AihBfqbTFNAjzolM/z0Pbd34qZIJEooa08TTrNcmw7cl08CzVz9i2Jv5f6vpQop6c0j9s/p9+/GY
e7T2zYcVgRBrmlZHFZLjVWtCDUKkb2qrJ0bIkMyDh38f70tPZRGj8PSXvmC92xuAvVRjZN6YPVrI
2DiqD7FgvdYMmMGSd8zSPsFF6KPXx+M1iwT49HOaZVdT+Yhtm1eQJ28PRwSupDmiVCA594kgbrce
rIqjt+hdwwh2OGj7bRy8PXP19joIfHcs0pG0e8M8n2RJ9nZ+p1jO7JwglGO8eIu9VEjquu1JzM2B
VmzyNVQHRZKHGAud9oeBCjcMDVs+iUQakP2TUCYxSXeAxoj0lnR9acOb7kVU8H59yX5NsBS7ClhQ
bHr4dKRzUPgrUgpSyo3r3jZJ0d8PypckpCSXYcluSRgq99DZ1aaQFdPfhZheyTYTzYqybc36c6zW
1EPlUDhldPbAA/Gs4nQiX9eYxO1M09275GxozeGIEsJtSJxif1DbY/p93LKq6pNALumOZ4yImDNw
RTwD3HZPK69IygK4an3Vfzc7x1/mQyPmcJYuKyY1ybJtbSSsnCerRCGPMnziE23ifddMurt333dV
9IOeTf5hkGgrQkkLWRCLjvFdPxSEppTRGobemlOFk9Z3rdEEfqQ8VGw7COd7CZQFmAjT4CdZln1L
koz+K/9yb8wNpOZnmDgLkUSa2QRFkbrj6Dj8PJIFIhk3wpAkmxF+EjZIDTC4PyOnMamcRK/nbadG
CTkO11IUEWvIwBcM7iLnmfRbiHv4IqnHKiCh/ozXTSPLL6H/AGwWnlcEQh4Pw9TZ4L3orCcQeKXE
Tw9HKPv1hl01xNyxGDitdoy8P7TW+b6OIuCyVHFZ5/CQyD4zSn7fckUAGocSgJx5OzljwUKfUBeI
olwQHl8xLjuz1jAa7Ign1KVNitDm0DPqzxX2qjAT+CQbwVKfwPx5avXINL4tkEHghlelvKGZtGsc
EESN/AVIFtlmfDsS0Vm56EDVUW2pV1Eqs6SGpTccIAuhLvFnRcc55LhEUUKw1WP8hnPAknA2ibzI
uiLmRo8qKkhW82vwKridF/kyr/qltW+W3MkSYrD9LjxXIn67nwTlL34yW/qwGcqPp1U4Ur80+kwC
vxkb473djpS4rt1CKupByxg3aQi5v3Pl3n1V0d+3VsHW3ejDabYYH4KZGK/cTVcPfBQG9phdIgJA
lFeZv3fWX6h+AGEQnsq1YAQENXhOWeKMjh69sgmFx3bxia/KY1nRMYmJ7OA+QxfC7Gva5gd8ZBT0
Z8VgECzzlC8skd0KgrdhE7KRRp5gU5HfAqoaXki0poaa7iB3QLjZeCyb0V61Lp3rEjPyXEMsU/ou
4P6D2VmWcuUh30jBeLCz+sMtDXQ6+fpKQSYsdQx+Iy+9TepsI/IFLyesNh2GC8nm8HMXeMniKAZk
pWklCp2L6WTA1HjkAH2jujSg/w9tLKLt8gP7FYfI50dYt+prnz72zpWb7uZ5gU/FHwjP8FB1aFn9
xc0ZGBwLZPA8IvuM/lYnWk2Cv/IF8Fzu16uKUANQwMwqjbt3Fo/ygTCeQLBBy/8YjDO3L/x8o+1f
0kfbFPfaVm+ztXMFZoMVJLcw7XzuV97ATJ/vmfhuazEm39jzz46m8VghBaXQoF2hLhRpTCIu0ABN
ElxvXs9GASuNq4XJ/f77m0dIMZSI0SJJEV4alkZeNlxA7dEpb6YSG8F7sz+CE28s36HdSbP5F3Gk
6ikb4XqE1fRCBS/16opekMEOPWMMpiSHTk4dUJWPkscl7kjM4JhwP9snymxMav8tuTuGL/uGz4DM
rhP1GVcpO2yg4dPraKcc14tr33YEuYhHWo8fiB0YMD59xGSuoPyGnJUGlHNGalbpGeAJfWJ0pSab
idftekc6v+Jv4wlHFWD9K+SkJq5OtE4eTnQexsnPRfSHv9rhB2nUaYeYDGR0EsS8WP6PmTe5UhaO
UpFWmpl6ZQH7BN7pXDw4K5oJOrEN1/TzU2QyvdnQRfMyA3LxScyw/Z9ccWUoKN8i7rNXnZZg5zwL
AtEbvHCfjrWanrG3R1YiIbYMk/2cCtWD999VkOk6L+69CFupMeTLMcLdEnyudqyeI2MNkD5MeNu/
XEKa1pfipACOPhBWWuoETGowiCeDU47ovciw/YW5YKqc4x+ObTr7mwSUPxBPr37wmAxKKfbo96Bu
vhe/qxqbZicZkAHt0LqnRRmIUNumlOLZ6szlfzd9JkZSUSuGP655pEwFtts/J3ZaubkgCFAJB0xR
7XBcLiXRvvz64Aj0pE86m8UO6I2ZehY/+uSnuVz7VKKxxxbJV84mw8XdhzpC91BQlqp4tgIOUMET
8TZRn//TpzSBha4/NdDK7czkmBBwfkmftQ4RmNzBWDAymM4zJOda8/lr1o3LHnu/e+qbueIAbtX0
Ps6Vf9KLx88beQVlVclihUbDemwzPWz454pF+3B6acjgfOvurMR7Nb3oBUFq7otv8yk2x4CNUoEx
eW0891FsVc+edkvkmo2iVftyryrUgN+MI5E+x9aqTaIWxsvOyY8IUcMPX6elavB9aLgrCxsgdr1P
pZSbiR/zwA9O8heXJB1BpfbUv33eyo42ORQtfyKvBz9CfqlmfsMFmbZNgThdBpMzCzJI1nMVBuSQ
Erim9m2hP+9B2oACwVCXY1yHVr45nzxQ/hUOu4/4Wt2orRT5NChlcHWg3r77JKsXACKsB4BFOU6X
/3940glxrg/1h55SZC64NQhrOT+WCg4WRCc/7REJQGBMSMtT44pbcCXX6aqB3GVnaRqIIjv0m5EO
A+gr6HTIp9x0vtHb2PWRA7vHZOeMSVtViZ+HcVPetdt81S13inY0uSOH2OssA1nUJspqp9pJV0o8
N1ug2I2SQ8tY4EmbWlaFKt1KNZncucT3u1LNGtSr1sAD5EzdAzwAisXwMEaiSo9VDiE1fg6lRYnI
f6kbj3iLBCdQoqMG6SMCPxj60jrsmdG8vNFQsdhbkWNIj73VLXXWOw53eEH2QBNwbq6NpOMLTKDj
Ij5z1Vrl8El/Ah1W2GFxJ3WQ1uyGzY/lX+BnbRwtibDlZ2W0x45i5ZbEewaWnE6YcFqIIcwCxIUb
7cW+cQ/31SHNU7zj/TqBFBuAwXCNKbpAYInByjdDqzUIGj4MuA1fWC/3FFLwNHPZoJDQ18n2iarX
z0j7U469XX9JL/7e+R1hrl5KMrgApLP5XiE1ufNITCKNUGbOEbpUSJHXYcJrvZuZuAAn7xbGruEs
kTzP3tBCGOODQi4zDNbeks5PhMeNkkeGM7/LC36qTG7hQp2nVn5qt5b+u8+h4SO2h2+IHwymr/dm
HdnMfb8fiOJErHMswVcl9zIe0TNzphjJMruRHpZbGy78Xn8ZoJRusf+xWL9XfMlCb4I10fD2yT4m
OL2q/LglwVmjFbimMEb9uOycEBnV32KcKdQEjYGDVpFmshz3FrXwCusBCUJCpJsnUZAx1hghNggs
d7fZQbhu9EBBFl9FxWKcHbdfCqovMq2hL1TJZRXGGwSZXQg+8Bmdgh5AG1kmMNy4dBwFrSxeGtka
RyoyqkIAY2wOqVmEWSRDCwac2g460SybL6Zuf/SEf8RSrACqe9Y7WjohS6PolLooZNmA7ZPqIeqe
c6h7NhyARjBc7qtnuSz7avGt8hmdFtlicyHrGy1rp+JqwIssAHJugJUJtGPlRdKmiAOFD/ChEz6s
XCNBvBaS5/5kMgrqvMlXbNOYI0CcUykhsNfr815Ya3X934RV1MdyZz8Wk+xW+iM9jH0Cw5akh4bT
nSco5EP2a1Moidv5L2Hb31EM9YW2JqckoL+4EoGMjrEEL8nD1pMPdtKT8SqQWXTISOyfyAVYAavg
3eIOe4DtG733ntFrIDSFjC0nAdCwHU+2bGOksgvE4ZgM/B5xmRmibTumGnzCKAOQeDZfAc1LsiUK
eg0ZvyuPFfifJLBP5fA80gV0pgw0WM3ilCblkSADlnYsX5173RR+x+BXPg6rPn0O/Th4AJwU5KDh
17HOx8Dc3umFAB1N/u/+nxEhtJMadnyot98OlO/zcBWtrFsyciYvvicVnyBy+yi150kU3hLmvG/q
Nwgb6f9Wog0tR6MUPDJe+vWBms1zSXTrVHb5iK/6uN5gsY3YDkfUly/Y6CBEx2pPeTr2RXjSk7eP
rnD4zoa3IYRlxL3Mefk1IozFr5iazoNLEyiR/qBnXmRwnh4tUrDNl9r3pCpCVULldZ8gH7Hhpeqv
ljlNMJXOu1TD/kMqVJvz3PMHwrGvXi8dTkTKnFlBqOxFb79M+yoRS4g5UtL5mUO68am5JbR8tJg+
sPtRu0BxfbMZIh5JcxKGcXotP3Nb7aqslhtwFTJxGQv0FZaOoO4GTsMtDJ9b8w9a4bG9AskkljWT
h7Sm+fNOWwdzeuU87ttQk+xoIL3e6uA9UQOIE6FH3wZWR+xRCaBsrgyyFi33OjdGsQV81ZDPVzbh
QpKowhWe0Totsfw9TPG6PtmySXJBS7sGElO06VUDHUyFeeRxZgkw/SwPlBnerd5XfoDmul9B9gaO
clGY/kiIRjmABIstQ/4lII5mNWvqfIA9TMsjxIQa8LrMjCYa3pJQVp9eCnnunkn5W0k4ko/2mg9p
0rrPBbtPFzgH3Aw8ahkb276NtGVP3qCaJmuawf1Nkg1sqqHlIqGbVtnvFJ2VpMBhDNUwCGOd63S6
+8CDBn5S+v7UpwKQXM7xrRLGkxTtbmJWYv1HYwTedBL0ZxDN/U49zbTnKQHdbEpuX884I7uyrsps
kG/jrbVS+Bcdn5uMRpReC5s5HxwLbXyIqhnKsh0f98psxbtlbZNvxUSjX5Yh6nq4ZEOJkdUuLQAb
2ZtezVc3HZXsVUSoua4wAQi7i/Y4ClJ6GxKSnguqJtHnBaKdM0r2ADVpj2y9GzXSUXSvhP8iiUzB
HoDmLI2JpzzuWYtAKza/7zXipbyVrTqSbVW8vETjckd2OQyqADXSQ0KMQb5dn0jhRisP5+IjOzPC
uNt53A4CKnMDPaOn7TlqO74+B6zppZJh5MDg25ebBRgIuW7iblex9sNj83n/jVFX6NwVG3iI5Wmd
GUzksp25K4U+pJxKdG8b/UIZB5VHiU09naJ2Bz81z/JgYFwB0HSGjgrRRHO7/5FmKTCNVG3byZWF
nEfskOLJgRc4xkjePfPQXgxy9I+PwDGraJgqvYADte6cFEBaeI0U6DOoNCt6wvha29vQyP1cGOTw
1BZhJ32YJye5KYOPPSEbdOcsJnZe7mjRELyTSOF609yy0Jmyh/uicxR+zLeEUWce6vC3oDGjVr2C
ciGIeGLapK7Z3J5owQKWvjNKR90vmNWn4iUOonnKlC1kMmIihdCyn3mozsN5w08IOBkgqBATDO/f
GDEo+35KYWaZl+sId7RgN3RH5Hxjoh0+flFH0DtnasjFWB9tWXyM4aiBnNIxI860JSfQQwAMIaH1
/O0KHxmHJwQLh01xR87J7bpEFKdIXdwSdE4aIdxO5otY5+1dUiOB9Fc9Pm91wOEfElV5GK5fctll
7AM3YcdK36nbMpklRTl7+MI84GyrSLQDlDwa8r5nuVuwfk4D3eb8RtLQGntGwIOcNEpYC9Qa5pat
7JWv0cxuZcQLaVZIWv9WWPKzRiUKs9WgnBXx/8e6DeDyagqiOkdjdnyEvVFSMjSfUnBgnzu2MBRK
FpYP8yqvHtBzD9lcd/dYpMOXzg0rlb/cTqGnelHeJ/UoFLi0I253End43XgOq23HvX2cN54PH98b
XmdvD/0s4z068A8NLk2TXUA42JHmPd4j7eBOfeBQp1wEwNsMFUFMSv33bqdLYQrJnyequgjpGMYS
A82pgxd71caWP8EIXP5Wf82D4u1seQIv0+/5z3dMxoTwxWBB41WCzivrHCSB+b0x8+TnpgOcCyGZ
NXqbl061gXUH27m/u/dKlxuofdbIle6NZnNX/WjEm/RwAfZO6iX3RCUIZ42+9nM3J4R2uhHqswgX
+nPho7fzhXk8tMPv+OIplQvdM3ckAAfJxkRLUefaDC0ViVzHzM2+gajSxnpvE0+9ydYXb3tWiFgT
R+HY79/Muqw+GqWfuOTYPmIe+58ZC8CRyMlHJdx6QhlsyFLw1LkRqTKhzarwq/koo7VDY7ouIvpw
Zgqvjv162ekY1erx9NRqwGIoDE2ihnTrGptQ/0Azpu05vBqp6jkAE+EN7kk7IFeINRqJKITBMSOK
NklwJg3L31D8lNBTJq8xpE0yuEzXLirVpkImyssJImIKfpdSbpIavS+tsOJAuG40OJAX+3KXEFmJ
Fh4VdLvpjkI34nIxOtqaTFSesO4r3ePof9TpWhaU+dMTuxqUdC+jj/NYnLybbhHo3F27Sc9un8qv
gKFkKcgDb0H8ycTSOXFwkLaq0V9lxGx0+RMcLLUVbZtIZYNQW4hlveEthwDVdfARa2Mln5awSXDI
nsw2wq/5WsuqLNW9K4+DhcKodNz9wTETLsYecWdURhbH1ibGjt2XKnrnpv5agSGYZZ6ByZ972kO1
J3h6dkZjVI9FCdFSqGF2C7FfkrO7LpAmUCyrdNvMIvC7RSt3ES2dMSHELrFrrzHms9Gy/pRW4BdD
xOiofmuueYIxhbbIL3OdyIo032lun7OGgv6guHYM2i0ezLFdgFF9yOxhyE+kBBjS64umAMVAiXJK
2a5YDbLamA/F+2t9i5/CrVsWZrg6I0X04DBR16ZOlfBS00QU/UGcaL27BdlvxNgJbchSRhPYPykC
mr1wQRYSYeD2ipA+5ydW/JmIn3gbDIXJ5ElT7CvONNFSJy+Ci0i5zghYWQcYCBNYLcMp2jNLooW1
W2oKpEVKqKxK8rO7b6wYiEKFcGu4A5D4tFP5jc2rYHMr/QwSbHvOxbj567yhi3kE6Pzs2/Yo0D/o
jUkz7p+pBDn+vri0GtTsyvwnSoDaE+v9co1clF2MfYrmVOdQ9V2XVcD0cjATwOfs35FJiJEYILvt
rnSmi5cYZIlUlXxW/iSBqPjWN32ooSiBWJubrCphPj12Tkxck1RX2eAZm5n9PgD7UFhUZ8JxiM3q
d21llDAdPzQLzr40CH+Y89N38kLwYjx8S5sT0aD1bdHi+TU+64ETLRpzGECcYVugv6+WAmMDbjPx
kgNKOKm1d6Gwy3r8//uatNphG1EXIxRpQAzbCeziQedc+tfR8en7YQ0/0n5uHk8M75AteC+eZ9Wv
TNcxBEA7W4K+9lFLThgheZda5d7b4Pt6sDgWXFzG8+yGnJ6D8WwEvwk4Yhsm/dQqzNd98RnqfxG9
YN1pupqPoyvgqb3WrDdBdF01e7Kta1u0IkLzONYBTQO8Mu7MOwRpLlV3f0KSbXYhBq7SgwFsXa/t
vEb+y6ibjhUpXaP05uHtXJTrckiDGNAO8o8xfRdIDGywJfCOrVDb68VyqsoeOZIgp576nzM+PMxN
dR338UL5zzzTiflIgpHoqIb7Zq9svxAJEIwuKQQtHKJ0p7YFYoTowGQQvhvUa++vLHGIth5cw1qg
EhRLuJ7IxOHvU1pvOY2wrE7STWvSdaeuuK7lfGZP64u41+jKLbEQsyEy08F/J1yf/ThXo6gf9Muk
HcqQ20+tZfuhDg9GwECCztixUZKqyqaloV32qmNTNscIEz5XaN7r0sl/AHQ6rpOAzKcXTYD31KIg
uqJz1/H/RkmL7hpGjaL4kCVUpUCv154FMHtC1nTJwhqLMAOHCBpQbf3eDt5MPkfdZfeTkvHBExXC
u5PNXpzhie1e8G6yZlp33ZB1QJv2abliZ1GbV8sw5dpsMPOkGYeOBNDEV1NAEyBa5JJ1mrcqgkLm
QL55Lk0WPYmflrWLzMhgH775b2GifgdTY0FpUqeApKYCl0cw2YekVnMmDprciE/c6ExyUSQ/P3eM
GA0WA8vGpeUPC88ifXzJ/gbu6DuBz/BuTZrgXaQSVdJF85z2ehZePUBKCYNpJ5l4CZ8ZOsdmXTuA
VJwU83Kvupae1gaP8PTxDSQY92beyOEWMaxCx/3PBg/NlX/9CS/qmIGvjroJsFWoaqGBgKfclG0M
5j+v45FrhnmqVwYKC2QObZrNsUNH28zhoxThHJDjzENSxY8P5bsi+u1UKLK6jjKtZiDWD3xDQvZa
Ch1oPRf6+9M7Qbaa2jrUQ4VFRZnKY7YjsyE5U/NRvLL2ElE692qL1dYdZl/03tzH0BCXdRV2GL0n
d9CeuZsg8a/QKc8C4fVQzmO7xgngbD2fD/Yio55OjcnWc+Zwm/URISzjAfx7evJwhVKYdOkFxCfV
9h6t+s4PCHBP8Pm82auG8oqK5IFFOAd0sXIdc45QdH/vaE6hTiyrmOnMstjRRoChY2oSalpCA2kG
iYzhUPeNpBAGpwZgKXdFu2z92n9s8En4dJfjXcIfl1I2UoFHa7QWJ6O4QfFqSnKAJ+9S9c11A8po
ox/vs0Ryah3NQc1qtFZASabUIwvFFl9nXZgeeUoLVO8uyh+eT0YSH92SCxFqd/i208gb3QtkK62j
ZU17B91FMAHYKm/jhtCWEgJ8hRr40aI8nqz8P0gZMoyLzKnkxkVU8DaCsG8rSedbB37Sh7foOU/T
f26Oxp1QDmbSVPGXe/W3ZxqEHtxqIX8IG66t97Sb64itLXE7Yuy8S9YgFhT6aezb2WBTBsBdwz8w
lzG089VqoRft7w+bjtqdUAsii5nn1ISPD0+SwNSG+RR9DjFpuTECGU+VKq3OUwwcyC5sHkyg6Ppn
1dbl3/1iazhLL09KE31kaETdmIo7tVJ1ltg+iflsftGdnL9ivj2NQh37nVtjlVcp1P/iG9BKFLxC
IgsgKBDSP7H1nHPYDwx7WevBZckt8MhaKDKMmuK6I+Ms4t4nGzHQ7CYSAVpZVNcwNKn1dE6k+Nds
NqSDoiJZZ88g49L/GH/JZxYqiEkiWcjTUgEKKZV1NKHnwTyBDYne/Egc7bYyk2+NFKclHsvhF6Du
hl4rY3LPJxGlomMiIe+rtK/wQixV210hAaD6pg8jZ0HnwjBLN4u2wULXxeI8ON9PCsjTmfTNFUGB
6PbEbws2XF5sKcXra8J+ZynPpj9KP/lmkLm+9vicy175yaNZgFNXlMkUii4r4Q80oTA1+RsUlXMT
L/Ha48P/HAQ9vtcWZeTDU524VH8dlWl8nnD7ggxgh+DxVTyCxURYWFkDeWe7OdHdtWdRXzxKZkwF
HWbaDiyuI1OLf/YBIVpHowBEQPVRUIbOT/ScI/eZsj6Irj4TrulQI+5Teh3CSm3PYuYpifGzFxKO
0DFFJ8UMKq70g7RZ6qC08UzH8tQfE+ef2ONx+K2kA3dCFQplRgJJuMPApZkLzGvjg9gyCnQNHf0j
C1GHqYAZ+L6IPSFBc/CrM46m+/886zpwYpUewYDZm6O67cwepOZzaJcMyxxzxD5L72zp7YIu+t6w
s1sKcbOaadU0tUCIsfO+SzTdbrY7Vu7c+VBZo49c6UfH9fcbnryekFkGBJD2P5xNWOx4/F/PD0TQ
Q1fvC87HThNorp8MCGUgjLaQ/I3ZNsMBWp/GamqEdN44lpmHqm3ryp/cJ23yfSH8jgroGbfBefZo
H82uj7asiyL1Lmne0z04eOERP02TPsJP8p9FDisGkFw8PhnM36hOfKWWV0PQNMurFm90YUUMXbAe
abuMeu4QUnGEGu16jcxl8m+EXcVlPldxz9F/Xj1q4X/9KGu7LY8aZP/4Uqndvd0IoSKWrhDReBAx
Fvhk5YHGYmflSjm5OQ4nNnO8CQwQQDQP6fWf2lUmER9A
`protect end_protected

