

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g7azmhtm6FcP7uNFjuXJjN8Z6yccOPk3SSjzvKB27peFKmnPmQmov5+YTGwYqqN9LpdyiUExk8K6
vPnJqontvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MFrqn2K0Cr7TmQ5al162oDGiY83d+AkTWOgFyXPYrTNznygR/tx44RAp24ytphNK9p6shs2EFMg/
Qqz0l8DCWiVEoJ/T8vMpnAn7Y+poGVGS1qAR3qE2njrl81VcGBZJeFaWIudhfr/DLTuuf2T/dWDU
YpelM3KbfYNPPiPy8PU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FZca5XZouG+/BYoQ8qrJTmnJanku4IprIWRkO6VciHehE5WehR0wsZJhfKlqLEeY1oTPA4bXaxmY
NjYkrop4EOwW8t47/hj2kFLI1OKUAE/TAhCGg/aNSOViUbB3dUomG/y+TBuDt9L6g0Arj1vb/5Pt
IChc5ZdEfRr1lJMTpFfP+5qmEH6lePPdzgPZATPB4Zrj0P6EyiEsU1FKBuAKd9iYNGiLCxVomaz0
3/RwK2Nl+/l4mc7PJt5Hso+4s1qHb4s2wD+OgbIwdH26ZkEnKVFpaLiuWQKu9uhDLGnsBMPf7XDE
p29f+mrvP9Zi/3nonA2aBKrTwR7XuH+ZYoakxA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jP68OjlYJglq3zpmKrXOhq7Sex8XNW8fQKp4hUNmuw06OOoKhQASNTnjtyVjAIk/VXb64ViBu1ds
cNMJybDSWBhnChfJq4h9PNybShGJXxSm3NDOo5wUHKf10Eti3fSotB9rVks+tNdTEZo4O97kgfdD
G1FNOqlsYcQiShEGLLiEQ2yYtgJBxJ+jc8mFjIEfPhAYy1ElrvtFEpnhkNS2LfE7xdWOQdO/XoKK
ibeY08pgncTI3pvO6TMbXushf0AX2S7hgfk8ysZrT+0gktqFrJnyR6oljS6VVPLtRNW2vo/cC8XQ
Bzvwwt4cpSo5KLS4XxB6qClZipItck2AUEdIbQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o7jAZIoXlFbFtDYmtXhfRBlb07dhBb6Wp03mlT4T0FXtvccSHWhWZgc+VUNwt6TohLihOwvSipPP
XVXpGL4pUVYNdQBCVpFzhMkt6jhyUgsF5t10yI5Of6YEfQrDHigceoBukM3+/zJHPprrPQE6FUvC
wXSGhBCXnHJs1R+n4l0714w8/WftPQhlD9QGQp1qT2VARQXUKBRxcRjxe9TcLfs0P4xnN7uHu0R6
JTmV+MHmhGpetSZGx+B2Wa1MQofUPURqwE70IwBoUhdXH8+39DT5I6x2+wMY6RcVATnhNd2BCgPd
RzAhwfrcqRiU9aB+eNNdFR8ve9M2nGMmV2JxZg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cl1Dz+fZIDYEIQuUd0pSg+5jknmtX/JERd+yOZ2SRaVra/4pU/eCTjEXMzhz4VFGYB6dgUxMsGBk
nL2WNdn/uaSPpi6mNF0UHQvZik4pUkYPrnRbFveVqW8i1t95SG0RW96uD19206lWrp5U1lqc4fH7
sfKHi8ZpU3MAg0DOO0E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qqp76m2aV9ue8Qai7QUavb+lhRYdu/txrnwYLzwTe0vS0S2OD1vxr8VeIT3bF/ZuXlTGm4S/UCSF
bgOPp7VqEOeGNfsSPK+VpQ+foQMENCQYccwKquBDSg/sLjpPK9uuoGLBLxjw2OwsRzplVFXiPcRN
LYK1/FmCP7RJBNgmhh/ti99a+WSl6i2YIIRGocNplQlG8FXq8ZTTHd/x2Gtdf/zGvJOy/fNsos6S
Oq9yJ0rMmbGeWbri5c04gZM08pUmXBsivgOHm2IVEZZFM4SBqrsi0xa52hs2kelc3iKJcWiTvU3X
0fJP9qNFuIjXBPPZvEYwhVtIh6DwiIC2viSscQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
yf5tjj9PaOYCh6LMNWxh2N5RKXz7fV/oLu7RSmcqVODLH6DyTNrIGggRnRqfjHRt8rT1I7fXqicI
4zPKtFYS3W15G/9H+BApRo+KfptqtWiIyKiPVu+eDNrjUfK11qn9OriD/VRoGhA/9DVpDNXP7aJV
4hNm0e8lh+TVRhmA2owuiVvAYg6xJMSow44OG6MRdQFKDk/q2WBwrjLs+77gE2yg1zSjDaw0hqgb
wyBOHwZyg0mBmFgdWq+TjswUQBEUdXtQ3MvysgzFeK1zwc24TssIc4HUhZ6MWzK4NmeqIjn9bxcw
AwKuNCzFC9SLyZqk/qTk1T9iiluN6LbOwNJSJTq9mgC1mPCDwjFJsuiM1OdcU0heJcpYvIrMXhJu
5sht7GcRID7GQIKrkrUuk6ztEH9za4sdonn+bErMom1QjfxEbJ2nGzLn7Im2SMk6XVnuGmFi86v9
3NuNCzb9/JA4DWk/uTLANcAvS5GHfm/jEitxrvjtBW3qp9oKjHLv04BhJ+czM9LG6e5SXfPI1401
Z8FkxnbD/HpiWlLa3kYkcga/4TAXkWLpyG1KhNfYwY8vBuk+mRaEuoKE1Jy5J4VALx12rEwtH+HK
FtE6oo5i0qtZmEcW3JiUL4dw3tOxt9BnVz6JomQ3sQAajTg7tGIJ6O5cacCMlLRu4R+XrTTELaSd
V29/aVzFZI6e8YOJk8rwK4pP2uevM9t9G2Eg7iCZhj5BHd7s94Lzlc+zBOXlYZkAT9LuU2xj9UqL
GSrrkXepuVMqffL0SNDPjA/0R0MAzgMRqJoATFr+0K8sQq31O/tfxQVABBSvycsRWRS1n1vMapK1
GiSk5WJq6vGM99vc1oRrgw2A3lTfxqBMhmjGRU9Rcypth0KuhoYPUJLxBDyNKvGXzDuqu6Dhppeb
WXlZ7+VYganM1MXDrBd6F2NFty31ky2XSKLWGmDy6uu8AO/D8bSX8MX9pDCS5lrOIIg8DDqzQ5Gy
rFof09V9uOoT/27NbwQjiakHNpCfaQ1tnfmy8nbfBTIyjBneiuCc+z9sbr4sDQ5sqAW64Ai3k4+h
/kpGzytsMbRZceDy4wd7RM+QfH7V2EaC3AfPQxbxqzTC5egcQaGErc+d93lf6EFJYaL1gKAPyzED
vfrXedt8Moko/wIWj7F0yUGKASGsvDC8QieWeJ6yyOGmc6J7r/SncgXFwOoX04aCxb74ypODQJ1Q
ObkOeJteDqtZEGbxDTi2cOwBW31CTL2joWOTKzNuH2jmHFC7+XcrIwmOt680OiGWiFre6Wc+MX2S
tYdP89ocz35hphl3JeHn5NKQ9X2BRbNVhM/gxOeKikwr/RMaOGATn07oqJc5zOebr35xRv9gGbxa
kfvz51yD40qKZrgscLXjSDp8uSXpl1M7SY29Pwtcj72paYcedV4nBGjgoUonYiNk1AeFvYUaz0bS
JAcJWdQOeZW4ito0lu3nEzzl7qEydf4V5ZDaQt3LcUmVMCQ/2+1XUWToMrX3DmXKoXlf3sZ3eTbI
PlVn/gisPDDyh71qX4ybPWwzEv5SFQoXXulsJTZ78zsmW3xUaqHbWgL29JBM2GjA4srL03aP9Whf
OQNYmD5sbiw76fj6xKS1GM7MIjC6QOQWIk4QqeG3zKjPlWEaQfmeRReJ4whtwTsc1VOv0NNlH9F/
LNGcwwTfGO1maVKa79/Je1yDKpQb22APAsvQpPF7Uw/zZJaN5Y4HCZL0JYQ/FSEZllAAICuU4BYB
GMp00ocJx8iHMB7NfaA9zFuv/qoQdEtF66P9isRK8KybL+Sx4K3rAqWTThL9tglqGkDm9DfuvkC6
0h/6K5nQ2uxAP7Da2ACZfHHPHbjhNykAb5HjQTYcF3thX8/Mu7AxrhErbdyhCY1OWe1Q4ZZYYudZ
yia/3/mCs8DhV9APuf7TWaDCpYjY6X3a7ya/OZxJl/XQ4adqpCC0KHLax3DSzg84+hoLPaXpiJtv
9LAvwTOBnmc8DYTFZ/nKlIcx/Gh8Rf4ZiaEHCcPboVqrgeUvPC1WH6kd1myLyTYn8sI9o+u2aXIg
4SIO9bjSr8kiaSobKErSr+5oXEJewQgMTLHgrBU2/qW7ZyUXT7D7Q5lsKYnnabjGmkE9QZyTA1IO
k0J0tGlfxdBNcGNiiO6fKyZJVJta63P+nFcGpC9oPe1ujANmwCMHTrywjGIxMl8Jhz7p7mJh7T38
way3Fw+YDxZTEJ4vkI4j8j5bg8tb3Re8bm1dhJXS4Z2Kn3CWu/dQM0GfLA17UpHkBJmos7/WPAQ5
QW6d5JZ4lDZ+6ql/hn9t8+yd7cbL7Nhh7/9F961R7nRAtfDuiQa/lrlRFzzDs33neZ9e3xU97dJq
+rUQre+LO2q9AiCyNa69ypBQ82iX0bU37SgktsWMfEdmzrhMxcW6B8F5/H6L/DlqUpFy5pbvGVl6
PGUXcEuZV72lZx7TCl0Cpe2AH0hh01WayQ/A8GGnVevVEcg2X8tJUY07gntcWIT6UOuH2Du+Df2G
UjUZeRgqLXLOnAwxDuvBCT2/ps/L/mkwm6e5dDbYW97XJphJMuRUrthvvyHmV5U3KoeEYVAmgIcL
XZYV4FfkJYNDwy6Eio4C+IG8xQtJmu0H8ynzcc8qESRMUjWi6ZJ9hjtecNb4WymRxbS+s+9Wfi5z
eyg8/etRPuTZsZj7UGSbiEy9CXLIKH7h6GJi/v8SNBnfYfE1N62QH3ewtUllGKW9lPSSuI6x7Xb7
RXoQIku4T4BPIaBo2Z4YsBe1d5is9ytOlKUGbmAWtiYM+kWBVDIdBjp9eZWtiTnzwPr6lXulbUzQ
u89gmzzmuuaRVWBJzqKCm8XGmk7AtF9QzNDfO/wZjiJbLd0NZGDuwwpQ2v4whBfzt3nf0xZfAnnV
gCuEhg8cM/U7OfywP+BqGfyCfp9pZ0r94WmM559/JcaWbA4D/IcYQhtb5b6pKOHPd5Dleqb1r9g6
2BUAO2yV8lWBM0NW3wQq+e8gwLUAufdFkEbEwN6TTpn3Z0BG0unILRbChH7rC6MM/q9cClaPDdyq
uHUOqGmkmdzV8j9p0qIot5X8dJdrGCpkHvU0m/eTlzUjTeO78acCVCLQR5Sr7nqJ+SWGdojdUfCF
S4vST9rd2JzgVsQ/c7HcO7hhkmYkw/25CnFn+pxaIl7+Y7loE/ri4frEzmL0v8H78qVxeNCb6Vgd
tVChIQbolKeAg95TxIfx0fvjp+eH5jxYEIZb3lbvG3psbScytp8CyfMnXm0ubVevHViV+l1W7T5/
h5nfNgoMhotwdjNdQMWwCUmUB9oPjJSKJIan2CNEmyV1vibHep2IWZ0RQHt0QZqXpqfwvIX2cImM
X4M9I0OpNUQUP4D+f0uzBXvXgVdaQATh+wIszxdELAo4DCmfXuFboKqxwb1R6j7/1LejQtr/Ueo9
ZLiOVvR+0xef4+NsyzawUbL8BgvEN7CF4fjgxDJ6YGiOyTnqNszIaXAxat4bAZNQ3138MIvkQeSN
u0EDWdzed69jAG1an0JAL5Qzz3CBT7nVxa8AlL/5gLUdgWUoot34ZDG4bdkTRZeaYid0JIMaMJ+A
P7Y95v4TcCwiLV/d1Zg+hIHgMCMnJbDnU9wC7xrZCnMOUSlKYqzNSCd4weju/itpdM1bWpdJmvcN
F2xvLY7sZvE6IHNKEmEQoUXO2TK1FShpH9o72Dz63s2jrx7XLydcLjny3y7oDvksIl73MQv9Yn1E
Fud4TLI3ShhkiQcdTDUnLmCKL3XohjO3TuFDiDyqRtGN/ooDMrjE77pkkv/njTownoSe4est/l0e
DpvCqqTXXeGEVrPmac102NMv85G2sZXF7aNbhLqvZA/mFm7cX9EBNEEn1TfZQhEwC+NqObmjuCoN
+SX0VuW/ISPvJ8rpc+Bvdh/xbviNzIEjrfyrtI3PusWOB6ofAaFAgP/RHOpiVcHr2J3cbpMZGmKI
J6H9ertoGEqlf/s9//miIVBQj/J1bWKAHTR7bbcEzjelIUtMAzpr5OqDPvmHBb6K7u3eukie35hy
6+wrS5Lg2UVpOn6KVmw0+l/egDDSfpmgDpr1v4/2MvYek99lFK9iZbR+M+u5ZdC5/6Hq70/W2P0/
YiLbFZp88PJxdtZo3Dukcf4HatbgtA7R+ribd1ax/kQkIV/QYIqqOuPKoiN8wKvsI6sf0bbfPWEn
UzoVOhbjm/V25mZoCNhEz8TPnLh2SJ2ww7OerFWPH0EwPGtHAc3PudR6UCWkfsnLXCKyGTAcRoo2
i+IqGSQdv3OeXPIhWhrPOM/TbjurCePpRvnYyYdnMXOl3UTgVPnoivgOIYFAnxEsFPek4CHseosd
75MtDyqHwS3n72Ta+rVJnVzXMEbIdhGlNXAm+nK/3ZsXCMao+hCVztkl0MMeqFVHEEE0VGYC+kst
qHcAgmTYWLvBPcUT/jRYtRCVnajgWl5DhiAZMX2I/PfCL+DLC62JMWl31BqWgi+G3bmzZOcUTunf
Shvtj6yfT8ZD9+JI+RFMC8mAkt2u0cr2kpXZY1UPSqt2+v0xFnJRb3gMwr6I9OoRtWC17j6VNwaL
lYlj+sSB+l89GtvodC61wH0df4yF4cyhjHzEC6FgHwjftmmwHoXYyrHopnUOfo/fXtjk6V4Prx/N
xIn6B80HFzcIjh6JEBTNLNns0cKP8RGQBilMXet3ay3baPb7W1qG9HrUftXPByoA7d+6s3LluZ0m
wdAxCxqy87CTngNCNQ+1jQ6qCDEjSJjEzoFdugKzsPkLdH9QJHh1/nRNoT2/LHV6ILtqiHt1tgam
Vcbc9jcbtMj96wNJ81VqaFjGBdbTqf+9XgVlmowPGI8MwkNCX9UwDyPRTMlpl6sZre7bjH4sYWeA
BOQOTRTOlVYRQHs3c2EXLttz04X+66wPFr8E6QHLPoUsH0Kf6NbYVWx+QU6PxZ+PqA8mTK1NYTS4
9W9uFYgdi2K9rHWPjopEsALDtABfvJqZcy5htlXccmPaC4Ha3y2uG0qFmuAAC/mU+vXyY29urDo8
0rxUrGyNTdojef9LW5pKT0VKBqF3/8M7SD3K7+SAWLg2BQx8Mt/1YPDCcDpUZLuvImBihPxORGW3
k1s+Ac0/GzDBYL61N4uIJq9ot6sBXPy8GIh4F5yrUSCwm4jPjEM6nrGfnhncPEc1hAa0Q/3DYKMR
gI/i8WipiXU+gan3WRJ9BPG7tXbKwdfkwo2LybHWy0ljblgQfniTnk1GpFrZf2GTKTrsB0p9fTXC
omufLOKMYCJs5LoI0TIzPfbJEXZaYx+ykEVrKmNGCqpFfXyFEb1K5Bp13U9dEuo3rujbQTTEDU4B
hvjl2ct5BfNptleZtEtn33yUxmOZGc4Kcv84OucENXYzMFH25T6DXDAIx0Y9JBfKH8JV1jcn+zon
XzMclAIEfUQn6ZdMipJYR1+OFm3jEZd5jhspVY4ismE6yPP+tl08m0JfxxKvFhZN/rlbcbxj3shE
BFXXsishsHc/x5Md6U+0egwvtB1j8YB//Fb5M65qHsKZ10zOM8cCSHbjidQ5IxKTKDyZHCM2wvDe
EbAo+soXVHFHOEwHEXm4ov7K6a/7//GocPVK/EDJiagVLhoK9JIvgh6DKyj64BytSSr78KmiKAyO
rQT0zfn+iQU8Pt6zmYgTIlngsEhtnYwCKSFr8Ly3pwx5GW2piviFTuUr1oCCD8+zPo+UwXhAUmKO
fTmT5jg1hb6qlmTemfWxzcvvc8EHj/MaPfqmIz7s6CTB3EkyjUsDLAqJDQAxer3wt+f/sUXheg2y
P7CFC+8CPt2zcDQCygusvXkDfkUVfcmS7FVHZGG+0YA8MCo2mi3s1Qk1jdxjzb2V9LhTjdoHPBXJ
nLHeigRtuPxd8d6MFSFvPZh67SFzElbCdsHpLioN3vAnzP+pMXjVhwsmRqOMFz3mKreVnrzZJ8CG
4NwZHeUGUTa1rZNgMklTFyvBMl62t80QuURngA4BisgU5Mnx0n3CDyi2XvZAh5wTvEv8icJNOPAK
Ud4z6Mwc/TCTc+cSeJkM6+iA9k42MI5oAnjNdOXWMuAsoIQsFOZlVRDf5PA/vnObuCDqevPre6Y4
uq90qq/NdA9Y/7FX6R7K8tSarowgPfjxdyV0ZSlZ09/4RNytZfax5rKoqzc5jVIITK01OkUcsBzI
s/tQ27XVc7lmhHT4LgdrOMS2Zq91aC4idYzfmVGaJy+GtU+ld5m+ziJ0lARK4bjXwdPCCtAWMdEA
3RcGw1Solk7dSADKVI4wkgbTMYPEXsbIdIa/piqdKO2hdp2nIu26oUsFlxw0hi6IQO9AYxysqiYU
rtqmIw42CokNtSx67AcPEiGDf++d8cFGyFWvwOPje/+DAJ9EWJb6xMiike2Xzb9lSlJLpOYRDnn3
d7seQUhHQfbgcZjntOJd+GS6a5Fvc6Cw+cBs26fEhFHBh+RKnw/bZY6Um0HIWukaLhyxtjYGP1DC
SpT8OHu4SEq4s0KVH6BoAzKzNXKMR9Wsn6AmyAA3kudAyx2Abh0cD4KAC16z84m+uEsb6KBUyEfe
eiEPKJYJ7pT7ajsHN5pomth0Cqb/JB01ibHzeYrBWyCAJUddgvwDF5Y9DS2orlx9eh+MHnsBhGpi
3hB6HkN52AACij3fOgSmzYc9LSMqcqHl5hwf5aF+UF80akToXRZY4sNalavfbwUCs8WPocPjAa2T
RDnNgzNgSJgDLqHXhS+8Vq6eRvcYbS2EYj9x+t7mN/3C9m17su45XsT+CQ/oxBWUmGGvaCUZbWov
jRi194jm5SPVH2jrbNj45Xwb9KoCCjIRdTJ2opMVg689mLYEMRzMnGEJg68uTBj9fVM/gSktOcHq
ax3xau3qIMoU/oFeRvmxF/LxglbMIxyhSWuzBrZoIfEmtEAAsVLg8Lb9Ypi+9RjtXBo4y17YsiB6
73qNeeBoNTfWrv2HWno8zxOCst0HC8fjGo0eohhCEjfKBahNykV3BWDZYlCTL6hG+M60NoBmPO9q
rSTCgCl7lofMqkGkxpRN7K5fjJ98Cmp+uun4tzCns0/wE0OLpzz5hsHNhpZE8fYK/0pQiIn2FuIE
b4XqhpI/G4XSPJ+2Eji3cp485LpSTkEFwh2vvnfnC4+qZo+b7XWXNTn5NTxMhkUFhYaIVl1RGwjb
8d6VurbM0pMqZqtA+70Twb7m0GQ/eWW9DmW5Gj8D/WKLu8XcABMV137cQ//UxtNrA5Z64gadNetu
s/05hlamq/M802nyueU0e5o6LOi4SAKYUxryZ/DMo4Vm1tVLNP963gUArEQI7ECTF4DyPkdMnzRg
GIRIRAyOsa4mEiU4KAVCive67Z1l4kN4a2Yy13a/eiHX7UNG/RW2hU3KqzBW8j/Px9mrdho77Ztz
/B12n4JsCZquO9dAq2dWvgrzGln3WnSqzx5Ie8PDVr7NzaLUcH7oEMCaL7Vr5ihcLs8V+6LrF4rP
TKxk24scTpXF6cxF7ihSQL8cWDYG08fOQfNoOT6JmTq+N1rEU/leipbL/cCKVq8r6ANjG7WMNuOI
giTPE+k1fC+5Jcn7LUUdpVExpWAMJ98w5MvMi4+TNsQ/zDzM3tNLPNz924yKqwFsdIOHhyr6JamB
UKEDPRT3NSxthoaLHyL9ciqWffiogYe/vvw7uO3t1/Wy9dtt0ZqT7K08M4wJUkPpXb8MsqiZK5oN
wpl+xzym7mc6BO4Ux7iM1w2j3/+TKF9p9kRMPNWkgRIE8hwnuKNwO77INsAGcFtmi/4erMDrCRHd
CqgghwgoKcI7cJOAwhApwrddaat9tBtn9tj1K0IJ/PMmVo6KJgLF3lsfXE6k94PA05trDzY8ki/5
Q5YmJqEzJblu2Adexxv8V+7FodYS4bcah+fw5JJ0UjkeN5zV/HivOrjugHXtKhs9ZgokT6gAZqrJ
LxlU96aZmhcie/TKyaunLoVkR9o98B82X2egXAj7Sdp/M0fQS6inLBxKsuMuRtbYvC5yB5R3GxkL
SeeqS/yMceBMxfjA9ZY0oZNrrBYFps91xW3nldd/Wd9O/PqwpuENK63131tTyljJKF1cb3Qx8+fy
Pa3Oe0JGmNQA5jgTS56Aj4A1atCvUd1ZZUh81bYnH6spI1TO/lOWOnLMW/mEZbYwNM6/RtpyZELJ
NUhVicLlU659bfjvO4esaoyJ74h0+0k5mrpT30SjeYBY7YfMxtPmiADPfSzGevvKiDJeKYp9Nh25
WuMDCI9PcbjYa6i75fgCAB1x8RtmqkT3p66vYqiajz2IeAxDT/fcbileap0quJHGQ436dOpNk7lh
wOeACY/sjuWelPrQ617DOYQ9I91s/JBcSh//Y8hYWxRVl7aF2HTNbfXO1Bc9vN+3TYCandXBYAE1
WryHNu/QXKVwFdhuEcYcFluymeQcoZBi1rayGhk4ilj5IBw0bT35e9Il4jXTWek12axBOHZHKeb8
8vHHa57YEg4uhxSr7LeESvU/o1FVnJllZ6u7YvDnV65rMFmFpXSUt6rQHRgfDn2MZEbPvG4fEtAs
xQPvVM+wEZ5c8cvHBcSX8bYLFBC6zeyPmtT1O2Hu2C5BSybR1s+2QENa5vweH4n3XFmCtESBidgv
Kcq8IQPwXVHhMYogq4j9u7bVDecid8zQMDzIsfCKPLKq9vIFtSflzwNB8KuRtProEkmdfjdNFF5I
tnwrsNku6wGGFlD/NqGkxTC0osdlWmuPgd9P3S3K82xsYVQOGMnAK3qJutQEv1Mn+4ds9JQOp7l7
q7NF4Ts9j1OCfDF2iGgnVF47YNbVNGsWeHW1i8h8t0JDcGDcSm37xq3s0X6TdZhZVc1oOQHetM4n
IsIQFruN8IT+rubiG/Io96CW6LCiJpG0jTlwQDbYAe9t9t2V6QaKdTKTN5L3FMed1pwRA4dXkfqi
xxd/5RksQcu8cWr2A2WXRqgVJCxRQCQ6IUlPaVjm9lHdlsFYp/NzRh+oFvXi/L8u8SZSxPCtb0U4
QhHsDZtYfMeLFuVkhU3/1aGld8LbvnDkOUiy3Xz6K9wa1n1JZoa/g4f4cxGWDmrvABmzzttkHZvg
kDWy46VB0ObQQJSvEcdXsp6qNJFVQsJhxPAlJM1nyUESTOb7gxT0yAvqGTXgAABAo+Lvg6zWlNmS
JkRfoduObCdbaTcmGQ0Ie1CdZkAknb03ef9PXZoVA6UAvDpa2Pv1xSbaP9a1rzRAlbHwBFuYvFN5
LP4huJyGtbB+QLT26/Ymw7m4k40XPBg/HeAC3+fK6kydH1SxeA4A18YTLNlJdlqq6xVKCYQrLn6r
kAnaj4Of0wPM80n+g54EahIflxasc8l4PcNdzyV5G2NBLtCR6xoki7ubtdlRuG7H3MHSk4umLw1J
2Pjci4K84KDz14WE4r0Cl+QeSxPT73mdxTpp4/W7wfsCeh1Hjj1/YisESZp48X/8hEja+bTsZKS5
nssf8EjHcadnYHcYHgthY5JqYBZJRB7waiYZ+HLz/PhSjdR3Qd7IxMs9QqhcVhAtl9Nr4haWr0Sv
B8Ams4ITZSYxvSiieSF4HyR/GHxVwXQwX0/9BzwUlfiasDfbyOzjoFSbOvIZLjdmRkleCEEyqgAC
otYlcUiKG/C4QtF16kKrxiRzieY3Ue2C1yMUVCTLXULrB52MpNR/FC/hbp80gow6lADLewd+ksn/
v0dwRXScFVidNErs6VKUgnK/gbXByVcnYhUKbQs0hCBQAHKQb2TgZDrSjwPJiJ0yjJowZpaSY+l8
F2EElTaUvWphCSjAUQk0aBn5Q8c2PE07uokufOeO5Z8KhyQauMhoMkAIQ6FMk3a7HvMOzzdUeA9C
6YAtYNtDfumzs6iL4HbgJLHPmuMXg1uRPRcmaw3IKqYbIvir+0+qc21At7CgAf9zBZ/s9i8AFnt8
f11p5Rzj9TnVP3Ta2XaPn54S9+xgUMoh8/t5KgOCY7tZI6yneTNkOhS06b+iFAErVxjzracvLAFl
qqz7YGYiVd17MIv5X5eRJGm2XJsaAw75TylTCOvQhmTTa2IKqtFPwMehMbp/M2DlVWbpFDQSYFEf
rdPtuM/9AIcZRiLS5oPY4e5d192oV0niRbLcDA3wIc+u6DKdB4/gdzwHRl6v7021JZxwBUqXu8tS
oAVnxF/sJyl2DuETPQPSZB6HmM9aAeZxiecHdWd4l+1iIf5aX04yKGX0rCj9jbhGT6POyeGK/pv7
/iISyYsiZlHTftMhQaQiMZeMcYUibabIfdrgzfHdIyIJO30J4BpgfzZSncJRMJoMgu/fq4V1yKSV
o6ynpfDYweCUrucOSXsyNEyeBClYSp+owwQ+iwEr6f8QeKyXwZ317rCcsJLlvOfUycoxLYfpcDL+
/J2cmsmrr4909i1GYoOTmtcKvK83sucZkZZObOyrnkQsf9Gy+B7kD5OXhvXnDwUv+1hMRWxeiPNp
BALO5X1c19oQC9exUpVsvo5zKkDz8Ak6hSqErRG7T0L35fqM/1aVSJjdruA3t3BwgLq04ZRzX9kI
torWTfbg/ABeATznNRxxxNZgLveKI1WMYbNRBLhhkgoUW+QkdSr0xHiAH4e3nMioxV7hA4tnVDP4
nKAFBEOMIzZT93ZsNEnVzkLzLNq4bg3ns4mzKCAyV2FaB0jAhYYwNJX/eq9mNt65c3aYQzfdSJs5
RvN/c90Cit5yNww7f5k5I1MMmZmliCH7E1lJGXj4jNZnYeKF4ZejsQyPqRahcHGkb6FXRIXAJxHA
IueSIgqnRJcRNE1rHeztSr75cbFpu6kSHYYURHfY8d1GypKKNs5vMm9zEVlLzekzyAx1MLBQa288
Wa1DuqAfoak8wBAokLOvoKDKaApGnmLw2nAVS25uSnIAK9wrFHVkHdLj1fxvkC65NIPlNqx+qyXK
eQOc+629IAGJc/wy9AEsw6VKtzijmzHBHltBciFCil7CdEGeYlqVIo7I2puPF88dS+/1hNjnemXQ
2U7hWuhA1DqSno23jUUaNTfqUyayOiQP4hj3a49CenddzgVVNbddYj8HRf995wdkOI9gelXMfiQw
3/lyrKFwaADNSDIMaLjQO4/OgJbPCJaW2Jt5YDfA1qkSjDoI6AXiiDxzrAKDUG11oSSA/qv4u9tC
U8w/seS+Yim2RCpipxWooAZblUGZkrslygGEngJmizpagicysJZ1FiYPtN0cC5EsnBLFvh+uTgar
KElqB9Z1dkDuurRIHtf3Tc7O5Way/gf/CFQXT2MIsf4UWz9vUmyfd0bssBt6aSmzj0ITjHtpjsUA
DhSarWf82dZPp9aX94r7FFdDvXmJBFPsOb7ujKBqpoMD8jq48hBnPLDlexXntu6Y+dp8UZernsih
Mc33Dunjo7/QH4JsONUHn2aVrz8hLsZsVVJ4q3gbmfkqpm0lATaY1OB6FZdZO5ylBbGCCl8+Cjig
x9UbyTWiOWRBEta5gKQVcVmG+ebiOvkDu0P5LAlp+4DL4sIus+dbXOP8TZcTbf7lXY6Y3l9EnAQ3
fSj88x6rJxqzOq/eUP9r+V3jdy5tc6cHr7voOHBPqffTVbzhqdK3pIR3GCcEuF4jIxuKN4aR/rvy
Xhgf75zWxoXcZOFcMs/yL54W0x31Aus+MqKgOTJiVPwDbZtRnGx1eweF31eWCpvHhnUHK4KuvAkG
qcdNJ6hL78k5FxnrxdGzetHfpo4aBEP2O7pUuEaImZjzEbX4Yvpa6SoNJvWZzYhidGArRiOzpG9C
N+Vp94vgdPdzN2ZfhvQosqgVRI+F/O9zLRL4oDUL01wG3uQHfRlNRckW2QPOs8gPs2PiFCaSmLO4
nAkjOpcSZG4ihJXHvfkUP5Z/QGIY/sZ7AP5/PHu4oWPyllSS/0OOCdjrHqaMkxAMOFU4++fA6m1G
Lnw+kkFAhtWwclKbK1gApXjnkXQoa2q5u0BaQcGtEF8TA/r0iaylYp7jRp4+hKlkISN4AQq02tli
YbvVcs/tqHKjSFEJwL7UgaAF1iaa935jY9gHJr1LNWepejW+3PfLb3F6AMb19eXKhVZIGnVk+3mJ
8F1IlOl16Wmmu9kxQky0PVCSAgHWTOJTDrGoYgOgO/VEf1fERvqduo706GRLvm1jN4MgARswZFpK
NCjR66ysM5NWKlNIbGvOQhX3TVlnYZG3h3wSftpyHjMx4wceLkBFf6vduVxmZ9GSWjWrjg7/bhCL
jgrCUWU1LKrhos0FQJl/hQmJVJuOpFkXX1Ex0wpfuJCh+Ax+DQD3NpZaRLXdDmkd1KWsg1zpZ4cp
q7mx+lEit9WaBgujV+f88MUcGReoWRTP3QMneWOwfZJ85az+7rnPUcCfp35Um3nu7E7LpDihzEgI
BClEEvyLUg1rys7khAeLGjvkNPV+jWKMve8pfZaQkyGxfRMTSpJxDQin1qcJYTyGGHSbfcEdxUXS
YFgEi6R7bo5bgEKrc0VlYB/F1WR3WofL1suMnDhGQ3HPeFBOM0RVvqlUHGIQs7ZEAHmqQbYQ9taJ
eExxhllt3p5nMhTiL7LhCV8VJQ3ILbKDQsp6O7jQuezlTqUjsE8GnZNQ2MEqLapvTzkoycmirzTY
kUJE9RQW6dKe990RX4JBwERJD5MVQ8bf10Lv7k79MJaMPLYxEuLqMVO9apPvZsZ+LpoXZCJ6/2xe
1L74q0jHgcGaG083W5aOCshlMnm9YCSHCrR8Dv8KreuWHjT50DgEVl3pnKUNDDcV/TFHsbsKOXMO
KhFRkExJgaSUFHMopasOtovNx0u2WR1FGldqCvQjcNc+M+YSEEGFcTpp21mXgzp5k+uCDj+BVr+/
HZYC7rXRymMWtpz2mtjvR+eWiIvB/jgaC5UgoA53ck9czRwcoHd8+pFSJ9zGZbgPdeK1RlQXXUDa
cEDlGTpts6NqxFG7DrpGwVARiuRvfPizBu9IVbnIdetI8s+0Rn7+CfYF5N+vr6pKtak6K410HRib
t6Gm8/P9bjReF53w59XNBVOLN0J3U/GVrd4G2lW2my2S5BFBBBO6pFvCIZyNOmGsG8iZ6rtllt1b
Gl15EYKQqiyJVwnbfY54Vqux2RyBTTvKRxMswct7HrmOf/wpneXxj/RkgSRSOzCDNReKDYQOdT/M
ig87NQ4J6dnk4F0ZDiW6HyGdRuwqkmpfgJAODfsArXulVqQGDELjwNKiyUEmzeogKvTalneRy6pq
BulUUJh3eTs1Y3TbiyB9nxubzcIgVdh/db5YFIC54fHKt9qpaliG8jIsfIwejFHp4mPclINuozat
8yQoEE73c/D3eaYsOwW5f7e01ins9meeW8JgfHLbzZqqDDjItUSwF/wD4NrAzTHiRDb8xVHZqO7+
rh77wZvIEGYnHlZWUE98Q+T/M3LoM/ujN7h472+X03TwjxbVFjTSjsGUaxYgGRXiVN4FhOH98ZZA
YhvRdesvd3BEZxkMC9JFzKogN4VzYI1OoH9HiGGhi4CP3gMoUt3HOi3+Ua8+lC7Fo22u4JVhW8VV
c2DK4+kvaLkNjXIg0paJKqBPQIWiI3AwZrDVMDAdizBTnJsS5CnHlN/qj/6mRMWmAjfd/MH8EXtx
1UVbSAXDYEkSOsZ1Z3SkKTsrZf2QTG4S17Rm+0gBelFqrOMch2Zze0P4L3Ws15uMsy70hdDWxoQs
Nqvv+e5zlXd42wXUJpAOJcz+rmGEOz/QgVwL5SZMMr5wAivcMwKupwwwhBCTm3aedQXXh1d+a/+r
JY42+sOtYBsEXF0wB750gt5Vh/HVaZa7YJVIB2LZ0dxBixMU75+KWN+LMtDXbP5UtLTS+8qNbaZQ
ZT4ZSL1oI5JEcelqbrySQML3QNccURLB4MDG/VW6E9MBJP3U83kN3ixWJqHv48lDPXFm78t0W9iA
WqJyGBewj2RH2vKL1ulIiv12JXDyIX4SAfQCPKY/q75CPLB2egB/XJVG/aEt0ckDshjGl2rkqtDU
gG+NgKnxw+91fM2MJ26dm1bHMHzwsa+pa1DEaw43eMROxscdURjGe+JLaBZXAhc26nXJxuWW4s6w
kfNLONbCbwiUOhrhO/F1ndqJEfFzmeG81xZ270qz8sxwzOJfcsfDH2hOoMtFlIVM3/+Fp6ANk6VP
p7TbRiexp6CZtMj3S7KDCJ47x+kefEXL9i/zQOfo4noRcHj80Cq6o8U0FVmwc9NJ0+KkTlHr9WpH
CVgn10zsvdywGLKFOPs+sU2rMHE0D5utXqm+QScoO7KqdmQgGbbbI9NPMDW3Hx9TE0MZ0LEiKzzJ
Ae4QuJvm0SdVo/G+PY99+hQIG5L5nt2cfj/yjGRiiHzC4zSMaVXaYrG+baisFHkX9PrXkTbnfQu9
S6O1ik/GdWAz/BLqVU8/Btseo2tRun5gPo34FwXhcWM2wkDRgyqjMDNv4jhnruYDjAf1VRQxqTSP
Bn7PN6zmI6Mi0KLC8EdtjPn1yAG8hy7QPw5t6T/64F8xkKyMyaOeVMmKcfy4xm7z6bAOrL+UaOFu
embp5xS5Bs9igAo/Z/EzpX2AbVa8cmSTfafmnYuU4jWiomBWXp3Wxj3h7fgf5EHNLqth1S7GuDc3
enoUbZ7/Q5mK3nhiaE7RuXi1iiJH8aznFCdBriIRhP7ThB+vCl7W7BVvwj1Bqv2BicXVqOKxOge2
pRrqdULX8RNHXcoppWrfUL2KtHeRuKw5L2Gz5WSNL/8NYRqka/K3bCWKEy8zhnNCdcEwP/Ldnb49
8a6/XuoGUVXK8ALR6QZNW6nlSegf4VBSnBu+E7rgLR4Z2PrLf5ltpQOsOm8irA6FcJeIfd8mkNwF
8VapTMdRGDG7rf7thNtzEXT2jX9SkXrNIqhnfPN2FOw19kToj741H0wngHm+jQ6h+0JPvJTJ0GZ/
HsKUyO4giEh8wjBobLuLhoBonQCnqeXXNwozOcOqMTcOqj+cQ1Dy2oM+cwV3Qr/EvbrkcZi/SDKA
gEB43ymDZxbWntJzsHPaqT8PblpTZDqCirVGi6342HqZnF6/FOcDLigdC/8AuOW0AwLK5rCdt18+
mN3eTaEinvlkVjXJ56ln6NaRBVaX6aCgb3aAMOTViX7p6hRyS7adTVm1ma5Kclo+E5Nqg1p7gGR/
SMYYL2bqWpfNvDmAKHXRlPFv7PmqI0AncCALSr1AAWQRY9M3LFGm2NAkxbbO+nNbThec4hnDn1E/
Wiy9Lyh8IyPmQdYMbShXnJ8yQFcbKPeOb2WKEus8OokeTLm6jp0YjYEQZJNEaoS48V+EciDOMuuW
OI3gCoc/4JWu7S7I3KhEH2yRb1X/sMojgq8GAkH17dSMX/zQESYEBRWxnBEjmlFom6Dow/xt2o1m
Ywg5Nvu3Y+suaM5Z78ZKmluYUgEz8brJKywtlFvtmXIaYVwugSFRTLlB4iHnHd0csY4f0/MmFiz2
4//ftltiNzdwkOKv6fPBNZO66tFA0Ftu76hGht0VemBIdHEdN8HWSgp3DGJVyK6AsuI+5rs9pGQb
PkUzk12ab3K/0V3djTwFjqZ5B29Gbf+KRxP90oqvGY2EFKb5Gk9xfp389mrnIqwyvPo1PgRIJiJ3
xpmxlqEU8FT1uDpFLwWvKs25Hc5WdOdQVbH0FBT6+RwfA1NpfIZCRNbLmCtxGymb+Ru332EATGOR
p2oRkoMq9t8Sx3eRaRooeFta5uNNasu8C+TuilJOO1JAT8y4kg4pbjBH/192MPbPOOgnyn0hb+7f
jgcYP6SLKuXrdNuLRd/r23XkO87C7tLgYgJYZQlvMGv/hShxKohMU3fd6CuVMWTJ+x5yNAbwZjMu
Dhx75TXQxBhnZENRQodZ+k8u5MDDiDGvyYXMt5IwGrudLo4k6mN0zu1qNv7eVUvpCl/5IedqKoBJ
nFbG0mQDCGnLK3zwbKxjCnY05u010zakKUkqC7q8cUNq35X0m5QiPafi90XuFxpljyD5u6ocRvw7
LFDex2opucnY92Jp3mf8THgsbPed8sejvp8kH9ZK7eWL20zeLnuyUEBhPVgxrB597nQV5FDhSjc9
yt5Bl2L0ZRiahh34dfISjsniF5Gs65Fi5Rw3+Ej7cnBbicpMxtTCPtndj2l15brwwA8y+u6TTfXJ
BnfpM31qxCefAM1PprqRcato+I+1o9Z1YuTH7X5EpDH/+OwcNOxz6yU159ltf3rUKKjfBCNubUNX
oVHLnSc6E20h/JQPztCFkSd2n0CTh+/N5iXCpXjirwtsxfn1xqmDfuKnVs9Gl1moGxIZCDdk8PWq
rSz+kQvnjbQBQigL0BOZ+C5kMApZiZujmBNGbKjUFTcakl5Jry5MISERJoJCAy6/ahqFJdSBU/Rt
UJXYBCokxYuBrymf4q/+PZxtnNGUzb76Y2DLcd/03BBGbDjETr79GAHU4/fkCIY/Zwxxb71r8/Os
t1iMTocGDQkgkiA5Em98on8+aQ66Kxz4Zzclj3f2xEWNE3Mkl2wrpnHuaInTbvITVamQ7Ipa1tbP
SF8pMcucb/XhVXhzjzifczqgtHJ3up55Wt4r8y7QwJt2+cHOJyl/2gxFEGv9x9tg/BrvEEpnjFH6
LW0PHK41XC4s595zIiZ5I7PBABAmJ/JkCO8rDk+P6xvAR+EG+8i31ls5PEv0JmOyNLm2ghG/1Sw9
me7gzjg0iN4eUcclHhAJCZvbujmRstQOy20uqwnOEgsSznuXZ1YKbP8GOzOXV4Y+dIlRXDDSGDuJ
5Qxobiwc9tIzwYJgmR9z/Z02tgDNNzEvq/b9Ijai+o1IT61iuimrK3ecjw7tnoc6vfC3rWLxcWWn
0sVt6TLGtiZjrOG6ncTMI0srSFn2oUFiN7xqxGOwHdcCagIRwRir2zXtxm8XTMkV1eK5u88Xvw03
dn8TLUJJqoyqQbhmGHYQ6Q1hJBthJZ4RpppLREiPFn7N/iowgyBl1D5jsLoEWWhyRa4MjPTm81VN
Mqi40qZVaMLAj+yG1nz6p/IHYSEB24Vv0Nrw9IqbfIZ3IymAPadeiigChn8W/cDwk3dYvi6A/l8b
Mr3UtTNbzMx40WorPfMwzHAcfPDFwuoYpsIkmYcDeTtgHPQK4mrq2Dh3ky39OJ/iZZL8uYe3Dd8/
gN6DfnqFD4Vo865veTUfA7tX4nWMzuhpjgesvJUBFWADYvGD5AurD1Z6dugYJxLgt/ScayKupEO1
34zXQ+vCLVoEAlwTvjGyxTrHS98tAeZsWUfROZE857OM95Ja2jYPXkueUYCBdgiQmHVxsx9BRU1B
FMPz59khvcirgiN7nqmL/aVcmThALCZ26dOMC6/2fIV4dOGefg3tU/t5yefFLtKfxQcPIY7jNNhU
v0/MUInPcGGGBEyyk9VzKQfi/VvZxoky/prux7P3G9lBco8158Iy+fhjbH81oJNhnwYjsOD37mBK
z3sy1zrAcnFpYqwswCkQiVcgb6E82vkSlLt+hrPZ2YIMWNHMM5kI26vGHxnuSlbLYsuqrmK7uB6T
Zb/zB0aBkSw5Q8IqwOfDH4f4f42f8dmKTFxbbI5V1AkNXvVSeDU5vqMqIrxVvnWb9NsgXytWjBfB
o2UCtAmV8ofb3ZK5Gg8OBxmgKTGOKU4v2KbBzrlvON3jvhD72NuZSEmQg70//yBZNjS7XCwvzkt8
AqzcTBYa02VCcf9ydbFaNPYCXZh+h5vrSi+PQ9SOrQR3IT+wRdFhnhtMniyA44r355N2C13QgV7e
18FK10AQ0aqZdAP1nOyR4W4O5mXo0eU5LPs2GVouIauwDnTTFMV/6Q36uKRLhpX2s2krJmRl2QRm
wV8tqIjDppfyT1Yw9NX4f+ihBW3Pdw7xx0/qQN2ohQb0aL/KD3uWwix2oWTo5cxeJsxqVHhJ7ojm
mJDK1svaBLf809bnAhIpGxY9dxvujnM8MZfTkyexU3HUagX75Bna6vNfY/6PE7/GQGFtm5sMne/e
rzBCrqqdh5Esl2XJjrSdn8hzFLib3HeZu87K8ZJvkz+iPQkKxN05vc6NsiqwiNPAcdA7UBKaKoG4
O4mXgsrpiR/03D8C4SHaWJPqUmUIMiZvcn9SZWqyUJqu71AqJlAfQrReLQgClzToiS/kMgutpNlP
R8SJi6REuP/QvvTTBB4QskJFDscWlAFzIHloIanHNG3yb7VzWp9C1TJpJdvD1Q/FUskWpIcQ3zj+
/NQXEpA7tj5wJLMAu485UUuPPLInx9RJtl7QNE79CPKkLtSjD3hhMzdBgYbVlTVnV1WF11IBGnMv
yzgCQ+UK4+Pf2aT5ZYRllYgC3pYMUj4xIibN/B7JpwYSr7yS8RmDVnHFN2+QRcEaRjjZ0+GynBV/
2ZmOlRYPr7AMcke9bPq0iqi8K71wuDsDQjSH+2MY89PXVzyyRUoIjkG3sWH/eX2jWAykAzneBF7B
tfD+w9fJ7rMjcLaIWnlZk4Lob1Bua4bxlO/sdLL5c/PNqWLFNQ6i73vTPu8x9x590E2djxVtl+3d
m/Hq5Ry8g5NBc+bt0y20cJYR8BziAExlMi1ovEoZUZBXNlVjaUSxvvUkm1gjF3oUOJIO0x/h57qO
4cIAe02YEym22lKai4tJeGNCoxX26o8f1fExE+7GyFWQW84gqP2lEsxfS7lDUEiNkhNcD4SN0q2u
9xnTlwpJ8kB7L/VfvSNwAV07Vr9bDMfb72EOSRq2HI7OhlJvE17/s84Ne60toyKXUPCq2NkB/TO0
Rpho1WOFzqKm+hhSpg6RW0bg91S0Jw5aXkEB59sMyW50OLZPbpxilx7yM3u/fsRvaYDpJYAlt2Nn
t6VjqauR5X+SVpx5Gsn8AmUUlwCaEVr8DcJ63XXPTK5fKKC2sVUzrNfogC4ge5lJnEBxmEBxd2fH
AS5h17UUGI6dJ8JnOvDITtl4JTBByfbNQ2J0wI660+V6YyLuFRHtY5PRumPjVt8jgVNpuocunX8Z
TaWGEAHz88huCgq3HI7qm9QDNpDiADuchyX0XD51t3WwALoQP1yV1COOeGw9tkcs3c+MZ3aE5js0
S2TYfab83PCrCB9OnrthMk/493y1aEtKnsH1Uydi9Eb8YI0i6iogU5sIbhJdO1P9E0swvV2/LIND
qTTE93AVYeazwf3YDyj+QqsfQbcL1W8Tf636hVOMWfR+LRuz9BiXYERoUx+Od/Gpak0p+Tzh6+ML
sYnd6sGqUf4Yx3VetQUQsg2JfEBr1Ch3PWowsQJv4HQPex63MZkEAo6NQ3VfO1W6kUJ31bp0/vpW
VD/nS0ehW8QLdNmeJhPOuveAru5meWbEiPTivdAaywyj0WVLSg+3Kso2SJyWK9RFzeiH41opxDD0
6Ccu+Ld5weAVm6g15wpNvgA225cd0lcJQzg4WWh8Wcdhra6ra8CVX3IBEGp3vS2D57tqYV7Q02Rt
+D9mjVbxJDJDDfEQHvfLtL0UjTHEAfqDcnXZNpR0hfhEVjvsihYVH8B2ShVfcPdxaYKANOKsrOii
lSkGgymL0V3KsXQeFlR3VmB4qrnwOQIodNw3x3xXOQ0GRMSNTJjeNLMaUullDbJdbpT1a5raoWDk
Y1FRkBfnZokHoIgOcyHe8gAdtIZKSiFfDmA0irX1evBwDhaBlS8iIE93UQNPs+hl/laYwD2J3s38
BhjLjKYZwZ05C2PsBqzmlZzHbCvboCC+o7AShAt8CaSeQbu1cfDxw95gtLPti5jNZwD7XYoFDQwN
ggW5gGAb4V61hN9NEZBxUZjDG85klDg6DQEXcruWxqwagsFTI8BvqxC1piHJmtGV6PZWE4OakjGt
1WaL6d8MAqh3w0c2T96Fxhq6GxurlOZeVX4059NgI7pdB+zJgDeKZJh24j6oYYjAtEqVLViA17Z1
ZwjINxkqykt2ErWJs+92i4BkmApgmB1URlRKgLoTALImulN+NNkkuJyJ8OXBqIT7/by8p/Abv8od
bCpzvJZ+cHyv3SXBIqGmjF+74vlyMqgEPqhWKYSGCMn8wtQbh9NRRK7nlcIJ5i3tQemimPZ3vdRA
uZiedNC3LK9JuCtj2toHJSlLiU8AG6f7+OSPpPi40+kP7feYrTeqecqTOsn4VlilY3Une0bfu0D0
3qT7jivQiBOZypnN28fbRray5s72M79sxEYBjfQXbHIT071IMWMoLbU2Sw6rHD4Mpgv/xMcppGLD
94KRgQqbPwb073jP6nsKFz6bOtct91nhwtV02Fa46cbO79AzKd/xjYp26R4yVWRgyfMlr3RH3ZG8
8va26R9oKUjQfwU1MJVLGxkX5v9k8yYfPpoD8w23NF3DBGeSt04krvQ8jCvIQ4lCxwhIYpb0y180
XyJtJaP4U/ZVNALg0l7f3Of4RxVojGMqLCs3rLJvoOcqW0l5fs9CNO9ZhQ5z+oGbhgBcDvdaUKe0
46g/fQt+lfJdnxurRNURFA3jxMn8Za7dC0GUDWhOfFjoSMom7kmPQMJgWhh3pLFL70rwmIZEt8VA
7A1/PVgJruURmyBBVdsZxENyQadryBpFVta0NdYNrTMqsG4OM+KPO4FI/NWwIyRi33cVceMDsa0v
if0PGfPs94enrOPvhpGuoQZaeYP2oqCzYCziT6bTffDD4w1Nv6HYWxLUSnc276Z3jH0QXWwwYDb/
mNHl2m8HCAODOoMDS+dXpH7q5uFwooLSG2Owl7UeHllOknF7YrW7pB0RDDCmpKnXAUgelbPjE3Co
8bkoPuyK6wiBcQ+vEJIgqe5tUUxrOtuKELAVyHETGGu9wXuC6+cI8WAplAGt1mFnDJ1sXNIAWEb2
Y+RbQHABfunexF+TFEytefaIKLvab5VxkpsXtzMIj6noxSTESQeObpbb8xANKPvHNeskXqFojGZs
qb7nS0/UA4rm9L1cNCzzDeTYhfr9OmBmFuz32K5AofxLJAy363XINpXejCHiXrL74hQ7/+IJg5h+
2JVb2tv0z6ra7K2t4KURr6nOU6q7bzeqSAnK5b6KagrZB0/ufrPC0Ufhc//qX678rfsQlDPG8ipQ
LKYn8hcg/GIilciYOLPMvdd74s8CzAUYD7odtI6A/orQ0yQSSuandyS21bI1mWFhE+K9X1u50SSv
QfWopJhXEpbcO7HEtanCm1fTzwNs97JjJWwPCiogcOvUTLcPyyifgJ1LSbQIwxnq9tROBe/H8EXN
njqbcbHtym1L0cZkhMCppVUwAeDjOMq40DN02ko/1rqQ+Miz2hLvmlFlKc/iJjFfbznWrtKp+N8j
uWcqJQ5RUWgHDmZvDHM+HwhXOctIaHNx2TmXp31i9BGHyQ7wSU98cSlN85hLo93HjMlpz932T/8y
94lCoV3FRjiIkLlBbU9jKJIYeQ+4nZL935gTC2dCA2CGpcln5Go7nNJDb7n0j6zS/gEtp0a0TGKQ
IH3BL731QjBB1/5WEpZenzuO1GKxeax/EUHo0w5Bn8GwSytZy7IsiqntIVOmxV+5y0a04NrMsZs9
kzBlmms9SMpoqGWmXzZCJlOcm6kpkdOzirn/CKf7RUbsUyBzQP5FniM52u2i5NFzUJJ7OmTl/6qy
TyvTw1C8zcJucpQGGAJP35+/bJ6/YRQLPHlWaHoUujh+ePn1yd1gz583WYs2yX1CjIyDl58iiO+L
Sos4fsBhXjyWlpjJ/zwZOM8znTDDI07O/cDCcM1rDAz1m4D3oOWkEQuF+6i2kI9qPcH+zKh213q7
b87EyqTCD1AjHmZQ5j3jfkZjPH2l8vVkeB/Ox3SpiO74MuCb6e+XkVJYhqKaUsNljFbcjZSpSsvk
skRDGTlwLJ4qqDR0+FcleGk5s2CpAz3WFhBC8044VlSK1417ZKkLjLzLoyYbP0h68xXaGdoXfarR
EZ+fWqUdCve/96LLS4em2KzQWFEJ1RCv+XPJzwMWrJ6jmnTFilSESAO/aikF9aRdw/YheNLnmef6
yohd6jy7leLs95VxAL/2Tezevb85vOVh4JTnxPkRNOl0LKQ4t0xPVH4kRzMef26k1tjqdHqqiQnN
cyL9GIEsFf+3lEmp2F7SyUkbH99UleYiUhwr5fh5bVcH4QrHWMFQkzjKb/yoGvwO6tttxT2LqCui
K9kKy0cQTtwvD386rZ3QNtSROUr8ubPo3m/lSMZjgthhkkUkpDf68WuGPo6DB5+OxK8eDBerngPK
XbRbvkgUjReU8zcsgMk/Y63Jar1CoWu9piIWQeOuXJqZRPlQADdudHRQMbcu+CS5pUR/vUfYnIX9
eDHJiH4a0szu0c3ezjPSiuknYc86HTolLZVdxIkXa7oOZoM/GMwOUFgDtubXyIi4+kqh8Hh8k1NX
Lv6+8ZgaP4vAilLx2tr1SLh6B27HqwpETQsXEmvsXcWhazZdC0DwFcyLcCFK/SxJ34pu0Xh9SjD5
QyB9btAJCAZ4p5kl3fays0nvtDik9XZsAFL4b2KZjU0I7vR9TFLE8uo+2nj+ZICuVXsQnCPzUj2k
EGuP1dHvYcAer+JW8/QWnwhdobkU3fOPjpOhqryDNSJL2cEKU5u+0T6iDjHvj6xhAhbOPt7Uve6v
F8rtO/LV26I/+Id3z8kp37fmDghP8/jQc8U4kYXtWAHBCcXfN2GMog3EvSJVRX8OrltuzHp1TO+U
dDRBuTdaYKPvvZ2uI7o99Oa7J7S50qKoLq3wEdJcYTvYhfTmvjNEttWEWa4RYn1Fi0RuVRD30lZu
4vvIcilX1L5weHvqaUbsUGjn6xTZy9HgOSwoscES+1bSwrI9CepPvYr16GmEfyebCKv1p58X3rkJ
A79n14LcvawTNUqo6kg9KNY2BCjGZHGLAgNlZsspwtoGtyGpliQ5ComBmbonsrZ3oAyV9HqDlswa
LWDY624QZXbGty9IGC/+0ucyDHvEiCqBU+Wv3eNuMmcFsB1nqoAS7uIzOldAQ+nPxiQftUicBBHY
YKFHPbLz2uJiQ0+ueiZsNNdlcdHekqM1Ai//lE8M+PS2UWnWJgYY1u+aUf7/Qvjnjk5012mQXKlg
0AzAB+8u6H3pTkuTIFvKWSBQXICopBqPCIYx1xDdGfVWJug2JpSbwmCRFaDPH/IKRXcVTSgoWT+k
xRMATp4H04Z4G7LG78MO9UUE6XmClFUiFTW8zbgp04tMPjop64lGnsRfmUjbrk2RkzdUik2FJV/Q
ORFFiq9yC4Wf8okUjRl1JR3ikxacfPWVKBOd1o1FCzwlMiZkbAWblcYmvfiZ5W+qUQ9oqqW8FQjM
nr+JIVmgYR5bqIlSiXum1TKg2ZWAA+TNKuVxZbcWdq+YslGrezo26a8pHBOm3m6HT99U5+9G7kN4
+6F2iVUJXJd/il181xwci4cVZxn/PROo74hpaiGZZqCj4aSkJtisYz7wcYimxEufblPYyscV4mGe
RcChWb9/+fNvHF/GyLPXvfoOFxEE01YJ7mtnQKv2X8+FfMzCqTrF5VP6ck/gdzk6oiCdviGN4PHC
Xp1atgIVcRh2LAbbSuKxwRh3KeLRkQjMHBzejIlgBzTHcFDZzn3AFUw+ytaXKhV91zOghWMBsaVl
gch6a60L0G2KHHFSE1/iryIntARDLhsFgxXtrtfMLngr3yDKOpQqFa1dchzYhS/GqsjV9oad1L0T
W46vPT2frWR1jM3qI204TtNT3Da90WH2+HTGNHl2gwAOTsZfk3iREPT3QxpqOhEZDar00HLRkeP4
T23NAi3yaUZFMGzZKp4gMDAfMZYyVG9TYyL6lMZHEgRn5SABM6Cw90o+lvnVnsHjZbbI6xMh/77J
yMKrHgJQjBDyq3xPkQSKBJL6vKTOZYiRCYIE4Sc2yTwTY75VW1El70KC7qg9nY7CxZa/J9Ucyref
ATPh4Ux+sQqEJQIXM9MRo13fJ4H3x4jSV/MCDfVlDzllXpBqwLf69cPTARsC6XldOvYzO3nqVase
oAUk+xOUypTvZBy7+CTGXsjWKsQ5xkxWhhB+1rFsdiqJMAX8d+ZXKiNgp8sAKxMC4whdLY5TSTIM
Mf5u6jZlqe2BWJ7B24cjR9P3uMX5HikCT0koR26AHSw8NHr5E9pqbGnmYCgsPrVDg0/6BFoYq/M2
MCBq/QdqaBiRxCdhm5oJymZxlN/4jx9k6rThZoSfe5mi5ztM86nOoSaC2o9y1Fv6Px6ZVFXZf4Xk
aKXKbKdsuQHG7eMPXjcJB9zjqSP98UE03Yik10NKwqFqoqrAscRJA3jwHgIxtAzFfTCxecX2sitx
XkhKoGVpkqd4g8wUPLjGFt4Bgy46DI8rdovVVkgzoydFyynZzVd0StQfNQGvFF0sNMNOFtQ6sGjX
jF1WbJtnxf+ME0kAYRcodCmdWWzmHdt+xVR5Ezx8rKcnxP+ejPf7KqtF6EEVuhYbXI3J0Sbra1Bx
dmIZYls/9/jL4hl9l8VRp1mnKKZ4g9x7u1dHxdb9xD9AZDZHYdxSkGiDwzdd7hmwGnSHybilwHUz
OzFcxcsA2PR4dxmehgBVhHe38N8Lsj4WiZCZEqadoNANhQF5iqeSfDTgxJbs2itssTJ7c+C08mHA
7ILIqStzWXic3/Pt3L0k0JMDXqItGnYJ2jWEwxV/qee66Rr3RL4sO6GN7mGLe9bxRJcWjlLGKJfF
HKg2Q9f+P4ydvTfW3lI/jbTPKYxUoiFC66X+2C3Fwmo3T5G6kxvaFipPk5Ry0mlwf/19Fq8a72Oi
js8E10CdDRfBSoJqyuvq6zuwg1Pel9eZrqRE/VvTJJnr4uFLcx/iTTQi8tFIhHuxCjTezUBvbq/j
EA13zyLy1O9T6kPZu3FR24mcwoFzEtcepQ/Bs4T4s4co0uR3kcIl/7cQONL0TjR3vMhN7rW47WFq
QPjCF37TzDtJbB509LGqIU//9pAJP6ZlKHiqy6PlaMZG5iD4/OJuTUvLaTOsIxIvXx4fYJHOlAFR
nxXOhB2qYvPr8Ml9Ft5aJby34enDzFyJcZAflGfPTkykQuDsuiCK5Rk8upj4dUaue/AeGMZBsz4Q
9eNkERTlNWHI33KGwMaqHq8NjZggt53B4EKaVwRndFG/HOiQPkIZlr9rWHlLR0qc3yTed0r2XlFo
GT1wf47RlKBLoFWUXjIOuWNEOMfrvzOrtjZDwZfvJPH+AtP1U5QQerM/JsGgD2rYQ8MLIXrjAyni
EACKC3zSXPYmaSh6m9ykpUDH889OIYP2NnTk8v0fiYxFBQGE/cw40nvopmCqtavwIYdsMyyvMGGh
T2DFnKieodGr4Rr3+0aEkB+VSr1tNjhYqMwFDpqrMjLgEGAcVrwslsU8V72NEKW7wgXZNWe6UYir
zNLb8HmmYPKO+YMNLQHhdqYFZakvWxZI5Fql3YR+tSYJCklbkmQ4q9pMZZ/2DvPOYYZEZAryK8FT
czqnKetqdI+Nya9eD7WaVxt40MN54waxK2nkAvkM5gjr6QaSekn8+P8stZnYzL5quPIIKr3oDyBe
/GEsvaN9NB6+RAMZ5MUZoMFa16wJ7I6e5OwMwcObyE0fmkhhXAhPFzgtG5LhRyr6LTJiSy2yzYh1
+wZ4dsRP65zfun0/tvt35/8EmthZxlALzG7/x8swi8aemomW5fU9tzgkGE59hSRKF4PIaDJxT6Z9
rWECF6/fYndmdWaSxmoZvLBEEFse5zvd9apzRWX8k/78WCgkw9hU7jlBGtMHROL81p2XkNGJb+QN
zWJG1I532PLsKiI7zuVCkQEbM4jZIQ8g8Q17Mdt+C1t+1msK5s3TQvUMhtqyH8GNqbPeTraMXfhY
LMS9ThBgOry2Rx5k8A/SzpNbkWTHqniyrqwdKkJGzmHuXnXs9wNeiPGmdAnyAA7cv1NiyP0BWGSl
3ZUUorMcxHklQldLz4lU47yRtU9gVJ7npRUDxCyc5Cd6IAHB7UcnAUWiimSIy/kGgZ4uelSGvprB
HrpzdHxK0lyjwVVrrL8RPOpfk3dx2QZcoNclP+BpVyz862X0otq6ibq1A8/J7mHC3tgNRlRoAdvz
u8hy+8rc9DxyFBr5KNxHa7+IG8hs0SZDJNEDsU1XsXpAl6Oxkm9KesWnDN8LNC8Xr/H2oA6GzbRN
yQqGNkG0IsGbW5l84qLC79RMhzOT63zJGFGo4QuAIbHOlpS6GArWBfavSeev9ZRMQy0WtTA0HnVA
JDsHu28dX6l9Rv7rzyaG2xv98vnHOW5krm507Sdkijcec8jhTfEuyeavtJ8OBDUjEbERvIN1qiGj
4jo8coBg1hP0P5f4QJ1zdu8dZPsm3VwqoLHlCxzGkpZ48kZ7HHVtujgBnXiGWB68Xjsdy7iMD10Y
Ie2zj9VF8giwUJqabrBuUKkCaRqjxAYWMSv39GOSAwogNz7h/UqUBApy8nSEyycK3BBiV2o2gELb
jWgPI6+Td+Od12RbVObSet7C/92fOOWORnaoKm9FimEpuWyO26xo8DvPzQDmQAJNbsIMiK+6E+mM
4XJepNZNaic/amm5TCz+Nxl/t5HbszyaYJTqYsTUIamUQe94rb/nXbWfskyqDzaK9jxpb5AsxO0g
KDTtuKDVlID+207tw0C9QbKTXU6UuukTzbGkPxP8PfVX5xBVbNrbH27yaSWOK+xaBCKn7UC85eCE
em7TCM9G/kkPfv4hIQx+PJHOPLSJdQbHxahEt0MYxu3TrkgSSgUXiFyN0vsOKlsx8Qv5D7GaZW+F
inumEexvTBwA6pRbSZCacmnC49iP0+ENkdhHLEnmXtlW6Bs8lO/hziQ1hJPmMBCvSttuSSJxawAh
dmKyEVV7sEYo8KKErQZPtmQXYa8yAErPlZLi2H33Djle8j7rP0OF9nX41+pU0vwUORo5QMkvk5M6
Ei5oQiS9P312zr8D1Bi8ZK4hk4nj6t9e2PheKZYVfqURDec/U1e20xQZbP03i1j1C9fShQQ+xRmh
x7SRDzxAx9xNzH8V0LQTUcs76+Z5Sqr1jfb6Xzlcu0dOaiRKzm2C8f5EP2EgsTzK7W1Q55P8+5qc
TMIYQfZpYeE97+QQFX8IsLb8mLZCkqvowSZzm6FPnPESiRbKRb7sqkhCso/jIgZycYzSyyGWYlrx
EJZaFb5UiCcJeysXEyrSyzPvAfM3NGhyBTT+GtWJ6xZWBaKRsPTnVIpgViqAR0vNuZb8uEHuEtNk
PJJwUqbGo33b12CA/ub5/gLZ/CF5HYILrwgp6Ufhhrx2dfVKHXdsjuWMEZ+GFu2LKN6Vg5H9Usy7
iMOentDt92ffPDpSuI3EZ3UYqU1Qk/PTthcQm6UDdhvPr/UwvavV/GoLZXrgiUWS8DTFubaHy+j3
AYFrtGhT0u0PifHphGQAM4nLM3OwvFkpc3XodemrS+DFfrycQA1vX3taupbWBWUaW2Ggxkq3MFAo
+jMW7/HClSOObd04c/YraRKzD+iX9uzej8rMEVs9eHL/fbfcrlaMOxjVXpQNnlumRyRxipzoNpsO
J28H/PbjYq1dE2uC1o/z4EKCxzopU+6HVtg9vd+1V6mPuzwvZWvXEE+TCxS6oV/7Sd2GubLlDjz9
6Uu9JqBBJj0x/nlD+Q5Ald8cm++zjXXNOhd8iRl+l0KcAzCDIF2BOezF6M3G7hOFrL7EwKMPrr80
Y6tsdvS7c/AcbNAQFD6Nemq2ZaKfbmyb2+ibK4Rk1CRGKzr1RC676U5j2j3ku4U/9Tod3Q5tZrKd
yHQTMw7B5e9HpDYIszNBraeX6KX+jjw1cZv5KCJ/qoDteOEzV3kwxo+taeaA/SVqZuJSgvFz+s3n
RZr+F0tTpOzKh5rUSmNOuNQsfZEnRSpKlOZnreJkv0jYgfVyhr0liEYIZKjbNwxMYrFaTx10AI3t
s9FROad2uJE5ApapYTp2/HmJDcILVBokCBXVd4GU/P1jEK14U86sIsGmFOxjWk1am2cQCeMUvpP+
8jztBYyjc+e+aXLHp+7cw+nvYNRWYF0IBwGfI/bZYEpoNcmbKz3uUdx5YF2W2Si/ZSFfZpwG0YVi
B/Ly0z1u2XVuwDx0HWkcq80hsomUzvOuDIXWxUN6jAjq8H8JWWvcJ3l70E7kTKAYMuqgGwjerv7T
71tKmckA9pSLGTDXQrEhRKoLMi+y4SBNaobQKyXdJ1lZ+f1C6MTR9mrqH985RIzMYCGXIN6PhwFm
TTgXWZPEYC72gkTt5hxn9veKUxQx1YefeWla+qEEniyV4oIlFqV91OUR+ZCZx1VBrmSojDx+bbT7
8ptFwkpQaJxJxxs8WRaKi49UwnwvlB1WoDDvI9/vxuUb7+ld8qPeVBifrda1inO1HwUgzyDxP9Io
HIqEHviSYYfpmduMDAT3RKZUMVUWBSC9MmhjwaffWalEPd6iZ0HZMDdavg5GIGtXQ3FGtHkGxIWd
GAU7AkCxXuFyYZ3Og6C1lS6hGzEl77ZE7QUBa7+7TXxAz5VOuOr0mK5YZGFPdEpQvHhslw2mKBuJ
P2zt3uNUHBS6wMj/K0orXK9xDQ7nVTHFuFkFBSpzXqa+X6nX/dm3rx/QNLlAgG1lgiM1+nvBhAAh
UQvV+WC4IY7cZOpLVIEgFHODkU/DsRG/fUcscvJZ7nVzKDgvEpqlJLtBr5m9AfvA0SEGAEvkyvpg
MqdpMn9bChxbhifUDrti1+7OuQMVdiS6jyCR2gtzexO/SgmWX7xI8IokYjsNMrOoq2h6HM630eOa
Am4Lcmojklzxs10usJ2b9xCpI8Des4Te1xcYqvE0cG1T7uFdpZWrm3P32iqafVmxLnLAPfQHdPuJ
VofRM9CQaBT2aPjB0JEPVBmvn0xwT0gwdwTlb8Z7Yu33DqhqQNPBDnOWsG5zjV+0+12Dt0AXyBt/
xBc2MRX3fJesD62Rp/r5PaN+5dVeGBn5Vq+P/iStMYonuZloou0xNFdzWaqvRvdyLXq02+JmrVHU
t+hvRcXIK2MCnFmVGC+O3wubI8l0UVDuhbCuqQMjsSKx8NrBhyAbJ+36L2dbOiVnHw/Cy0giRrjF
of6ftyRy8Y3onyX/caaozvoBOM7lmADD+dXNwA7Q7sD0I5H7rGZq5cj/FboIO8AAZFxpSrGS5Wau
oLOsK/tzVgDUMhMEYrOOE/9FpmRj0yt3V2rmy+zObLVWbfroNX4p0LPI83eeQY+llPGHQJEJI734
8cKnuih4+lzy4AKstu74XJQ0WoTJ270kLh2JBTTFUWP9Gj6dZElCAO4j/jf1j9djSTD0lftVwDZd
xT2GkTJ3tyVmvAXAWOE0Q/4SmxzRzeLVW1Dj5ycdNVMv8tMMJkPmDEBSDXChWOQ06KRmo2nVujac
5jEWel2Jzzn8j2FYNsjMF1ADstIlHqnSld84GuQF2ZSozyUu6yUZScpXgHJXZuXirFSKWYzREjZw
3hjiNpxhjj7KkluuGiphcTN4gwarRTBhAZpXgvM03mYQJzCzts5iaRvB3q/8cRTDjQQ8cnMbVCoz
4JGojK/QUFiGOM+OtMCLQrxKu5CyTZq7dUTh0TibypWT2ii1BOFl0Y++mhNoxNc4tfZh9LJ9Ic3y
E+Gcs3fed67BzUoWtnK75wb1RF0O0/3DjjceSJlhvCtUSR4i1Qja78QK7EaShvmiqGeqtLQp8t+H
hK9O9SBa2KZPhQcudpy//WKp9yO1NaiJNJjHmpo+nVDleMA61+HwVvhWKVwx8QHt47RQLvFW8a5A
h8ZAIFSHtFvdlAivDShHaOjznAfot4F2idvbMLEgoroMmonzhoRRYmUhxfpOdj2UNnaNJ84m6dWS
5nuJXTOZ2x05edLc1RRAiqGyliOwRyA8I1kAO/a1U/7w+bw6yUSID/keYzu04zZ0+cBMNomXaPJb
J418TXeHhDHKe9I84OBuJzZl5TmQmiREhGqVk0HUUbZ11kpf77Jjcb2Oisj02JzN2fB4g693mV7o
+kzGVvZNqqAG+KxilDLWn/A37435mmeoktMCBDziGEUVKgxe4gNQ9LcDBEMNuKn2Ca1NZYrd7TaW
Sy+vkgObSxqwi6puME0mBwgUdg+msmOyflUr4r7SGo60KseyadkTYwuYFHsvdX43MAUcJVNOzWYV
+bVjEa/Ia3wv3z3XIW576lPH3LaMbtWmSfb3dhIRuoXeg1+sKtvLApyP1Bkh1amgy++B1vVFLCH+
1fnfHd/h4ggIvmsl9vzwZqHsMsQy9omMveCmOvqJdDRGh+GPapOw9wWDIBs0cro5noEJxFhPlDB+
S0dAJrmFr/KdQ5zkgui92qQSEEmTZMRNq0xW953l7PvNikO6Rjnd9EJSfeozV5EeBJJXzszwmAxF
iqS948dsDDglQnLrCdmHpzO2ppkkskMcXkn1hHaw1E8iGjTQyKlNo0anW1tFecip5j3afMDB6Wv5
H2wg0FRGhJjMYvYRcZChzeh3ybdM+75+vgytI3Kl7z3q3mgWFTdeFCGIHoi4Q6FXBdfDmUrvrDb7
T8hC6TZ48IAnwjRAVRcCpHzGCA1yiI/UaeDjEWlZww9LouHXjxggWMgbEGGkq2hsMzkP/O1nRGjz
3hzSdhd+U4SffBli1LBiplLTS2aXIe6kx8/loHywPly/UmWV9qrwJ0e1lqOTxKVow2PDDw7F1eXA
bWnmhLQKLipo1Tgrshe3zyC3tGDBIRLdhxe0fmH1A6BCWU1nxcA4GrojkishNq3fSa5MMWgjoUs6
TMQciSTxzD3Zo0lHwJ/Vn/DEbjIjp8eFycN4iZDUZvEN3jsjsLBtMCJDvM6OMFV7h24zlDOQ3AWm
ztBUaMl2kAc2sIk6UFZ1Odp2XKGi0xB+Vshp4d5O1bwN937bY08B9rUxZ2m3rVcr4+SeBuhNLJBJ
6LfKu/sq9xj76CONHDDEVDsuPxe2X0Yw+b3wjjDWd2Ui2vOKUJuWtjWvdGx3dZIywh1ZjibbUWsq
QoiEC0C0Arepckxrob/Ypqu8wiQnrpm1nVpVTIlqqWhbE4OyVVB5JADHhx2SA0wDxPlXmiQwRXch
TA+hKwwvf0dtunptroc0zjCo8uG1xH7wCxW4moI4rAC0hBN1YYpemehzYNBWqG+/uLpS6cOGh0+5
FdIvvYbc4FQMJRPkKZMVkBBZEW9M9wOC/b6SgKIQKigTuHsv93ExYl9f6UcOYD+xx/tqs6MiXacI
iKK1Jpoy/3xkPEnsgrUeGv2NaCOpEoNPCmrdDmq/xxRUfhWwT807qNREBphlf858eoVpBOegIwbw
kIEjsebl1O3oDPhxYSdMXoIMCerDx6jeovRorEnf+ZxbdIyBwehqE0fJrFV9ANeUyRzsNnb0k0zi
Sq9oVtL6A3OdyJAw0USYvNcM3MxOR3LN8ekPgtg4PJajizVi4NRtnQ+fLo6kc0nZ1HPcSuHdoT0Z
FRbTHzMn6+D4eDM06iv7RuREQ4q8JfMwaiGC2Qm8cfuH6+vuzsqeg4Ge6ka53STvJcxGm2nkBYce
RkqQMbI/v4DBKIHj5O3L3jp5lwODs88zIElENXMmpV7Ui+7KAqnwZG4UvQ1AD/x2MHt0q+GWUmNq
nw2GZfpw3hKMHH9YjAk2WEU/VbgIRw5/hn0qfGDnzYJhzkMefSHqhWyydyTGSXWqhxnk0eZzkTGR
Ei2ZtZ2tvnDnaxRJudDFH0qo2SANdzMMvAVZIsb3lLPUCLFymlBf6U6Qm+/6jUkFMFCbC4Ufw2D5
4Lec+EGzWzSg+CV1MXmQrWzCnQYnN03/S5dEbsg8HXlMGVpFxdhm3chgqmCdTn8sSJwP4EmZjoyF
daRHp8hj4b2vYrzq3VcKrWcPPEhnHr0aKztcVqh+EYL9/qJCWeNPbS2lS0uYxBRBy4RGlz5YbStb
QqqfbLRfW6kIcHriCzA+dulToekfGHwFVGY4mlJhMNoi4Tx23b3c3JMl/vdIkf4n/4qzs/hcMmMD
WpcxmzEPjMjtGAjr0r0UNZi103R6UtbDlv/lgQzOY29C4QTYXTOKOFL8c07qHLJ4gBK+xOXm1QgL
y4fVuv7T7gjlLTZ0a+G9QFMqmNcPDwYkx/NjVfvYQudPWfULpk9Uc0vX9DUMsgvMIVWOu15Po6kG
pvSjiJauYZgIjFkvUy80gGZBgR2EX0ZZzixwcvhvMZAXZ2bS/+af2C5Nzdc9h+H7j+1D5jyEM9X9
IPOMsf7BpjJy/qfqqbhJBgHmo6qYJls6gKpxDCu5dH5OvyOr++1rgmAmQANHcP7fZ2mMPva+PLMW
c+5o8EJGMblP1JYO9YMR+uyk+jcZ0xijKonmzLfeOy0uhSaOm/8fIM5er2Z1wnovR9xTw/HDZ71C
WkDR+G/8Xf3jFGeCzGyTMKApVOnOtMu1YC4MnujmilOGJLscpqoRxjS/KRABMEdYY3Uy8NHut0DM
2xERTZMH36yARIB0iZZxiMKnWGC/zZTI+OFH4L3UC3xhwUEgGGUHcXUvXZ/yyQmm3CeACeVsr5oZ
Wg7+trBkdfwVMgE8xfltpERnoH2EQl9FlXK4PGZ8OId7irMRhsY2AQxq/eCnMgTZr6hcXHr1r192
TwmfJwP2vi8lMY/mMK1ICuCiyedcuL2dKhS3PZXzqzGVm37TyS4cVO6JAPKK8MhNA3TKYyV7mgUf
s5NdX0djo7HWSIRp0j4cmbHTkOYHeFYELPmSLLaGx1H9NdViyLI8gIk9JUBWQa9N4d5mKEH5hsZ4
sgm9hO2sNeYv2KLYgx0+bcZauyykANc1KksR5Ypii0mfym4GWELkD1HD05N4Qb0d+3AYRq5yI7QN
SCCYNmdcWtEC8dwCqd/FwHOoUQ6DjTYsIL5j8ozQcy2GuYbMZQU+j6sUUQp0vPPhM69RtLR2aG42
kHwB72W7mJZpjPxBtSAL9TZ9pTrLUj9MqjdK9pWgN1OCxcSEwckLBqHMXNhL8LMyHosqq8MFuHnK
V7+YFSzPS3pC2q8sWOgVM6K33zVjNhwj7g4BwSg7gIjaecfKHjY+Rzp/9KS2m9FxjjdgQtyeFOoH
s9+VXFjNrwb5W8bsnO5cfgjX8kiFwbxC6jkDMUfRvhEqN6riazJSBkNTri4AzChED0zYHgde3lUr
4WIpfYXrBHpdAWeRxFn2ApHtrWtEOTsjGyRG+qvs3WkpGZnBhj9hMXN5aKGOHQFGWaHVX0cdJFn6
jMi1duIGsiEh2gaiGuizYkDkMi4Ls8DgrLh0tktSbDi86A2R/cfHHMVL6aaKNJ11DDQB47UBMjWU
nmxRwWqabSvg+d2QYF+shqkUYoYXcn4qNPIDD+w/2g5UolA2nKzTUj72Ligu/FYdXlQLrSc95NXu
goAQqbQW4zhv4e7g+1MtydRUnLRIdZkh7a86+JUbWf28LDZxuNv40c1E6OIEKZtdaoo+XjlexygB
3URsKvNLaBKwg0WSsUeXz3JWZf4t4AtmK0reQkvJT2SxqpIo4XdG5YkyJDuu2Dm1hWdPG0IjUVQd
t9uKJjhz65XRw6/n/0HtMSvLc9N90BPSFdnYOG8RQvTwomzK14pa9vhN4MOKYJVewXFoI1iWv5bu
12afomDPdon/Pdvwg5UKB7scBX+0EuSBcsNM8j3SgTbOWU8NjPVzjSBKBXcacC6Dt2LtkWHqYeC6
vZSyg9YBeeC9P501N3wHfIh06hsikyqrApNmi0kGpF3MfAL+BEToZ6wq2nJ709FoHd3NU+oLQMAr
31SJkZqVmA/8Tbb9I+qOK8YuzfnyBBQ8CvKbp8NSYAmrd4d7thwUmYj6sLlbW6dWbdmo2upalKIG
QsYBrvFnpBtMwzs3Siqz5CMu9CojTyW/Y4eWhB7PHrQB2FHCcE4ps89ajj9VFRbumxvz7pFTD4X6
WBI7U3SjL8XiDr+NOATsbHR9euStIvUbkpnWwMUQUByuqSxAXmIMXkMBzMgE6cNYtt9rZVYxHQBt
D1uJU7CRQSZBhkAN+EzqHUQw6mXZ23b1Dldt+KdUCWrbPO83YN+BnG4lfWbxL8eqww0ZSzNjU9Qc
7wFqEKVfmxMnNuMvEat+mFWL+tuwtnV5V7tAOAlTQv0krdfxLH605w4rRsyFYZ7PLr5aWaZHsYgf
9xlb3YauSNhkH8qhXHhk3KVlNSEujgXjlhZBn0khpXgxskIaLbm6EhKvq6kIam3vsZNAzkWGkR4m
Mgc/8RwiBLoP72yUquc/j5TUfsHsAqUWBKVr2KNrCQWarGJxuuEp5JJkWa0eWnU3BOCC15WB3Vmr
Hf8XlYlAPl3CVKdRQFyf/PrxCRDhVZQXrIqfv+kuq4T/Vp1cSWYsVTSG0L1T0vgbw3AYpreQoYCW
XswZ52y/QrFCA0V0zo78MpxN8Wnjt4EALGQy87uvHYhn6VGJOv6J/ZVgzvRz33+G73f+GSWZ82lB
iwwMvhCihyEmRMq/mnbEitDNIl6nsH8wapX7VYMlQ6DJXFWplhrW0TGmKtGZRmJe+T1HOZFHQoMl
CznfHrMJKh9/bN0tlKmj9zZqraGPMRYo4MjVIcOzIqhCUrN3g3A5BSnYVQzKT9Qkr94FVvOiiWYV
yOtCoRGArlLoqTsV8uJUb233U7nK8GZYnkLjmCrNXiWqLwjhmC5LeFSaUYMAtepCSx9y7V3tKK5e
Fyc8surlbPCY+4T2PmK7ANxAOR1mdjzzOxxMjQHIaDbXOUDvRccSRdob7YFSAZIoCqO/+Vr+KIzb
O2GYT99858buZTdCVXexCq6fiwCNw+iHi2DW1FTTX1azHx4kZT7CmSfzPsGBETz/yhEjnNQG78a0
eDMvqSjVp29mK7+CO7kCgpOp4/280AAlBct7+uCeHzzUN5I4rau7N/PZ4w0gjPIdVn8BHoHfuHp8
ww1P96yAAuyUEj7QyYQ6aXFnLc0LyNuhMXwNGl5skPYU6NA+42ZWK5let4sEgcoeIc5syfYBiFFS
rq8hzw8w4+YMU+7Pm2SMM+HM4VlPjPf1atsnxntSFIajCE4Jf9aWLJk7c6UIrin89plrHuptrXpo
z8DmRMf2y5YKyLY2VC6yqZrad0cMsDqTZmIBd0rsUuEEeL29aMfYXIxdBKmsIMX0W88ve0SLiCDB
RobFOK+p7VYSab/bWoD+iwrzIaGcz6at0M8p71t8dslWmNfKb2EdbG2nxqlI1whBqXer05jaUc0m
KF6yZ+WZQBsQqwwhx3pJ/pcPMYLhICpUqw5s+HdOdT0f+BjK2yQ/RwNKEtysvEX+s8RVKEJBD96U
O+9tf6KMBVXCPVF7nxj4pWPg5tYTaLjY5AyX23M6Q3dVVXh4sUgE4BztBjgkvH8hT0WxQBswessQ
m4ziHqoZXOf//WbLoGJBLAw/2IJ8W1yrrx+RrmZwaksYg4PNCqQqK9x72R6wIqeRa5jXyN6WeK3G
xcxnsx7E7Ni16f3NSY3CvKw1QMOhV//bq5/EmWaZ8ZX8eC9M6IHjl50+QDDE+2ldMUndEly188RL
yStUu23ewxwOgAjP9e28jcqH7iTID3ppaqoSHZ3ZLpqHEG9uw4mM5iwCZFokXK7A7scv8+wjffvv
/2Qtk1McKMMFuvdgUCue7x+Gk6WCDL48U29RIzikBbss91b8YIrgE5OQbX0NnVLrOt50lpz8DC5p
n9SE6OdTkf96KqZcae1sX+hQWXG5lrnVui48f7z1s7hYFh/H2nWZakhC0M8HpR7M49B+4UNznWAx
9VYLqWfTbpjGLo7eaqM1zuOBA53ajD8/CPjaMRaMzSl56vBN8A4sXdap8esN6sRb9/GfWvbF4D4j
GBzUugRIn6jyjH6qmTdeXMakUDM4oTTdzky4c3i3+15cdcBE6YXmtqzzBCiTWrbklwdRbSr/CacU
N9ARicYjY+/DO2dQ8eVlWTArJ5ijudu5dD8nqpRtHUWe380UHf7mt9PHolrILrt/mEUhquoLGYyl
ezDhO0N8iihMNSWDMztlwIMhBeISyr/90spO7VeKPkRmsLO00/AYmW+kUFOCGrmiwhFaNqnaVh2v
fyhQ0Yayq9fDh/H2ITn5iJly9gWcugzg/+Ns8nglhwIzUMW/8nhQAFBiNm5xz/Vru4qVK5HKTQAr
fn4XSl/Vc1nd9s13RDGs6dqf6FwRRM+0wO4Zcik+WoxxOkgMShPAMdag3DNOYl4llPHGfphz/dmj
92Of5gKFtuOJLDftmmd46v2W1j8MQW7UMpjJvqUQOv9GcDynhNNXDOhbVLgxiAasY84lPhIJL3Fi
cOyJnmC8gAQyar+6e2L9mUlvvq8NhfDn3GKLYBWw21BEDTkZU8nNdcVCF0eG+zDZZWVuvZEMZLJY
wrHgjCVEESN3tqSk6oLPjm4cO7uRHm78qaPUDYYEHrNdGgtOLgdR9Vo/pdOhbKW+GWiSxGkQNIs8
vLEc0XdUXNxXPTGuMLUlxnAUo7DvfI9czhy1/9BhlK6HEggc+dLYIq29NkDzUwpjlSoeLuFOak3A
BoHS7crL6OEBVkZfz7jsG+WYAOONFCN3ud4uDEv1O3Bekmn4GX0IKfaslF3PmBNaHm48S7XcjaSk
bY/ysdyR5B5kv58Rmb+p3K8j3ZLx0Y/XWnB5tyCOpEQHWdeYTg6uG8B5tbrfLfuF8dvCjuwrc+Y0
pNBDsOAtRMLIH8o4jbmA43C33UlRF4yHQewzQT/xq55KmLpWkVd9SIyeBb+gM+MiVLibsLlOwK5S
2cyNAfamLFJ/C7zWRso+zjgyK4iC9YN1TcXDCLCo+2VVVVNKmFOK5hS1/l9mhe/8DRss50yRaJqI
BJ6fJTgEWOIM9ekWM9m+Hpmjfa40YJAFOzf933W8EWDFuQY32zp+TdgcPwtOfEcnX1r17SCwdiNe
4hA/J8TWhvU6EmXfa1LTEg+qxpiQd00/ZZzblPyo+NnUaBV3B2ggDid4zpQEBWTcsmoo1zGQTmk+
CHlgdhDx8IvKWnIoU9lb3yuF9b4LqWzclsy6lav1wzCxraIlwRUX+rhv4XBcadD4gpa5UJMZHIGd
5fIqkgVI2Y9G+OCLnMQDl1mEKtHzzU2lUjd8LH1O4zpkuvIroIufm0lliRGZYist8S61oHLAX+S9
mOE/igKfpKH8vxuTaPslogmooI8BAtRBrzDempQ1U2h17s+ynj5EwMfsRAAk2W8e1qGBtkG3iJ+T
ftPOamAmJb86UxykaJCXIrOGoZ9gGGUz0iU4RcV40FOKy48ZFDkHvQgSvL/n8BfOA8oLUeIY0Laq
/4uoDeVkJ9EjvUnIR/xY8qNFWDt9tWDygnt5cie3ED0gpUxRU3Y9IWFlJPCJqvf//qnOLvYATD1s
vaZfaZs8geM9HH+pm5A4Y394/+N9oSKK1Z2tSpvKcqhHW7MxuaW9tkmgdmkNp52ftLzicW/cYZtJ
nhguRsw5kfa01Ug5LwnxMwTnzNprQH15qBP7B6+KMG3QkJIG3OF2jgLPYvESDARSqCVmuDCYjKXO
RmevYTb9Z54X1GmpMkFc8uzYKM3mTD136uV+h+OI3VujJrfaV6jm2VgKbbUbcpVMaDqTKjqH/AmI
WrEFiIjyfK9HkaGhIHLJCc8V7tl0q6OSJEKPUBM45WNmC/5z+FnkAV6RjfhoJIVfkxG5Id2YrXke
ACyrYvo4R2K06B4yfNfuXWOvRcNj6fM83yIj/0d8uOvTjlRPESw9LmjkUWrYfa8lLk7Pc379hn+g
ldqpqs80fGifH7BgIICGCqn+sH2JQB9v3l0gXNAhpaxV0Z5Kapmo6YFWqugv184Op3/PwHPkmeCn
lx6hutH9/PsDlmp9QjvLOyQL0ARIv5qm9xcL3cH5wfgoOvNqKqHkDE7MfhAVTR/bi/naPSKg7sWc
74OzW+zwYW/nb74UtlJ0gv60cV6vSZfXMyI3ZBNDX+/WKCx437pLEPvHyLT/Doc+Hhvr8rM8qrbh
SgrxVM6R8z/70Xg5xXFUHPdrx3wnQ+iEoYnSwtM4XbnVwW4pAZU7VKiXpMH8QXWNzODlH2RV5tc6
kewASFfJl1rG0woWTTqqBCr3XYwuqh2RVVXGWi3w1Ik4DwX9oDwFJNfB5BMVpp8ZjHwSDBjNV8zk
4EGFrhjvF+LMAWrO6mXVOInFL2p8PnZCIE5MRO+OzoOpn9ts40hiJkiGISm1o4BCajk7sr6V3afn
P2Ff8gWfLgsw+b4Q/aK8yRYwFJz02ofPI6BXDRhT+GlBsMw9D9RNKgVNI1sFcEM7O9sujOLQ5RQf
u2Z+dycCDbXqpOYhq56ZQHMpgmXxe1n9mYhiPz3AmIr9MlghC26CdyhaEjqrkBGmbGm+TBpWLc4m
bECglnTkAmv+5qEF22P32YHOtfop+i6YuRHqjfaW10NiVig4a0pl54P8l1O+f+h/WiujJg6gnagv
YYKPADCEHvDbmR0Tl292NjxSyk6j/FGZX6oxPSfj8P8PHJ/3+imtwFuLHmxOlSFN4g5u6aoMRJgZ
3QXx88A5rZZcjx1oUUJ0RIGz0h1L8cwwddDGFebOCa/WXXtDG8+TlHzq6beAah/BA0vgsEP0daUM
1hMXuyE6RhiVtO8ibTcJyyqe5lgTMZJWgpBrDO+1DWSQGyXq9UdakFjxwzEdtbxNf+SomNL+mNtf
D1Dsjc2/zBt19oOR1jSufAaoHcQDaaasT3i/YlzG75hjTDz7weSE8Uh+FJkZH8aFM1kFabuPET52
OElLItBd+RHK9kVzbxy/xLV57vwh7EOCqPy5IthugTrTK1uSR6024EsWSjkZ9MlS8ZL623MoKiyc
Se4Tkjy5rLMe/Ux7OYSMw4Yb7oTFWygg56liVUq+qPrjyQSPTIFj1nplr65YfYlIZQFc6gXYxWH2
cBmTmaYodS9LfeoXUPkZcnGqxxTXuwCna/6a43r/MXqr+gX7KdaUNZrnIxaleNJLQSlBBpIfSbpf
j4dn9Ztutq/MYLGaPsghdOg6n6vMTEDUE7kd61eEyO7fuy8gjo/RYiOx5Lo2vKH5HahexydEn92z
VDbXeAR0p+RCCSqu5Vy6VdS/JDXJzr0wBLdH/MUNFmzNAnT990eP0M3nXK0ITFTKyc3q8BUY/eUd
fQDVym0oqRtTJUbzKNW+V/sG+tMrDnAVuee8BiHR2BEx7jiXV3O+Gn/qCKyt8Hnq25RzouXrcgNJ
Y8cjUuka0/Y8dxJR3/CPWOFEheEglH35z22w7/lF3Zh0HVPVOLYhcL+xbmgRRWMfjw+YESFkQXUK
c6rAnAuVbj6HZFoHLPWDZzPoNmzpLBOynotGmCDiEMau68GxsxQXZ5gRppX2EAXyUeH1s2ty38a8
jcG0S/lMZZWBzdsXbq3JIILVkHQ6RypW5bqdXdGtgrsdYiXWyErF3qpHH+X81RP85uxYgkW02ya1
dwadWx/IDHzRrJnezNTJBZPy64JM2wT+Ad/0OJhaAeHjDUDmrUyIrLc9CghW7pWa0LSWYLSbGsBW
B8mP9WtThy4HGYqCghb6XZ+FQXA3EGXnIVoOZXKSe0gv1sv4KYaZH1BQdeyR5ztEGVNoqciByUns
zL7I5Q6NCubZ1mXojqbcEOZwOfoTe/63brCq/LKTsYNIsYb61tDsZSuOeDgi1429XKfAYiITUCEM
fUQ5qWZViKuNjIHKVk5U1Zxi7HR2Gw9LNgvJ9J9WmJnuQxg8zzp2PbESbhAWgCgnKftXmSmmjs+J
MSj/FCzv+7c/Hi5w3jhO272dXEUFiMP5HIVulesyfGqRrnelzb8yjBlaQ1rfK+5hlRJ5+7YSDojo
qNB0GLHdUhqTfUEuk4XJ6vgarpxuyeU7GEoGJX8PLaBwPe9ZoDhQwqRwmtFqp520cAh8u/gmdZSu
8SxtvQkl9Yu5+N4TJQjCl1dX3JHpNIOxrCwwopWybOiFUXfyuejVWIF2nYMcgkcbxeUsoQzpi17l
c/g8S2pCf9zuyh6qaO8R/r9f/RaKu2Q2FWGDvzq8M2P4BDRmDMuSfRsEcLOU8jYHtTlqoMzqluag
mEa2OTxcdRhMeANgxRi6g+aTbco0e/iRsFfCfPE/Sr7maCswSLc5qz1slC6OBb3bL0BCJpAzzft1
O8wFCAOYXIAUPoYmpMHbqJte0Jmyk2+XbGc4rC8KSqsG/gH0pnwhiiFVy7jmB/Yc07LwQWFNeUBP
x+MXvX9DtjfXDbxhu6sQq0OorJCXCkuDzuDi00bAoGPDVpAlXXzn92rJ72UoiSg2hK8SDympVKux
ZS20ZtZtS3XJ4gTFUfY+MdCk+qWtzlf8fI5/J4dmZOz2/Bg2VnMSkPa0Bzgh35G63qIKdOwrPB1L
tQv1tXVb+dyIKY30NC5WTwm7EU4qKvhGmUsOx9ABEvmc76NSIRU8Lo+RI8u/FKVIN6Oe/p6kkpTt
lSKSYUywa+wWv9EbSQLK7R91UamfUCYHtmCJDWDWKNfQqbbAxTS/BoUVA/ewZ6ix/TjwSs8q907i
C9bZjkmyW83uVMP2rSg82RgEvRhQLdA/0172HK/y3QB7Xa1c4FGE9S5q8oFI+X8GRPm8zh2u3N69
YCWNOdk5fIWAk6dgYQbqf98TaSJhcHbx9RQY9g5gmBaIBQ6Ph3zTBudsbjK1ayd0DQW7mQuo+jKd
ENAOkATWRoFunOXMeCI7a/GBSf7h9hqsoL55yISIr6ZPY4mQafAAOjrAB7qkXtaESTUTRtOPrZOU
AhFPKWD45AcqdArkhVQklED1FuZqMkbU3I3i3o883XZPBs/emHWRdUaKf7HsFR1QjwY+hlIUNhat
8uoT8tqnBV77BGLNiSG5m2T8SULg2NQ8jpRpatqw4dK+z9AXM0AhLsZ7VHD+IoSLT903XVo9nvBq
AVRQgcpRpApXD/FH+1fFq+Tn36IgyxH2MlRkwGN8pERe9oXgaR5HrCf+NSi4waRciGJZzdy4rWUd
z7mCNP+q7sOuEy+v347VkVf0tKse+8Whtq3oC78B81yPFe7Lbtvr1s+2DfVuA44sx45WHioR1u+X
iYRYOohr/Ap9XUl/ZKHw2yg5e+uYR/iFXiOpGdK3dwCNpfgAnD7jZAK2V1LJBn3FuldXuhB3XTq7
Wpp08C17iadXKzz+TppqwbDdZmxJgUQoWp1s9pKn8jUDZyarTID85mTquLoUY+Ulif7AVK6+nNT8
PdWcRYl0YYCJBU7cbhDm1syRBejz46pt8hic4DkoMTbAUaeD93ySXqh36ig1rtDa8oX4dd553rS5
EdfSvBTRUPXo1lmdTm3wHo3wAtL2v59VgVBqNB7/c2XTbFsLbPXiSAdTzjPZ7HBq08qQASPMbhLg
RPcjeOejTkEKoBkYGf08n2cETudUE90IvekxqUowIMlG7m9Q6CSfWqctkr4SNqQ0t+xkE9Cr63wv
Tk04TZKXCufNDFn6ASB4T/BMFXsdQzZyvzC/kxpfRXoq6A3clzQToWJCE8D6gEGbWYoHECdk6AUc
m/ez/pZ4e1Xw7nWM/wBhDwKPzSi2E50ethRcyzEpnWdRaCB51xZMX0JLUlnm97I29aFTmrzq9LmN
mqnN8E9xGdmyRFrNf75Ha9Z5kuyDH/Pm22HlkkYeVDVexBmuHhkE5BZedgpdyt0kS3XAJIQiKVzW
vO7vP6RCwm5Rr67MfUg6G5Xxn0NW2FsfxpzMUEKPlttxr3oNhRAHj6jhHNKkAhcYkvCXgkZusr0K
rgrPA8AgHdJcVWpG0AtKp+5W4Mt/F73qe+u1tJdRY/e7HV8e18E1TKXB0/IE//2pBDo7VcW2o+BG
OPHKWW9qf7n4GUYw9b3lSxvt0+FilyXs60DxMEMoNosw42ymhr30g1pyZq5VY0gSl6j4R9ffxDXr
rLUTmmLg2MYV0OB4PcCpWnLjw81t/14+WZJEXb9hA3A5IUXlMe3CgDvsi/X0YLpEvXJzPgY3XEdJ
i/9bxgM0PL4J1i19lP8q/zbZ6bbDvk1l7LjcKWUxXSwaOv4NGoj0pYFs1j+oCxizVHZM5L7Kc0lv
5CcrU+ezMdcCxz9D9smWMk7a1YVlmKMCZnd9thj5lxrPh6rmX7IArjajIfHACYh6Hr6hUVKAkHGv
XPvYZ8BOYgHD8SSb6rRJYvbNaF9bCff84WhZqlOv/qtmHtiMBboMlG4zbCXu1lGYK94ySp0WBTJa
i5Q5rOr+2n9yPJvxDDXvDQ683zAqUCZmEkJXqAngn+w7GyrBiYF7HTK6U/047GLnSrZx0mb5bymf
jvsqxAXlBe0AngArlz1qPkce/ZqQKFFKa6D38CE1NYeMQfm36T/9hW3g94+SzfBBLC2sUFwTchNR
ft6hW2h7zl0VtCPo/tr3KXh+EM+pjwOHBWPZNUmmmX3+SXjqbIXfo1ar+t8H9RocYToK8sA5TsIE
SGwWy/g+NZg21JJdmvNBhwEBrAtiyThCiOqBw71dpFeNZMulHMJLq0LqH0Kp/f8vnnZytP4p7Tnh
FS8NK2PSC4CjbjYHs8J3SXmpNY967vX5mAsDAlxTTlAGgyb5cAvS87OT9ieARIsrDU/5J/wIZRgl
IRaGQ33xrEEo8hN6XqEN81WDtyr2ey/srsDfMDRt4bKxGsFxS+u01j017WKiHBdeICk9wVZddjln
IBYZyTp+4DnBg2bY1YYxGZxoLLaHd+VPJMe49fcDjwMOm8wb/HrptH41xLft5Q5FRKHTVm54fKUH
DzJSsZ9JooEY0EusaeV6J4FSmQ9Az5aqC97O3T9laquPP3GS79la5wZ1uT+mRrV0oO5fA8o9z4fn
crTbchreqUwLY3QzJ4lknA1BHL4CGbE3OuBtrSodjPOhtZAU9cYRFJP3kKBWfHj+GazHrVuKdI7S
k/xxnvyAzVFEyZznoSyCYhxCBixcIyMTZe2oDlO4/KmzJvs5yFxjR58wClS8hBBNJ5SM1VZnIX2b
4uSl/VkpHrPq87jeOuVlxDJQSR7ZB5xE/fjvlV2RztsVvbW2U7cNvSBAq817tlPoOxPBbVEt7MeK
iqRb0J/Lpjmjn/214H0QPlfB0M4mKz3WqpfNMzZvPIG+R387YJm0881L4+ziEKq4e/U601npbe98
tbwzh5odIjLw2ZuCpaXTlMJiIQSofQ46jmyq8OZJq4mcL3eIfWz2rAda0wRpJtAoMfuFv09JllBW
ZOYNPgez0Aq5uv32SjBFKECXOaUftnMa2L9I9kWDLfBR7gJ2HzD5WKb9kMpdbhoDidL2pAA2y2hg
lBct/7veKrlK0zFVZQ1W2E1ZprqIaFuUydxCaAcNbNdvJlfhCB+0fLIQvawBTtcVupFPS8+1dZls
lSrlMRn0rnGMMmP7hpn6/jOgD7au/HYfs3LM2EVlxfNh37WjMd0S8G9v2HqOX2jnc/yUg9308Le0
0B6b8adJWYeaFjcDK1qK+jKLB2AxUBqPx/Fdu7MzWiBn2Vck8o36Kn1WRpc6ehtoEQldVHu+iqYW
MZHF5eHvgZ1lS30emKEOrvykDJA03EIKuws72snLf/b53umC9wb8Fykv7sP5DFNYqNU119/Efxf2
we9xS9Cpd9qDNgNcn707rEW5W0zjYMcpZeep9aX65TBAXC3CFrih9700JJ+cw90JDv97EHjUaphx
x7+2DvOFzkeD9bHGF8zGvRtmKamr/l1j+vvzVtW1gF6N+RkNvRLMoFDvbKHT9ft/8nFf6pDTuQF0
PzPzc5nT1lEB1vwhbcPdfk+Z7qPhVxbPydc06ydNsdL857cIGeAyWOq3iiNATAExBv+B+ae3eGU/
Cvqz1N5rB8Kva33PzzHRcEPV0eJlyT8xTjUEQeU7PiNepIWIrnhgyBZ8xGmefzHlBB/bhWhgt8uR
0FsLNwj4uOI6qPWlX+11mAU+Ynyjk5JpILqDJvmdcSwI0KSlfSBERRroZcfDZBBIPJD91N8cPEMx
1hK9mix622NwvnQTSL8aepTgrceQvqN7vwgiCuiC1hiS5o312L7gV8YuGrhzQ4rcBNGwuDjD4Bfq
I4CYl/VYyuD7453DYqdLYH//9+srrCt2nN7g7pC5d/VClHz2JTpc3XlE90sLn+lECrblAf/HPF2W
ZCaPMDXVo8gdZJtAQe6VHw+ZrVI2w3CxCR3sYBvR2DBeh/X3ELHLZRUXvYrErexTzhrDLKw0+9Yv
O1lewL9HjcgZKirBDXPTIKTst28P0jTvkI3DNaPoEkNOTGBc6k9jKvNmLl/6VGPYctyR6ekxu4yK
OME7CLKkL4au812/xdvVsmKpmvGwCY2oxsJM5707Kx8WKjlUXD2iEqWAG1aTRBkvLAmmnbMAoOB/
3BstI0enwHLalpwPay3eToMzFymfPTkwi9LlnYs8OTxI+0A+xVKYzLA3V1nw2WnR2ip4xr8EGgUU
scC/eniR2TtOlqv7wrz9iGHAiF077j9+RrmH4rRgN/wXJ4i95ckBSAJvIqOYgeexr19DorZUlbBJ
3dNgmICZsxdpt03tEgOnOPBdSAAqK+yCVuis2dJEuak3MeqsPIbsWZDQzoLzFQjO1tV7ctEckOee
Lv2w1ih3puOoEWdymP1MuicqrJxKG48phUaghnC1azY0wsyzEXBh3L2wKuDrXXr+0Jlii/1ewRuI
5YzpGrd9RpIiRlSwLBLj5nAdSSeyoVoaCs5B26G71dzLbNZPNPXrlxpDVCk54fUWgmmrCMp7dEMY
7aOpQmiz5XinTyyVylTt3rPVAkXdQRTerdC3BGmDm8wKIi48pie9BG74Icw07hnr1TbeI/NgPZ7s
W6qEVk53I8iCP0mdOShrs3EN0sjptfHWOVZz/cfjkgw4qzHJERx9lJBv9B0IXoKwmOQDSs9B80Ni
Mb1WmFh9MIZpG+t+YdafxvD98bUM9KtxCf0PbzGDdOjzQAuuaqsnEUT37PjYX41KGQ1Ex/5soQoG
7yGsHEqB3mnC9IgD2gtGdeIXmFsdyvvR/H8BYkluKOVhxohnYnAZ8GlJCHE6BGs5+M7hZEdTYjPR
mBdbCOUwo7P6BHB8p6l/vRuqhg1gpHMQUYUNiAcicbunOi4QFH6yRKllSts26fWRHz/fnc8/VSps
5peo81JKvI1NqXy4n5WKAxrVgbLmYYJYTGWEJVXiqeBaVX6CJxHGyy+LJuamW031OaAbAaEEObz6
EZZVpqJYXalB7OjIUciLzNyAb/r4XiXPxU9VWN+KfaExKCANyFLrR/aVSGGJssgifquve8rVMUS2
iyrOqj9/QJzvxUkrfElnGnzvGuIcRLuZkvrFqUAkt0Rx5kIej218tLt7sd3qqXs6DPzT8ve9TcvZ
SuAladESCpWfzOAeTnBRqg/fhl1lNTyZQrSMotTvJimCCYccoKEcLlM1fCu/vqiNgZbeKf4Kbe34
OxtXAZaaB3yw46cP762juEOuFqXezyI3n7HuWQA78ERgAODsto8XP8f+izhxrlFFNjuQuRJ94nZB
0AnMZecR+ble1Am2EDMbE9Nu2bbm3cyo62wJ4XfXjT9Uz4IFMUttvoZAGr7gYI7me8vbjusnSN5V
+SXOTgwqccv0VsRa8YgPlYxf0BR85NuXl9CpPtjZHS9kr/Jo4zdkl8s8ZcMx5YANBKBMM5jOH0LA
2+BOOO8EbzKx6SsEiKXBS2zMy4pEm6XxkTnxSo9AXMLslq/kRUncehFM9pqK4QTfjJm3KlxQcbSF
zc3oR6ISAdo4JbDzyoffRJO2sJOEIHi/kszXLarW7ecafh0IxIS190aQMpavk1GBX3zQlQ6PxQCG
/pis/iN7Otc/hsaUI5JTVqnM6+EYrCwNi+xhtCNcPpdg7pKmChLgN4UwqjmvODTMOvFRIcPqdye9
gT5voVkdAtLMICeghr1wXSUozIcDCYsT26sNbk8Xrf/0N14z3X4//OeAKNzs6kcRduEr+lrNRuJW
uUq/vF8InD42mN9abJea+2PW3bHziztLu2pylB3pK6pNJv6/8tv9xKJ1sUhNNwv4C1sodq4mTpye
YOh/IUl0sZjYwK9MC5THswwrjG+CEJoAWkn0kr3mRqNekXsM+tjRat3TjX+L7iqAugxKsHgScKvj
D5R87WNWvc1JM99NvE+ZezMtQ77XG4jNb2EfeGghD4rZi9LWBN9VOcYJqL3ZRHh/1yGb4K/OWSYs
6IBX3m8M8scr17FSRsZXyCvJlDs394iodCc3nS0In4kj+Mfy8aC9P/SWPkG+IUcDWVjXcNKunDLx
8E7acyFTXmJ7BpF1xd+XxVSH2qhYccNNAcHBys3pVXBldbX2blhHkjvlBx7oO6HY5J4wkezGE7V0
zZ0BMZlsUedP6jpE2c9686aHn3G5SXwoixmpd0Ai2HQDAlbCB36mebIZrzqipVd5vKcGb9psFddh
3F2BCUB52FCvwKUck1UGVML+Qazey+Hlt4aD5j31CN4YGEZrAbuLxzxNgyMImPznCG69Uksd+2sj
93BjMpUTjlQoKViKmO4LD9DS0sR1d6zi2ybYYUEIDtoGpMSnrORqv7+q7974aX7+YAjl/cPLwZpS
vMBcEi5/v85o+GvqgjTxT/4nmUl8iLvN/jTZY2Oc43D3ewIODMRgCzaXJkuI4PzLNBLD/m9E2S//
gWTHwi7ayi9D+YkjB36t9PFWAaG47ULlWdgZpP4FQ/fPrZwsaVi2ikCMAVfVn+O6UAuALUHwWyr3
6khBTEkzJEZTOTeiMQAd/XY1Bl4lGRbghZ8KB31dBKpXwONt3DXlNSxjWwHY58m38FD5PyhSlGEg
Ce/F83a+iBYbVRjnZ9MeeAhk7uu9U+Mhv5Qptjmtn4f8VgNv5mRq6JjpvM27ItU/dg8WoMHRbfr0
DaNwmoactjp4E0XW75Ooon2fZyw0A86+XjIIvIYiztQ8uvCVqD0mVxlCp57T82/meA6LDJ6BHSaS
NobgNMkb8wB08L6AW/lpeWuil+zt+C72Ijqmuv/+yHNyUYz+kYj3YQxdKg/ZDmCZHCj1KOy1WYb+
m0g4/mjqA9A3ZOZautjSFlhh7vRT/n4odNR5ActR4YDuuaLwjbP+tCrCmuGjy4IsjutvzqP9NIY6
1S1lr2cT+aW5mlCUWwOxmjHCdcyHLYZLUXSCYkMV7g2u5CeufBsfJyDDI13wY/GLYfXBWxrl+9vT
tjK4PjPbs+3JkcJSGRUfidT4mczI0OpaDeD7zmgkNMlOt2mJrphA5QsLJTYK/lsCY/tXHsucWfyJ
IQFIoW9iZpDEJJTRBj5AdBoPOqeyKx0ItlXIVUBxGFkGsmm8wfVM8nyN0RAJFeJfnKpqlbCeUvS/
woSc8bIy9kWssMyy6w0iVAaFKTszFs1GTurxVqQSxEqDhAF8XYZEWl8YtpX+rMxblhpunZKivQJA
BYVmPRGXLpdbmoUGVULszdMpWcEJ36PtKcyvAtEImoyOx8U86/zEz3ilm240dHIkxjs8lIAEZHRx
xkvM26aXuZEur66St3JxY1swF3v7e5iN4MIZjRYDDRN3Y19RP/gPYPOEZhKVaSZ8bwDbZV3IyuWg
kk/rc/M4hC+fdGB8n5dKJrVpBKZmLmCbrNsy01ODXmWRrD3NvLriKvMhEg/E736D7yapZRlgB7ZP
AmYABa6T2HgDq19uaKffQZwpEekfPt4jetVyYrsxUYYb/gW9mCkXILiMh7SEqp59gHHEJWA3R4g6
X0C6v5nOsoEZR6eohM/O5e73WLTP17k8AmXC97cRPFSGqO9ryGn208Kxctpb4N6Eg+KzecHNgv46
ECzTnVU8PYiuSsLtA5F8vaMNqweEHjVQPymWcazoO+LCJvKgIJuBID2CFP+6JZXMeQABCA5TDaxk
BKvb/KKjW+gfqP2rFT09lQT1WIcSHB+ITwXUMBNYjLANtNMBPlkSBDISy7JeQ9k3q1d6XNEoTiBh
/yomvZE/hJyfMGYJygDejQlCa9N9F9opAYyGfKp0auS0vbFU2Ddp21LV5QmDAUwB/ncKwojTB43c
YwQKGlLFWrNvTyEVxAx5LOq716LQ5aGw8neNrTmolHq+ckcnydXA1LPD5w1bjboGnk1nY5+09m/h
luWbklnEZQX+C3WofxjzE+P5dfTfSriQBZflZYUk15AeiK3biZTOYf9Ke8WyHvWkeC/X3tMwI07m
xDcuY/7bj1jibhRE4ugQgKGrUaWNJ/8Bco531+1pCjXBLtzkTEO4dEjhX8zNFXzi2rrLOzPBdDhT
Fymk+JgyvswovLDPJ0OI4Io/hIwPXIUmlGd9zXF9WGw0MJ8bKZrd9WPdZipEaad3yAm3S6QHEac7
qP6sYaWnoQU7/QlQH0sOvnw4sQqMj/Y9bDNF180diFG48+bKJoByDS9z+ZJgfvn7dC8mDn6GdMRt
mooCqmWzx4JuzmJyJJqbVMnfOdk/wApt4q3+ylxhsnfDCIIx+z+IpZoHgvoecKd/zyRDU4KQDfL6
NQc2ofWzoRn1Mnwwvfost4kIi0wrcb74oM3GLslXORh9TvevooqCrTTqCvwmGHXZat75Hdgl08XI
C/8HzwGCjAj29jZRNrYmPu2Pv69XsIYIsGUieUwBI6+Q4nOeplHWmTcy/Sqg4tIjDSnGmJT6lLlh
qKfsJe+kKDeNatPLzNfj6aNb/MOaTEySQT7jZHZzo3CUyKqsTmAIfs3CI4f8KvCg1ZAKgFYVvMct
pk38CFzd0DHzILYZgrRsoK76X4WXuBzukDA8HNQ80PW0e4KQlPWmQs/D4FhYW+YcAkhTy/Nl9ZuY
2tUFllgVAZgNzZgHImb9bmxBAgkA7aZZF5N9pw0j3kgLD1AcDEj/+P2b/4/Bqn4SyFYo/+9321yn
lu3y5bPHdjneZSiOH4A+U5s5StYmG5x5JuFwecE5+whZx8VVwihaLyzHp6WHQ7Bw/c1lmGVFcJzo
YxzWmifQb0CzMhbzsF7UimgnpLPBv6G/WexYwNhdsJqFR3LdUscUz3mYE1qdxREsOpgYbPjNhAfm
rGn8jp6SGTGvQJReles4tjWtZuQC46NL2xICl2topdQ36TUc+js7I6+8Bza03VMXri1AoCWlKp58
mcvWPaeXZnwVFxkDtMbG+2AGfDA/NjO5bQAx4nXeSFfuI3wBIp47niBNmAZhxSDNgiotaqxSukbo
gaQ2wDePqWGjB39HXGcZArEKPn62/MTPy86ck4xz94WY1tl+1m3Q0D9p49iEGC2Z+X7aTRc61+oM
srB4FnVhE/OXMsTEf0pNSwulH7WOa9QHm9dnMQjy2BTbsIJCrcw2QDbJO+t4t0Bvb4Ud/0OklYtS
DFm4qy/ZKx044uT+TKII4Z5q/CmB1ngTLo/4PjdvW2Ce7cF8XjSR9kfGNrd/P87jXMzN4HEy4ilr
PJXkDF7nRj9rc/yPhbT6k2CviZQAuTG+OtPITeML5f8vStvKqotHNoT37JxE24DGqCusy7eM/hiR
CQEv9EPOZodeTI/CHAyCWX0x253pNbvVnXO0OUB7xwQpLMDZb1h/NQVkxl/tzEIEeqtCLCVy0z+J
K8n8hYA7PZYWkZ3xro13uQXHJpBpivmoeicizpI5fuCplIvj9rMuD6DW+JmXGF5/DmO4iS7MgZ6d
iriTtgs1tEL3f8ryM1uWdeDSgAtTpWbNylfiymZGmew2PQ9lP1AyIeqC/wyQnHnnieuFVAW9bxZA
+/zVAsM0dhfLCHP0dKS28jVSFYYUAy1yKmVCV82qMBFXNg2KhcV9NW4YhRsHf4FW042Lu7aaYCEC
dpI32sQusOhgWWo7eDWH9U2LHPUzXHGhsYoF/bczfhnawOI6S2RAO0a6l4XIvwq3y+M5LAoT2w6s
NHUrn/O7XW87cRoMNAAy5QdApK0Ji8Ak5sOct9RnTXJhH1wxLbBSyM4HeDrcqlSkkN7hnBHHGHb0
4Bl+W+38YB+Mzm/ZiU+a95HLCne0R36zdmWq7GaXOVU1Cjc+wC22cqdckw/HFAha+t3bjArBWAVw
nByXWM0qV2W4ZSkhLxm0MfLnvPlSjsf66NLGKRH+weRNGqia7RsVJVce6IRaaPSqpI0/k/C04ujU
jnQI8v0dny21DDSqFVGYEg2nt+uDBZAssWSCVe6ImCCFCqzRW6pgeShNP8BCxLvOSqUArdnxSMMu
jvUu7iGnzG20JNF6zASynAl7guO3V32yEt/jeN9e5y2opkCK/h1zJ4FMPKB2ryfO3MAzSWdy2VEJ
j9utCg4ov+/0YXySXuBrzsUiMcn7O1cflKGszIRYJVbQY4eeCOaYpwvraBWMSEOIFEadZRFg7dFu
/kYtPtWUf1etJ7zMJGmA2Lx+x1u1oAN0NfOREZP2mSdTre6TDUFj0E4qum5OsT18fif0I/Yv18s6
ovTeuH7duDAg2A6TIxV+MsLxySgu3mo8Z5VKGq4UVs7aseuxIKo/me/SK+G0/R5E8ahdb9QoSoIF
6jIeh7CP4sbTGu+b0SWE38okRSjidzGUxfmAXe6sEUDaJkR2mZGO6pQYrqvBVnFQhojRLbU0gcps
6IShUnHCKpPk8GIOxaqFqZ8LvnwReQ9DzkLwM8Twf6Nm7pC5WJuSruKFhB7LH3K8KXz9qIRzfZdI
ynhmsdRogSp+KoyxHYH7pBM1hnXfCMNnNZfxnSS5BALzObjXWrXXum+sP3kB3rrJ23pi/LEFSmhd
BAhO+O89jhik06YHiSSRp0BybvRkc3IaEGt5Az78dI7D+9MSTzDSejPKmqASJGI2SOLv94+UZJAx
7RjyoeoZbx+JYy8RZ52xvcNfiEuAnMccmhnH6j/1aXUOPOvHOmAE61eYDswnwkhIDIO6Jh7uq9qq
ZWJv+Ylm/VEqDL2Ia71VMSrGnJ6opAS0po9DdXuI1X+2qeSX//KOPJanUyiG/bDVdYWCRb/tkoJh
kL8jAxU9ixs1q4kwp4Yl1GqP6BViCWSLra37vGlybCPlf0i1j+01EYh4MfZtKyirJ/T0ipjEproh
VeZShfqMIQACHM3KDMmbGhAiAiYyUfqF9AkAGDc8+Ab5oh1sXq8Ni91dSl1+ZU6JFgrYPe62PkJv
yBQdpgJ2NFcmvHX9dD2XU3tEAaPi+Uin7XE36w1BPiFQ9eZYATdzeq6cpGHbG/WswWMR17vYyUyf
yuNsgxaNQWPccA5xiOr9eDAX9s2kYtlcAtSKYSAGcXIAsTA7jmKmDys+F16mgM3qFpd4iOKDv/pL
KSuIKJkx0bTCtizvj2g3fbfDtUsF01gDIdm6ktvluoSU09NkqsMxo65X6jjcm8UHJKR6AQiwT7Kx
gdhZQnK6MKt3R6MtDs6hdDrHYsQVw2iGbVM40r7gcEJr2RmKHn/flpU+hZKS+eOObZa3CGZAk0UA
bPJ5v9nFlTCy/RmjSLnmN2wHMxlnsws98hafKFJ54EAv6ZYT+GFlTJx7NwwqzqKAjk1z7urKK8Eg
6pDhuMqYoT+I5v1oKXxjc+2eN98RlSpcupTPQgc4ucTpPQILdpWgr0MZJuoCD+xRq4Glf85rmQTK
UmW6bgN/TfYtJZXoo+u9Ebt45QxDlIj2/a7ESGjNFD9Vo3YoyCpqEZVSsVNdjPXF5G+cP604r70k
KaOEHz0tCzRA6exLuBFvA6ehTHeCdthtPYyDharlFKmaWpQSbSUarpxpUmv1VvXaLP35l9fvo5LV
jS7ECZ/Ng5cfSvqyaYiferpHZ/j5aU1CtB7aa1WDU9XoNbF4H/4dI16Ohk2POuwu/G/3WlJWrEmB
OurHBnyvrhOWBS6U7PRZV/lmJklJBOvz25p5a1nrztHNd8ZlsxtCKPbRx2qbozycqLbvhweaO3RT
/K3EA16w5I74Kx3Q7Kh+XCshLnWW13j2ZjigQn8+d5Wcs9STwTpe5kd4vXS+Y/4MaRHANFLR4gpo
RzClDzbiEYcEPXG/kmWgiR5gpY+/1OPWVxgj92ijcum91s3AtW9IxOgQPbSOVE0svKTtmx+gNgkC
s1UcSPWqHlsZeOwJcnOOOmQqhDD/ZuwcSawwVLgewtfCgkS/RZWrzFzHqxH/r8U/VJOU2uHppC49
m4QirHOSaokArqKYQOQ+LT+e4vsUHM3p483XeaiORQLwTEW/AAJEcPD2awEChrNgO5dxId+4GLpO
iompaTRqJ8KMvTFOa53Lq9QgJ/EyfPqwG6LABq3CkvZnFTd21fiduWlJb8tibS/ZymtsKZTYP3wU
k+yIU5GuYYnE42tfbMOC2g67dNQ3s7Dc/Hq1lcxH0Y/hSfeYrGuzKb2dbwc2UEyC2LTqikNfqHFV
k5/nLnGtExA6iCk59S0qAVm988VUfJIhtdmOEZ5e0sGx53ByAswcFxydT4srjnF1YfPwj7qskR1v
1Ys/Kl3N9DAA93ayomLyPHs1QLAUYYpaqbOOP0P0qW6ucXDtg/2R1RqCNXQojwmaR/QwKLA+YbzU
n4FwzzKpO09HDy+ZdfELaoIHiLTVZRq0LOD/HYZycMIJXOTinXQovtAPnSJe/e5NlJcT05BMj5b3
U7UVWSVR9/FvbSln8iccWzqlHutFzeJinWV2746zOGq9KDvNEiMnmlXZq+6tKvZxpWV3rnblFLa9
ReA1BIlDUTso/v/kx6d88YNozeBRfdpUTVPLMv1pXShXEsSYhwVWqGs9GJrrOuBDGCAR0U//wA1x
Oy1JvFbi/P0ZuyfdXzpKSegc/PyxnIWUOw5hGraWMjCuERlNQHSv5AtguCIdBYCfZ/BCPTtCtJTA
DkWWEvfgeAHQ006PjF4lJLf6e1ARvJFN8qj7MuZz0iVt+q2Xb1UMBEPgNhjYd4EoK5gifsVUPO5p
Wc75Sf4vLf30vxwC7utR607pgVm2UGR7GhAnYGoTqL5psEubGJ/+aBhzEhvAdY3ROPuRe9mOWy3Z
g3hld/czMTPQm8NRWpdypemwxKHNSk6t1adenAWOI2a/Yto0nfCIsK5Z/hpuXr2YM9f5Ne1e5K9u
xMiwJu4Cg1gcvhtG6EHmyhQ6Dl7fu1Z3xTIPK4fEOMj2kl0g8b/Lvd4AgXE0oY+e1ievb27DvjI2
2LF/Iv07ki0cTu0noZCTzin4zkdXMDIEDWt0KEVfehYeszB9vPwCvVplZGzUi4TEx8XeP+KC/Bs0
Uz5iwtGHkUamzOD/HnnETLXF4e1oAKWft4JMo6WYgTxOWZq38xaXhu4BhV1RjKh844TJsTJLsT1w
7Vgqj9NomOXshkHJULRpBrC4pq06KGONPEo0RFXSDSj8KQRQk8Dzrj8+/9HfLMZrOO9tE6Rtac5g
1VSksI6cmExWETHUVyy/vbKHPmmkmApTHuCEqJmMLPv6elDQO7/7yzY8cw4bCI/onnnn+gzfbq/p
su4G0cW+kIa5mCsswNiAqXLDtoG0rHxE83eyLo2zCLZuUrd9A2JvZHe+O4e4t0/BbVrAu2HYaA+6
tgeb/oBRsPyTDeA4rbZ2JXMcWt8ZO82IfQ05EuuI8gTfpnkyOC3vUlsu9hruvFF11pJ7RUfvXaBu
uladkyKitoDpHOYfI6lit/KTDD2vwfRopBwbIqkUk2B9mSGe/X9kJQODvx9d73UnDIMN5WPcPXnV
ggS65pZCbJDwUg/YJDaO6xP3nWj9/yf9KnnXjiFcEdntJ0W/kWEZw9Id/IGofNAjPKSrApdaVeqG
Ipf4LgJaWy6VBqDuZXB/wAM9litpyzk+Nk0/8amVyaskF6rBCMpxaaKzGlz9lZRvzPrUKQe7cwvN
9MQdev1bioVb2ICQPR2Tgg+YK1OExJxJo6G2U5cm1GXWxfZHkkwQ3buf+DONR3//YY3tSO6f0t/Y
hb37kuOf2ukB0oYA8SkDh8VQ0Wz4zx8V95KKtsGHUQX96VO9oQd6sRanaZEWUPzcV2M1JDD/cVnJ
Vi1gyOvXHDVLjzP5PkVdpUHw9ZzmKnlVQTBcNJcq7aN+9bACisuBF2iUBIbZgUz/TqLplxnVcskb
he30tRr3oi2M6g0VwN2c2F1ixBQzjxX0poHxl8qrCXcQKQ3EaVFqKbeMMt5XbVK38B5FDjCOQjeu
reiTxFuEz5vojeTRp7CfTFeDsBpPB2q400sAA4I5q1EPdHeQADrl+Gp4z5YfpdAd5Ip5gDpAz85U
XxZdE2ASEheTvk5uShgj0h9H3aJmN60laPw6zFgSybV0Y632MdJCr/SLsoPpJ80G8vUzXx2/ryh1
XqE6W5bNEOQVus9sI8o5gGsyyuiN0WlVP8YkWezoYIB0j42rx2m3lGruwE/KKi9gTWz9v7+JhW0Q
iQpshubLFk89lkpO/3rNTpjcQbhOufW4C5jELjPT+A5oiC0JDrkC87uuxUzAhTYim2qoAquNlCSv
XIavFxVebod9F/FOad8mtUaMm//8njkS4RU5Ugl3pjZ7h5Moe2zE65ptIyT+UKZ5+RfF9lAdkPk2
oyMMfAKv2XvqVXnP8XW0KzaXM9RYVAZYpocPmV8L1ExK/5glOMilHmiyPacE/1Lr0Pwb4JAU5hSB
UzGKNPn59R5ZB4jS4K4T/VXPbC8kfvbamRuGaVxr5NzLnUZWo6EG3Kaa2Vxa5sr4ooXflWPN2aOy
WrLO8Xo1WYhM3WZBPNmaM3oZlgReKqrgwqYZRpOalmqET0t7XxPn+ve4nXLPBQXuwMv/coMwpno4
oXHV6/7wRy8EZM2gBUcTFu+dhePuI1YIctcKmV82qM/5PsEeQ7wai7LmII3Ns4mKU8CC04vwoBDO
7LeYs5YrBQBHUhl5TWcg0WDVkm23MhXOFyioPuhm/+XIrqQ6JhKDlXHUvqrOPw24Pb3PVq4uqZ3q
+pShH59mPVIwaRmzvRrnqcdxll7CMHHxDl7N94cGzfqCmBvNrt3MhmVJwR0Z+gGE1aHU+mjUhWly
7ys5N9YpP+kiJpQK2OvC4jN9HdiyMHql8f89FYd1jJcUsh9Zud5HQ4KoE0dKVT5HTcWcI4/4DBVr
pKMo+yrPfs/M7hj1KEzjaKRQuENlnLB5K3eqAJtVPDArPhCVrFLb9BVQH/FRFLcRBps3KwWOZbPr
1JLrSfTZ0b9v8oI2uc6F3c0l0tuTcG9CeT6DKcDg2iVIH6HLu5ypWhcYXa78jV8y64hE3q6QeF52
niDlJsY1Mu5/Rb0r/HGAdy4R6AVWXgmdGu3bCCJOdihalT4G4IFzRPOPk0DgPP+KOnEzk/R5Pf+L
AKSIaz4+q8DtRS9fIG+EWrdk1Uf5LK9Od6/L6sb1JFImYUu61aEwg5ILjfego79RfLpaZ9/E7yLR
+bGeb7abqVsgsJsRlBceki+Yt2jCH5Gonil7eCjR13pDuC6Mjr/MOm2ZY5+Iej6MTGJca1ym78eu
n8uL9a5Q068qq6Hs/yZfaOG5vQWHSSlpSGJ0RrYd2GcSP4slDjvm6+AevEeCf9hhWAVM0ie/UT+F
//H+PjL4+BKvMX0hB9NdnJZ5vT96SLRzz613Jqb6En1Q68fochRsHMUPbEvg6/y55YPHRwRPKvPI
vpIONzIy+sqlk/E6yk7v/aLzBvKeaipaWKQM3A02nDCjJV5yyZw0mGyv+hG1fCdz+CuArrggSqJM
mUNxmkLKkF/YRrhDxlHIfqE1m9OlvXLbKboQLtMZz43Bf9baI6gf9ZhzFxkrBifT2F9uibCQMi9w
zk3Jw3nftHIAbmfA76IlZ3nC/31SXAbbFAdVdZSqctG3UE0BBNxmHymwPzpHeJc6QyejqFaapce/
2p0gNWdqKm5Cedctuh3QmSbVKvBgFdijZmbm0MleAf7IsWR0O3p58KpeeKrqQJUi5+lgs2iYEqZu
rjZSb5vLAlq1Zbi9RzaSTI+wFDSEfcVVBPrqxUGQRS8dEmSHOTDayQedofESAFLLXJU/Tki1EHFh
RmFSGjmUfJ64CsuS7otvL2yuUM4WLRD5Lfy1hVBYJy7k6joy5yw4LYmUKmG/794q5jtkz+gByrDq
EA/qoEYf6j1Qn4x23GU/iXOszGAIzWQ29x3YIUDpsxMAlvga4NQckmkq81NcJdEXPSWYw28UzAe7
SDd5x50jlrmUyjcMskh0KdNlcFf+Feu58dgSQsyz5SJfKiXCZS/ZbQjmZHQ9TjSjXQ7/q9yh0/H7
CDZb9lkbjfclG4p2napcgTLjt9hjU68xtYMMj1vPxtVFmMbpDEbvLixSGU+y6I85sg2ffWt0GbH4
ditsr+xTzxi4Ac//lvxBd7X70CLZcW2YsuYkVsWSI17itvFcAfxc/JeRhHUF1vPP7yJ8sbiIMpRE
KdsTW5LADcuynan0iDHXiPo/KC02LTEX5VbJ+WZSQkqCo8/zAgHguyjoPjayU6NVG8CLyCdWS/eP
QJjkrgXAVPnk/uDEKgtqjdhz38ET+SNgWrGacWYGjKGS9kqvSHwFkSymYCucilwZq1R/ABy9SQe1
dFk4b8ulS+wQu9yPe20eWJCOlM6wM5gIeH4T5Z1qHFLMWdQEEatE76ChY7E1cM1SIw1TpBFF0gdn
fjkbnPlw7JLA92YeAPBvaQzoXsca8IpCN03y9gJ5zIjEZNlbZ+MUwFyXAEPs/P2yAd6hLCpWzGq8
wdIrthFugm4OIPdKUpBnbLkGi1rrF5VCG03dFwUM36IST2DdRImIknRR1O/rc0QV296dVuV7breY
ekZgyv5KVj1i5Zn0V0ESlD69xdmoocOORwnzGgcqF05yBJY9qH35/QZHoJ2Q+vuPUrnHWldYt6Mp
KnxBaq8TGAO9XACB4IDkhHrxPswAoW2QIS77WZil1xxTFgKgMO0o9Caxbui6RCHoQiT8dAwy5F5D
Mj65qX15dL28MDiyeiXvbX1IRg0FE7ziiVpIsYjoBevA+9ubOo09QXfXonajryh55lX/Yvpkjpf8
0wV06sZtUouPVYNtgQQrQyjbv0VvWoySJF0H+RPSWpKwTf9tDtNsgCRUH93+uOgiRcix2VxYojm7
AGUqmDLXdOIww7rU1tYY2S74IQLgKkwlmg7z+vZUdDjkul1ao9/ucwz1FV6BT8obreg2vYFoPA2a
SIiJpfWRzkB96f9B6OnobiJ97oT0xwillbvtyHpKH/qM6axZULyWLtmm0BdmWuJTqpLOG69oZynS
/QP7hrhWQyHKpk0EbqwSmbSywQthHIolgfEjRwFbMkmfwOnEPphdvtEVa7HCBzL9pOLTXupF17VX
uHEZl5RLRXyloSYGOcxuTG8wCQXefUKKJgGIt6GlUgSb2SzsbGXO0TSuvOIysQZBIGlntGbivP7p
uyzpF0c6cva5wnWbfXG9VambBwCosOptd44SoGiYJtDVqPhtYp4DsXcdODx/DeRhFqxZ11pUd3OI
ioAM61IrqmBkjSYh2ut0KkZyPDRDmkYRqA2CdXI06SNY9UTygK2vEkE6bfom9eUeWZ797wWooxnx
iN2EglqKy/EmIGXCsx8//5Gmh/zkLUtvZKr0NTa2iSliZCLKf2+7gphM6vz0oTyTogGk0Ymb0qhh
uz1lM9FnhhJDXuZDWIy43cPnocX4ZVTVIlzOP2kGXkdPAhLi29zCHksZJOcxKLZh1+/lWg4Ll4UZ
0incAn3mGg3zQzxei3R2qO3jPTzBcq3nqa/wpYTlzlsVcDiLrrugcCqtyVBy2nl8TLLpUk7h5kMS
pDBtAVyTay+EPxGQNdXETHRxBKohXcD1+DrXgvqUnnU0eGdT2Og973ieR9OM7LTRyTP8wlqVroxW
wKJDfC7y9Z5nSsKBVn9yDdEfPj+UJt6FQl90UhACklqyrPXp09HOff+D6yWgFYxN/CCkLbiC479A
qPuEqbcEUpdMwpatvqfcLmTCBgyzzad0Sb07gJIhT3j6nZxEMzEJlEwPFRFAumO/oX2pMr12Q1FI
zW6ZQbkNHPxPXiYh1JpBDJ0jH/SVcqc36R7DjXGPyHhHkx3H1iUZjVkmLEoTuphDouwbHmZ0GuW3
Dys4vtl0yb4+NvBonRwjb/kHFm5v/5o6CWCwG1bsDcaNVTEAgVucDhAvBF1L1s4ywfczQ9DbbqZH
fqtZyNQjSrC3v4+QmyJEHwDvtctMxOUq8qLfZgYKX3o9bFFS77SKc8dnXMQfkQ4+zmnxsVyIwOzk
lQgaJta+HCR6EFLshV2R2NLzyhfh1KZ5tmOEEhFcjQsYf3RywW6dwC2VuRewcIooHSe2a/49bM39
WgzfWhSGe/KWtTGi8vYqsD683XyiELfbSb2bTKzqlgs9Zo2FNZ2K0XNbF5tIdrRimSJgKH3PIk0o
Afwr8HEFqlH9enYeH/Vpg94AHRESBuIWC21M1uhzQAWxSR1d40nfGXDQZMOVIU2Ylnqzn+HZvDH9
lLZuL0XglcdiMF+b+GtrbqKOMj3OFFd/xgZyiDtg7HZH0kwstXL4ARRvBzOMLnKmQFCu5hMeKYu1
eSr8P5kADpnS+TaFw83mrRUQFISL5ovbgFkJxjelAxzFlxAQGGAX9iLK/eAQBw5l3V7XYS9UyvVM
335EkeIOvwwZZblGJaqWSzgHNji7cRGkykHywP4UoFXorq2unqqOEHpylksdMlCo6FdAY7qIfQ3F
LdmHI2UivmYr7BXsSAWIAK+sfWpFISuIo3FzPqEIq0aaYaMD6r+FklNBL3oD02JYrhHkGPdO5HjJ
DEE8AAlR0mTO9H1CHzO36BYNMKjrklAkKDaenLB7WVK2z9jqC8vxRIazdw0lXYxvctnLHAQgiugV
pj4bfKcKdLSPOQkL9bpUwHymOT3IR5rd7DoQlAWOUaDt1zE2opUML2XL1oxpEcjw1VgvGJlKoTNC
e6BgeV+PAV3fgGFwf+EVQ23Nxq3F8hYp+eC+H+3nwoIX1VmbZvo8Vu2ijmQX/BNQ23DTdfXH/iN4
D2zCst2U9v6LcWUsgcv3r3tWOkb1UbKPaFkkcVZDV7Gdpb06AAFqffozpqJvR/dSNEo522Fkql0+
QkDLDgzLVkHtjqAeipm1iwZhbosDyqL4Y4BtuHgrD7uv4+nSEn7S2C1jIMzhsqP4v0/OJHQ/YnRY
D5W85YUib7nSvDDWnJxFOkWquN1PaKNrEoNo6jb31cGONQqF8OOTK8vRdAwaT9ab+Hb+cnebl1EQ
yy0sS0OYOrMp/0mZGXVH3ezy4rR0yEeIeiOZV/sEyHUbMd2YLIscNwpJOhb0x/N48Jm9ixhddM59
8wv1YXTL7sr1W18+8ReXOPpD/yaH+1K1jRsgOcVSpt0fAHnYUb0Bg2W3p1yUhmIdDCqCF4ImzSbG
3GISE5xicGqV/ZcHUIlxR0CdCSAMTAGZ4xS2ayfhxfR6Hu3rshaTPeYyPPB00muUWo9b2VIfD4DN
5M8qqq/YiZqYxlP4qbYEk3UXfFMCrJNyojgXB8TqS13FGaOXog0IMFnh/0bf0JrSlCeHrSpRmXEq
RFixlSMzSj0L2W8W3nW/zZTKXYJpqDYtta/JGlaArXTnwUWfjKViVjV0x8kmi1222+r5Ps/Elnlv
c+DqI4gpCezk7ABGHx/AYFC4GYcoSABT67guqwlrVHAbqMbIpmYkugY9En/LtPkTT2Wd2XL1bVAQ
H868MO6SCteo7Xx0jIK5LQ35z9wiChVc5ek3e9E6JaD6TSb7jArXzKPsVg2F/fl5Cp03z40NXLXA
DkZos4ePppFO6eH/o7zMgX8sDuSRYNtFB/GzcHyljN0Y3FI1XtBSWa6DeQR1S2vhTTcKTSwsLlrX
QU9EJrLW3pHWqRN8Qd1/csgOHeCVKnFssKdRCLhPhvUbMK4bUALeXSUR2NWTBlUi9P47RO2TINCG
+xgQa8VtbIbFKrl3LZDavBPlxQHTuqOmduIU6alFB8qbH7PRnZ+5Z8w7i5QiUKCJWqVasf8GpCjG
rxciS2s5Ayjmh6Oqv/4RcbODDT8pS6NaZVdNT/6Wa6xkpeaig4xqS3PQYKtLTngx24js8NkDUB42
I5HQEv5T+EpZh6AiVX45Yu2zcEaFy0Ja/MvUggRFTpeRng4WZ5QaWx6lGhqPbl92BgXyLejEeBim
YxVQDX3SpZm2vu0cpHBmBMLQ1J6b0KZzy56g1MVvrn0faf+vg4qG9BX/S9yMuF3IuCiuDIJ8v1nv
4qowe6OzV+yfAU7j6b4nVSzNfuu+//Tie8NkVBW/X7N71OVG2x6rnW7Zg62yhY4j/q6XwNb0whmK
TCUEuzK8+wKePKg6T/I+5vQlxeydM2ilj/Wa76BYjgBe5zkBwFdjGj+9wgePzqGrH+7jbZpa16n0
WTjVqeXQIiBm1jj5Pg25R6U/++3DrXVlhDyMZaLnfolsjI2qXz4PxWfRnA++1jlU2t1cmrfgguhK
LdToEE0Vl+TERQMRYcVihv/d6Lx4QuxnOY/cka0utMFwzTRBsAS/e1DdztelT9rrA4MPRLO+kO/e
ogNA5v+K/YIADQX2dtoxv/BaYOxr6IGx37j3gs7PeCo8TlmjSvPNsezc05/rl2rREwCROK3NDDLo
4TJqZfWOgZ/QL3UqROLjLvXnXLD4e5UDm14QkgxsowdQHMoKINtFpBSwNO8xqL1MBiE8UYWCXYMT
yf0fatflLJyIx1ZoQYPQtSawShL3FBLP15cy3PA9GMXxs6wvp0yoZhHx3XB6a25Ib07dzGw6JEVY
sxU9IcpIFawrv84CpuT58E2ELIC6d/f2o9mTgtIhOzpijSgWJUa8zl837B+W8Yx29dyfdEMfT3uG
bSVv1giNh6e9az9qlRlaTY0R9zOpCNx/hJzd3lk+M26/CL2h1JVXJBESsbMNQJ9fia7JSnUwBtbK
gjh1pzBBxQyHr4jdd70pWKhh9kgwGsGbm0nmcdWuLIcJO4ftObSa33d87rCNT6VKTQ+By9jQZSP6
sgLKAd8oOAzVpII34UwxYyFRfG+Oti5RVAt5xNIFDt0+3PFvGHcBLZx4vx2iNRXzCLze04XyT3Bh
Ew11RXHwgNjq3sqvFViNiMnIsuAl6VARyX42RojgnzUjATc3zsr/NOgbrue0Q+MXKCcM11qdIo2A
Cc4DP4ZZgLK1sfJW0uJRpO/GXyavDwOp2QBYtnyYti8f9Ai3u+3nrB92ooJxWXxUFBz87Ip3rwqg
jZKHBuqTjrzuFuhwF9E1VMvOGCmseOBU2IQtBKsmYR0ozsNpkqVr7q898SsaAeVaADTnUsAMP/Oa
RJAkxV/ToVYO1qNT+FqEr/r7ZwA6m/koi8g1L9bdfcIXCZWE3GEdwZSN47ysrx4ZqrU0/Inj+Q3n
NhaajMU+PZ1sV0KYEqSTzUduSYXqPIrwdwu8YmIxzOEnGcXoGM6I58C7DVBVSeMCzvswQmaj3KBe
cK+++4HXDmXFXqplta+TbPXfGiCnvN84UxjlZw2MCHheZOv7143GdOsWU7omjOjTMhoz+c2//uL6
FYiiNuvXiIOWK69Oqw/YSKhZvdnMap2Sk3BQXrH/p3irBPuaFTFfN9i8I//mcm4AZQlMSo10FKa6
V3oqUUW/zfmEGc9Wnr7XFNOAuj0DvdNdAhLe78HBksQAi6LG/wFM8lKBt6cT240cM6Tw/n6TpEXB
QwIiKoI3D0ejzT3vKyGY2xcVDKXjVQbkmuZaSGhvHrbmAxeh7wX/Zws6mQQeJLw13YZ9p03PPE6R
Y4ppkcnV24aeoF9PkQB4JXVgMUIZHP6yNmEA0GPbWt9mOEB903FkX79euMFj+KoCVS3anbbO75IX
k+GZe2aXYWOR7jjZydlZBi7wve52H/ZHX24/3i6WZ0hUpLX8ZP6DSLOnq27pSOsSIJDAS1lvBj34
GzOm23q4TWjfqlEm1D9pabM82A2E52XDrLWFQvWcHFH0jwcM5yRjdvvSqQypLx7Ao5U86RRPvxmx
q6uAv0bBAA6N2dtYhrIwr4u4qCASe/QRadkDXEolAm8vHQs7rpe37QYaQZwl1P9H+ftWvBzOT/Ub
GnJLxMSMizMggb19u2XJeqOkHfifEmvZ4FhqY0XUvJt2/w228IW57s/Qh/QixNlwer7sc52XbHUy
dU0oj7cMPAtutlwE8fYrH1EXLF97KtSgIQDbgHe5SztiLznOnxIyrLnqBQY7kNFUECXuj0Rvd+Dy
S0DodWHA/kkoL4PkwBgss4eP+EHXuxURZrJn3DWNqYukUAoHrZRKFG5Br4hwILY70eRdelTpZ5d6
ccSmRebWAtwU20hv0lC1CVxY28Yzb8OAA8DLW9/RpByn9DZQKOpaEGtHn5vhn4kErtuV1HhKQ5oK
mwPLRlIaX5e4AkNXxsCV/gk7Y4F9vyxskW99StcbDt1cMmgKyvOFhT58A8L2Kqr9bEmzm2BtHIIU
m5VJoCgXO5oEI3NpPRU2+QHMyVEVgICcdyQGeI0AHX+JQ/cdQGr+Y9ubTfOQqr2ORpDaz7m0/YbM
DvzMSwxEw4WBhwFXORjrjzxpkjvZbUuXVSxOhkzzoM00OaUwoHDl1CyOVDTj1za11CUltUiU8RPO
6sGCfSgN2zCqB+2X4jhoqrfcYc1dDr9GPFbfFpDBY9OJqojsCUQfLPHgCP331Tz29JneH3NFY8J3
2A8WN2FfGPAuSUF9reXydP/io4sFOWOTlo6EXyf4/0xhL9EM0bORsBU61NJMuKccQMj9eL+yNdua
N/nVlNWVH8kvFgCeAxMxrsIrHTw43hhHmx9diTVCJPlgtebcEJ4e9r/2HFgpy4M0R0YdPbby2T9G
bMlmZxY3vRDWtbXRmT3H4lD5fgg4QV5JZVRwUFy0B4JTd6BvemoKi4PrNGobARi03JfArkCyioWO
zg8/+eKnOWKWTuxiomzIJEbab/CWYJZGehzPOjYJJXIg7j6NJ7Wd2qWBwVZo5QaTFPshTzhMx9gl
BlAbb6VvGDUeqmZOJNpIb1qSKw3mrr+EJC84GKmomG91qEe2+cQzlgqBUysvGUI5JN3lDSSwVCG6
gsIYzvn/6l/EoK3F/CGIlptGxlRClJNQtcCUaSCogpEIlrixx3Vbhegc33/4LdCFsiqMFXcK2+W5
qZNcjKdH2gf3s5qkJUBsovNymPZGQbrtq4Qdnen3gsDHE2aO2PKiUiBipdH9DBAtKORv57+Hmgpk
Y2JPfxIsivfQXm6MbPQ1KcsY98I9zBKHJikwmA8twko9hZ23rEljBPHi+d5215uj0Tp/gUHv4FIv
LsNJIJg2a3rSPQSJyrVNN+7wcXBMllh+4gMntlz9X/qFO5ZMUptjpNX77ajPsA2GrhGUh98CSBCx
9OGKIJa3cePqA/HVc5zouS0T9ZtmDBuMfZpzieT5n5XRrSmHoJTIsXRpiUXCT5DGq1F0HYHBiEij
3yGgKUsc7IAJzObxIpIoPkbT8nzUdJnY6pcuw9Ag0fPpNIjaj5i0z8FY7h5+9rE+AvX/h8/ljZcC
6JYhYalyfLOqWzXMVka8c8DjNoPGLzm1sAPwtNIUcqP5lru89Hc2narNNVowz47/050LAOhasjrP
wJLSkXl+47fDkYZ6lJ9DRy0KuzoS8oYmxObhCrPA6Q+lmnofWSOezUhmFzO8a+WqE7NxUtLebFd/
2b2Kq7pHxAzyMjoSHROBEwB1Eu6Y3of3bQ4iibD+3zMxw23kBSuN9PmxvBIlZ6IfsPy7dT2ZPav/
p0ryN1mFJsk249iFwPpLbNvSGXca9/J8XZXYhWEdQQMOiOX4JpdPwEVzpXUpO2eDvLOQxdrTQoqq
DA6c2TbrBcmTKWF7krhMByMrevWys6ANjk0/8ZHWeGLllxFzJOnMgDGk6XzGO22OlPwRpPre4Bvl
/83i1qtz2KAmYwIaJvlZSBq4WoCIcd69UI+GC0kE9WnH/RFWuhgP7zPXdBPd2w+gB5LMGGLhP1v9
hDI65fD7/DVFxOuLrsC7p7IwkhgIkCzVi9o1YLSNYXciOrA9CwQxAXoONsVTai4TtTact1BxXqiS
CPk10Kj6aIFM7mgNB0PID985URefmr73b4DRkF2ErHpaTfzXpT5U0wa8QIAJrUPveAfw7aOioS3/
+4g83BqDlaTRLxRhGQa6GryavTiIaDPMN8z8w4Mtfdz/Tq/yzbYyzGa+GAPejolGMnTg/RMg5gjg
6zBkd+kAJ60mtOHfEw0cZr+VllWdRonUxIMW4hvp2527rOqIvvhZSSJd2VYipy6VrgjXv4uBXAUs
eajXEY5ZvX5cx15XzoOEPnccgDBeadwmSpEakePW23GRKPV3HKlZfelovoR9cQ28nx323eqvVSr+
Xqu0qXCZufckoYiIXw9piQh1mHzXDDxI6iiKHxVA9ZOuzKSFqtWJNhQCmKyIm84vtuIBT8fNwS48
u4XTKEo/Y3TE7qiXfX0bfWDCorX/4mCTMi0CdOiV/S3oQa06/ExhrzQN3RMJYSZ8korSXPMPB18x
KBxW+L251nZrcV3x/cN6G/C6on1Pbn3FVnuT5HlfVM/7hDfCR/AKcwLpfWFz23xvbT4dpWGvSpF0
BiBtwTpKpdfmA+TQsCnGwMIInqmI6sfF9vdZQlcozFRI3NEyaxnDSKiGwtWOPXQ8Pp7dCHoXtl1e
LpObPMz0kduHlWW/0/LwZOHWdif6PtL/mQSFKkQiS7CmpZBtnsYpev1LuZcTtoioOURcmdfvQNDa
VKWHdWqapLAMwLZUYNmFICR1waCBBgO5KyjoJlqzM6uFiHhbo2hFxe5CAHVRPOkuCp7Bl4FI1A6H
E27N591OM4AIlDt7NBwECs+l0Wzx3YsXQ5rXQ0fcR7C8ssJchKcITjBnw3I5FoLS0x3aPiXaxnzY
E1BAyqIS5SkieuI63Iji4DklJs6Gv0T4il5AKIj3ai+cxjTKnGHMv3MLGxfKOOZHnVeUm2NdziTE
6jpZb91CMP7gxijd51ZzC4G/ZPKfy5vs/tXKDU3qjs6YvQtWfjidSSOYxmmIIahkZpwPtRt6h96A
KdJM/F2SDaChebcL29/CDt2XmH7bjWbZPKvmTugeDfAL5ckO2VWwwhhBaOgWEVodfcrwqCqd/WnP
mdOlCkwuBJqaEhfoCr4rnjV5Ij9mbZqJuzMZAnlDEKH/M5KLCja0K7IoHjNvoAh4CMAPOg2Y16vE
Y13iKSCEAMHI+qp8gHp1U0SvNd9YQjJ3t6wgycNKZHRL/lWErIGX2c9StmDr+l5d85Ged1IfIPOh
ev9cTmgXVbCiRilmvOuM6Iv9sxbcR9D/23hSfxFYFH64fZF4f1otPBLUFm5hNBxMbKM50ZckgBWz
dH4733Nxo9Dz3b6eLpt4D0lJ6KtkZ4nviZNcecI7X2yfzkqgaCAdapktdY4oZFcCfTjxclsNy5N8
evCCzhSEhljwU3Q4hWri2whUMK7N498oQdR4970DIm/8GulhlcmY/4bTi575Bb5ElNAJJKVi7gzR
9RMOjIa5Xhy7FZILTF/0SOPDSwBUJjKrmF4gG2eL2A+egiUafL6zJFrbDEiXHF3pVbr/snNkA+yI
whTeEjU8qx2gqlgUk6/t0qw7XhCBkK9FEEKrwlKd3Oof65RnjbpAm25uKeoqB0XUGnZZuE5az3y3
F+jvcMslc8aAfKCYJ4CooQcTSXgjxu2LhXzmKte8M+TrG7Oqrz+GdC1G0OdGRbROxez/M+VtgXTO
k4B9KD3cIdKxjQcsiGdpQM+/4c4Sw9cz3UPpldDwyy65zpW+asJZgaeOYrM9ryx3I5QvY6pGOgsi
+/jaccj4lX4nL+GxcGWCbgnBLXvC7VXdU7TQ6rkEPj94KW/wDAYzefS9omND+CRlLZc82NaCt465
DqRFbTJ8Ol8K2SxHePvUfYS0UUMJhQNsbP4Kpd5KXlN9nCli027amT/5je7Z0VaMzpUtSAYfAJe5
sAJER/HruEP6US4h0qoF/hzRo+YyJ7RH6s2XAlHA8W+Q8n4q1OtUnTV/DSWHtpARuz6315C6PTa3
iVBW2ddPjPU0eRzSzYwaoJL9HMztonquP7Fum1tSVB1TsZr/lRbZm25hOh+slhVh/Q9fYIKxGAx1
7Wsz7pgXMUDI/Q/O/Spbf8NonyhwZrrzR4iwZ7lFR86/69HZiicUV0pS5M9iww8zHXQfxzY9fQAi
qnzPE06TwjPTIfwg0a80Fyz1qWzQ+ZxuL1ngZVHYy98+ZcReoq8pKjueuk7LM01DBUtwMHakKgnM
0W5JrVufBqEWZX9Mk0cS0I5nNblqpHx4XvPSkUp4X/n9Yg5ZtideqPnBjGB9jLmhe9PCRAlr5iiy
GJfJoGilZbn45LA//ZhSa1eAMrnhgsFt/1Pbfv59xrtxe/8A4Yl7LuZSAqkYJOBcymNtp5bjfnHx
B/Laj25cJQQkvLDya/9nl99frpHRnN5dDimjD/rZ2B8m+gC6QdeNNBM97YDYyeDYWU2pmFQbp0e2
coNdFkJ6S6JTvzQsU2NAhWB+OxeYX48yuCAHko2dXjAJX8sc9CSS66sgoD7UGPQKVuZBIsYicu8J
0XxEBlyHxW/XIH7A+0zV2xSeFsbN5QDiCnIckm+R/LpIMvGFwytoJ/tzfO0w1EV3ttausRrZlB8w
Ut0n4gRAbdO5l3DODYwoyFYOh0zgsPYF+JSev7NOVo/W/6cIFdEzGyOKO+9W2Bkxy5M/WUKbKvA2
KfCRDcM6Lp9gumRy0rj14vnZgWuaZwWAYjPxStJl9pfPlqsFkSoW5jvMD4sS/CJRszvR4Kt+k+qE
MSArnN61f4VdyKolD4sf+YnNQG/H3AwwWLlz9bCGMDWNweeWX8W2XXSd4hqbqT0FIDfKmcZ53NHr
3ATaAk2X7nsOf9tyhlsUR41Fjst2gpZEo5/IsMiyuCONh8kG1GBcxrZ6ozYXSJ1fIvkeML7R6HvU
AO8MOS8h+1rA7todyVyijg5NTVptxE0su+2Rd2IPRn81hz5Z5e1jwjAma3OsZXVKhZy1cMVNtZzz
So0xOysLVSvWSKHp4ToybMO36L7aD1HlYSz2BYHH9MK1Z12fC0si8KvELsx90mCoBIjuhzdtmp/3
7nLvmiGEe4iT+8wwFVYrwdj0NEFWKpHiHd2yFEQXchLPc3XlxpWIQGS9f4dKoJL3z43JIID/AKdN
bCIvd9ROYXFmZlte2lUniKFl6WVH9vhd+7LmfBv6ivdsoPvNUSrHAfA0IZsPOjxz5NFzgn0tnF9x
waPmJU1jDtQW2NiQMigSAmilQZhyUpfdvBJqqzjEoJpNK0vNIeRY2zuFJ7zgD1I6AbRs0bInngz0
qLmY0aBTWvQEcS0Fxc4thmu4TZ+rnmSw7kTLIpe5rGN75FPB0EqZ3c8N0/ni2LZ7O5HvZH6JOhkH
75WX+Y78YpIq2ClLVDl23wbnEUipU5JR4dKT6dSfFNSXMrv29r3q+27FsCVd+hkSvkolWaqVBjyZ
xs1Q0tN74Qh0VbHp4ED5ON6kuri8zHx+jrl5bBq8Ine7IF5trrEN39qZU6kpYBh3XF4xP+vgSaAp
RuZKIzQXPnsPW48TNIIYw48mF2FVnuv4bEL4oIj+jQ6IflZGk0HMjBIpQltlDUWvzkaEi69PudAc
hwG+IANIA5V1mTE7Fofzcm6nTMQI0PV9uUIOMF8xMNQXe22pGta/TpK6f1jo8Q5B5Wrjwew6Zksf
e8mYp1zR1y118dHs/nl0TmSMx3t3m3SCkHmAODOWdiZbk0qY0m0em7JXCaUtRKUpZcgREa4GUtlP
aNj1ptxeF+waPI8+fkgWNBuz7aNZPz/FGFboVM62DviOEG+ljBIgJDxKmsPBEhKajV0TCMgKlVh9
zFQIMXTd05EhCdSNwJeFnmmBeoAjXj5CvLkwSn5FfOvJNm5RmZKRMb1Zp3RuV/cW8J8RBCAEBXiG
SO2CI8ZtQx11X9oTmO0Vw78aIS/NaEoxTQrod4eWvEDlW/DoxMO6M5qXEyhTjJOibptQshtML372
PQFKg3cJYNAj8kVNWENOwG9DHEIQoM1Bzqi1A6OXaL0h2gPe34SJKNYTiqMI7tVsH3aM4vNbtBzV
7WV8XX/ZU2ma0/zKVKifb9PTF0Msno+9u9on1hYKnvHOMfzqFbPS14HpSbuqzwU6VXkhr5NJrtDl
UV+SkV204+fTTiNVUDs/fRSDtaFs10yEyaYk1k03FjC05dSbPXuAU6CpCu7XE4SJ6fpMDxSn8dwl
7taSvbEG8vXAlK+aoY8H8Mh5J5y5HWOdc0UhyLDSnueBQuqruVGkWHvyyKO9XXtL2V+8DqY6L1VD
daecUFYnjTA93jd3nvEA3TN1tXz0nWcZuKbU0LKDjyZuHHReOKLlvQfJZOU57Npgh4Lq07c53PJ3
TIsi3yvU2FkZ/F1RSclZMSbpx5ZuiPbEgQkEFY+8AzNMA+T0jTYGmMItDUlS+nxBqD25MOHaRh4v
gw4BWBEZJVptNWgfNBDgJC1Caq9A0fvyAYN9UxPLn/KgmuxxN38SbGOUTj/4pImcP+689IzddD9H
WL/VDbwrIIAxKpuxDkDu+ucldQTdf3afCb+TNDTvQmjxUjIXFVmwSXXBHUOuaWcBomWyF/qP+XO3
Ejz3GcLWeCjC1aNhUmRry+ON4+axcIZfO3X6/CalgyFfStV/fWy39QvzniR7hzmE3nr4ypoG2lwx
sAiidtuKO5Nevk5CTf3nOLhKCR0SLsQmhF1gIrTAj1UdEoIn44AFEW9ldZru1COE87i6RsDU6m4G
6hJCUF1MdlS1+p+b+FwSDjSUARINsfsjLKVuKROrD5rJNsMb1eP7YOTNlLDGQ6DPb9pYYV7PUyQU
C0MRKdJQM8OyNMJ5z4Tgya589MYy1XnumE0lR5KJIfyiARanLSI0ZRgJkMVwD2CzFqBpTAe3FkL+
f8AkCdfKXiTq8kEiUcxoOv39+YB8ltVX+9WJrOozXG7MWZS8x6U87x1/znbb+rw9beou+S/13yPU
1KMyPSWBodYlSrcIoU6Cld16I5HArBivMtRcnEfnvTGModUU1jn7Zd+9/iJ6bs4IxvDP4QDgucnZ
9Sp4l4/3VhH3O8/IRciz/DOOb5I+W0J5GfYD99yY9t7rHLB2zoePthoJCcX72PBAvsMDN9yv3HoU
Gk5wyyAlvnyW4SJ/C2BudzkETPMHcFqvgqAGu4pqD/Uktyja9OidPY2e+ttIc2TxbUksThYIu/Ek
H1X4rwzKfQXUKWklM5A33gaMWtDnxgL48QKyJ0ZIzxc6OM/lN2NqShRDz757pamqGaQ8z1j+kCcY
II72Hqml8ySCIZK9LQTZvmsz3jz2aSNTIAxC8DLWiOww52N44dI8UvLh5ki3LYPiAJbOgYOgjMsP
fXlzgtmiG5e307HCyUWoq6DJzfEoknuLLeZ8DQ9B7GnoyajRLCSi9vvJ2ux3atLG7Ri88NknjS+k
04E451xkxielsh8tBjtee0KTXYpC7lGMxxJTPZdAsudc4m0E5jFuAzJTZ/c2k9z663INZKrFoTCF
jaBYRci87f7QgnRWDTX/DIm0SFWG21HptUycP4axjtnBCZk2SJbZDjUn2TdpLqNr8QkBDt4R6tdM
XxHWbrSkIidrAqcYPh+nI5pT5DJG85oJvfuvYvjELHZQQA1c06eGUgl3PK5EcXSaCCF9LzQLhjGI
efk/GXunZ7feiNxW3gJDzjSBZ0RIOQbHXmnua5KHM57ywQR6jlbsvAmVrmFm73y/ncpeeXfQVB4K
r1ckj9ufeSb3dAQgvvGsQh6ThWafhn3zhF8Qv8yexWouvWku/37lM5S/hSHWxk4Q1CGUHWqWQnz7
Nmd2kmHxL8LWFrMavwRavLz/pR9N3xyuDgvUSF6c7MeeYBsPPqOHctKCq/9bcWavgYrZBEVhGoQd
VyVZcw8JSJZFc7+UnPXdb+rKHuNllS4uNdD5/MV3wShoTTNiCQDlVAMp0fYiFd6aNKMh7Xl55zgj
FwHM/xZs3cMYbieZKzhPXLEJ1M03mdZ8Q7m+w+BUmZQEdm3vXbaXnlLpFleT/jlbeRvR3dNFeP07
x2caMM0AYPnNu/la+gniKjgpTa+LRwk2y8ekjhe4R73DRg+Hr1tKpv3p1r5mK3Rwpg8wVaNxtjZ2
mkpBoUhQ7z9h4CMdDY2XqlM4seXUS/iBmlrNr715y0AEtB1pcyq8sFCq/shcDP+k273rnXNMttM7
iLOTbjgGuNSb4qjizYj/kEtQ8cXpfEs7DFRlT9tg+/91Dj/kLKzX3+Fk0qqRP61naw0kcORDxuK7
ovM7Dd4qEJCh/KhAw0vXVmSN2iW7m0WvZyf1HL9VOVf3pZwqVTzeKcNbkHY2wN9MUs6Y10jAocSn
1Vf8nOaaHz5Y8KWPeAE+voPnwDPUqg0sTnNkyXAkYRbzzAgPMhYbs6uGZtdV7PmK47rNu3XcY4qj
QgmM6y8XZGVXWiRVORvzjHLN+deWTOUCzem5UzBSeyP06jW6sVYX7oF14/ICvh3Mwjwh1UHJ0XQF
2oroGfsAveZjskLf03dckOjKu5dQOgq6tQGuc16OjFgiOrp8MwulFRU4aIrXeWt/cjIiWNJ3wOG6
BakwcBXxfxBcszfijXy/pDDebAm8lNEAT5XSelJV9Np6E854s4qxFFsyToRuupGplF/0gyhei4Np
mlxrUpckfVFbYmWz+2wbh+ulTArvOZLv8s7M5/gxlweadsrZmn35yakFc8/vC/cQl6wU43IO+xZ6
vqvYZvg7wn8tQjv4s06BRa09iIFOy9L9uNNQC92UVeS/4Ea21YjbHmGg5tc9R2POWWV305CmWR6l
pC4lkBJWLlWnZBE52Ef18wkds5/VnduI3Gq4hYIpNNTlYFEDF0lWBtfQotKfzTqrGKCVxCkP1A9A
azT70WSPyQw417Jq2UWgjsTCAk49tMQU6xXxufYGMAidCuqx5liKy0QaDiy/zt/095Z3bW5g7w+Y
MLMrISuas+HU3F1APMtV8s5e5DPo5fgRFpkZbh8Hp/CrHos+nMt/gLRNRyMGL/MxyhFVmRKeSz2c
DjhkXmaD3crDNCYFEwLqzjfuwKqI47ZT2Z+FypLszIqTMgvbT1ZXj3/WybLjl9dhWjr8raP/vKmY
1ZkVs9tuUZxUN7WN3qZPkGIiUtVLk8P4Ax75zpvzvGPb8ODIFtpJTJ19QaxbL9wU9HIjQQiKIYYv
ZoSTzY0I8tdd50NwevOFNFwBFvntIsSPtsNR8PaQUz0LPXf25p7YL+4YkC1qqQD/hHLQ7mzsVe1O
tfbZq2qMQKMnc6oSYR/pP2hViOz9o2TCxzfGxpwZLgaFpzTcH1BQmwEhSVAE+E8hxkwbyvr6ow8I
i89SLSE3oNCqQ2kgUClKDZvd/fIQQ9NgPmlB2Zq0xZt6Gd7xpctTOCUqxiv/it27XIN2P/qnaNoz
jQ0bc6quh8yimIBjeVcBQ2nzOixl/UJDACn37NfxbbzyMD4pyhDC++AzIzhRQ+rjvo24/qqiyqA/
Xbra5EatNDT1BAKR/grvpIkUBuOFIoVlawfjO/F/nIVGLYrPY7YWr5nKEO3BmeYr2UPoU8cPpFgV
1bTQxsr8q5589uWabXcIDcD2l/jxxMUJ526q9LxInM1cUMD1FLIymWDIoKo/93R3UQqc2hacz5DD
NobUWmj4TME+Ov3g6dZObZnCu1RckyqlFasdTkpvhORLNhzhJYqvOOSTvi71YoK7QL3obFMxF0ay
aqFOfxg2PUQ7YrxJinXHA+cBxV4LQ8v4Zjo60NL98ZvfyW5TeTHYYV+13sV638trxSX1S9g2w50K
YqBzFPdaM3tmAjuxkuvkxj4PZqMbZwsT74+BIKe7H1yMmvtfOBIkMkHLqpif8CuklfplKJAeipqC
CsiNIA8esEQmmzAdKxasHTK2Ja34nEgpaVuEY0Q6vKg6N/G7LlM+ZxC/bX/votexyC9h32CJKWIH
UphhIsL80tjvuISshNvmtu+SXS9N5v9eJrr3ATkMHk5zRQ+pwjjmVp4m2efXXwqAUeV4kPi5OgVe
y4N8GCcijJP1chGcuqZ2EkHXK6p/2oenoWP+QRuZi+RwVFFOqzDrL7G/NxXwuqT0fsF4PfhI/gkp
jdfk2kK3oHdkcilRoYL1xltuTMgf4jjxgvscSlIM1BeoXHC2URPZtFzMRWZiygRqQWB840z6nk7p
wRQsBkpHWHpORih6NVkUhVb8rNYw3wLqRiP5TN6GXj9tevF2W931N9grsSeh4eUVI0Rylqk74llr
RDQWOR+B+6vNuQ+i57tWLEIa0wro1PWJPS5soV8irPkCbByEUNM+bdfQDDAFlpHr1QLRAWZcoPBh
DL11hVB8DQZfbtXT48XEi/ToGlsYqQtLJym6HqCEO6oXTCMsvdeKKtawdMeuDfei+UIJJqovWjtu
9p6XH5gC/w86hwlhLFF23VReBqaPxv44j5q1gbSGV0OD2rNxRDBYuK6H0XAwzcrol83QZ6WSWA51
LWolSEunCtDGkEx8B1wiM/3jnwz/3GopiKSLq8wosUkcv+RrL1JhDJER5938BY753ZovNtBWlygw
ALwGKbOrRZ9Yv4VzBKZnOV/lHKzt/CJaqNgxIkTtZozoYuuAv+fVlsKO3Fkn8tvWAdIK26EILZdq
JXiYFNHFYcdfx0jlZkSskvf0RxNWhFaH6X89ew2o/kriu0yD5Il0VLRAyBbItOVKU7AVOlUfJCWn
cJOv45S/eXOQS68I5JVbqpiHR4P9Y5vYlBf55qL9NQlYjZ8vZmGK7BjcCpcF6VlPSwEfGC480Y0l
jp2L55edOk8bELvzjoB3+ySManH81xOjQCz6Yl9n28DU4RiaenxG3X36Su0YJ8S3/ZtrwDdyVSxq
phnHB3a4lRmZfmUI9kJ1iVsayLnOIsqlKjL7wy+WekDAxWPO8UeCNydhNHifyMawOyI7NuCAh8Jo
DMKTIVvPcxBTuecUx7m6R91apkWiIeFpxD5KJTp/6scvHbBsysaPZjLjGm7L4akMZW/LhF486hpJ
kMg9rtXrVe+9GS81SuDJjpcaCVBULPGe362AttAuDioeQ6LK6difj33j2055R01Cr/MPlBM694rn
N9AIHBFbOJs7OGDvOjEfyJZl/wFETBAmKfBGgLGFxJ+3v+5k7k3j59qd6ryO+k6qp1vPIMXMnoAu
6QWDgcPKG79dkRt0rOi6qUn5OfAuZPix89+t63R9VSsE7tl/IBYhldELrFIypvK2C6ZOpHdNQsNY
9MLQNFsPdKVPK6qOTOtyrTJtz45rsJlueUvIrUdFvnnYoHfzrFRzLY6t8CQ2TDzjj2lKEr/wOApY
mplnLIeg+fMzadeUyBf1pGUtzbExSzwN8U9ql+Vnjd0g69aCOleAIO0UsD660AQ68QJHYQ2ay0VP
uuObuMqNeiMALAr71m8JV/9K87jWuKXxAb2azZhqhQC9PNdqU+f51Iuc0NvbIR+IwpYqR/xVuGq8
DoUdhmS+kSM0MKkmi5YUU5cMxErXHY65veVkVAX9OKwqfnXMi509Z9lbfHgqKajtWLdWu1NGJT9R
H+Hgj7ZubPkMiENMlKkS/FOH7JfpCqJgKBBTOZNxdTngmBsFord3sZWkJnT2MPQrLepFyEKYvtKz
2Q/GagwCzLllQXBYj8LlTcE1vjuEgUfOlDViT9DiHhuiGLhE9P77f7bKBB7k2VTo9CG/kgDxubYS
D8tlG4OT+6AebIowN05jNXXUbUzl2JfNIM+wqqMC12Su0oHTsR9YQ6+Wb3laPaB5dVF4zwj1pXnI
UlmdSLF3POSAqh70y2OxeAvRz+wGP26Eyz+NKQePxlm+gSOJTIN3vKIme9ZcBvM7jB3I4MNrfRq+
SgIImgQPoHAWH4V0sO0jAKElQSkE1K5zrt7LUZD4W/XxW8arj6WNcOEpoJRC7OUfQY2Wxz3CFW9l
ooOA4PTKRgIFy7BDu7Hd4Dba6+2wdvO3qw3IJx0CiaH2S9NhJhdt/DWtJ/aXPOzA6RfDpGHi87ED
GztlpVVkCU5r0nEE6kIF0SQXqlbV5K1fP1Mzep2VqsmK5/6jIJSaYB3cRPB9cOoEz06hGz66P1PJ
N8F4fXVaBmv+VhUzTN/32/v5BrlNYqf7BOYZX5KjQSUIpYgedubbScTHDUxvqXx7wipcsLPzo5z0
zw6g6t8W+PGGNitYdp0BgL/h7GAHmcSTfFc3WOwk9VdLdSgQAj6IgJtmevOUw4bQhIsBD70D2KZV
hPVb06KKyHP7mGmbrHgS2wnWZCjNyFCgRciwfXalP6t7GoSdBTy8qBDmmAh2D1fVkeDp7T79Qv5T
NsUJ1SmLefSzXcQjcVoVfvUAzMhNfkRxC5iHJ71q3ApXs+4YL8w/S9LBRNfbL6t1i4pX2GxsZ5X5
XVeUhFOA5RLZPG/iQQynTy/UdL3BDIamQIfSvDhOGL1j3Ft7rkOeh+F6GNSK9Mk5wBQr/WlRT68L
GxVQH1Tckj8725msOncF+iZbEC/0IFkIFxvB8emUMTCpP7ePGMYO7XAOxRq+mKCo1djWolACQdj8
9358k+mlNHIDfDTDpbQfk8qXkBtlfYPSofcQcnGDQroZ2xF2VbG+abFHfbjkIlV5fq/Y88r96fUM
DX2DjgXHyyR9L1D4h0SvdfWarYk29J7ZxOhono549A4RNoSwvb1cbWQez7CPIvag4FmodsxequML
m8H2Gx5hlybrBFL4vLOuFPZgh87OW+bUU5J9z+tMyjB2OhDeTmG8ibAEj0s8JHBygo08WGZN9ggE
Eu0YzFPUXgNszqR9V7gifvv1MF7eHokoHkrDviBNs6nCwsYMsASSuQQAoYusSFA5Aw6S2+4viz3G
M5xZjT2HQn1XPIsd9oGbkPwVTqRrmQ5aFEHQ/fc6HVBj83aiZXOF2lQ5d1/AWsOYBaF4GcA47P7h
iy8FykxhdI9dQ58rKrsS8xSNCHFAbzlOutgPBmZhQotCVesjx1i2PERFpVgg8p/dqrlnHCiTcaRn
IC/mS+p2JU9Xp+B5cLorgXS/DDqXv/JCGQzTVZtYeMDD32QdW0txSYoD+ODhto3Ge8ozqUFk7L8M
pUlRLsWXIOKq1t/fzfkl6Kq/KRVUtH+Cw9l69LljD5OHbzBoO1nDMPQyEfwbP9YpJ4jdtTXT20mj
M85S1bTy7bk+3YZ9NhcfZKjsQHwbBwA9gjq56/5hYi6l+Vymob0YoorAcO0djUzEFk13SyKk2twP
n3Ls6LPH39C8yiLxV1uzDB6015PyMKwlFcEDvCV0AQRwYrzitpmDKNNTEBNuOGERvXT7viods826
4InWBxIlJZWDwE0JyZsvPxfx3Dn7tMIOJJZ1tQVQNFCjT+YkDSphqo3Xl0dCz5eyxKp3IZexPcVs
C2TTuMwGHNqnE8jO2HCDWvdH0oHW8124Wbw6ggiWA7QP7hrI0yeviAmneeMqnJjOo4WMjdq5vLqh
uYO5aaVuYLbImWTrCbOO74/JtBUB68uiaf7cGkHcIEZCPsfBk9oOI5djx5GyHM7sziH9iNL0UjcU
v/I+/jWMeNZ9SmwP5OYtjVMHBBD2scghk8/S/J9wjsCkOZuFuKm8AA95AfQdFHd3CpFuE+7J6Yg5
k52wev/iCutnx+Rdlw7ib9tvkheIiufjfq0NRUNn+/GlBCjTvl3bzAnxG/1eCK38ztuzjRWRxbw4
GT27oqw8sJ+o6UjEbQvUqw8GHl0CadiNFYkxWF9YraYB6RYggdo/gSznDM8b3kqhKacrZps9GbHm
XPjPH0P35xV4reRt3uoh7XS4ljyH1b5YJOBUd6XHmR9InNhDiJMi6g1BhHlEA0CDL9zwzO4VLMmg
4AbcyeRW8VBU2kcq3/C38V6gf9yHofAzYWOrWVmcFVitT7aTHDlLEnVBq1Qojrt/fqawAWmlSH0o
fbeWu/HKkDkw/EzdszXMA/DwBk5F5oYO4+v2Hpp+tJ5Pwcw/Ol4QFHdX9KG1dnXF2Ha5qU8x1dXt
nsLcq3o9JJy0QXEMmucRiJ93Vy5/vGqvHONmbSrPwBq4YSrQXv946rZBN9DRhLafLXEGmPe6O9ta
RglMdbPI0EoHnpVY65Ng5itfzpPV4IxH3d8VSin2IJg4pPbkOMybKin1EmYlDpWf5NPUm0+DkfL0
OnzUhqGY27AIjrkSXTY6lFXVmxxTg3NiSq9Z64rQGMiu0G/I0KwDr/UuSwqsJGyKeEW+jhwCht0C
ck1MMgF1oxjwovEmfDCB8eFwYs0SwhGHT0+BC/7rdpmjNVJC/3A2YV5Y+X9M7Ik+twyCUfFkO8iu
cSfbIVHQ7H/er5LOwcme8CxBp0P1lQJWghMafjtROc2/UvmFHKruGvnbEMze5TNo32ShTxcTwcf1
tkr7AnTl5hiT4k9PxGBe7dOWHXnq6x1GU5sts2lP+t53hujKs5OSvCscXZhpIdBZBEEuxJwWp2IO
JyhCcB2xjYJjrNQpG5aecw90w9WTibExhi1OypOZAtiqo+Z4HggOKVEamL720JO9YNHgSQu8fx7T
4bTWFLCjpffAfJWRN82EJN6+nfF7r508n1oHWHq1ezznymY7r1wRoBMZrLn3CX6fZbXe5bTNkWSF
SJsH8BxacQoseuc0TuK9q/xjKDmzvP6AtKJNAbFViyZqkSSy7xFO/S2UPif1tJyS+VYYcpXvKDfm
fmJfMNBe4ij3NVkMGmxe9ZQQ1JyU8mtjeeqNgLREHAr89HIiYCySxi1PMctxYDbGQK2M4NIXLe+F
Dr36J4FUXCHnniif5ttRca4g6YRYjLDMlxrk6cq4igDgKSNsHRfEEpsJ8+J9I0iMc/zy78ZvIGKS
B4LLtcaYGrXupJpC8kKL3SoalFhrKhKOoKXhl9qOj0Zt1gDh3Ebd3l4nF6KYBKzYF616oVpkn3lU
cwI3+cda6BG+OqhBQXlwg1D8WN2WsxglXEI5FV6lPPMgja2oWD6PljtphPofiaVowyPVK/wraxP5
xNPRbs1luNyBnVq08hPJ56r0l32vC2WrxRsg5/6LfchWaoVgkIoxPKWUD2f1IJXOj8DnyCm5MI/w
n8+DcrsBLrz4rcwQWkoYcAF9PLKNJ4eyTEFSor1xfh5h7Chja4zjjflQ7cXRoQftt4VUTTDU+j2x
Gd3Ran82MJnNHSlR7FuRwHEg0FtZqVdufv48uyvTTb+UhRKXNNxUAqFhtMfeQyOHevhTPTM9O2O8
pcl7iuT+pfpR0ohQN5CsPJZGMpr03RG40VtHiq2JxaoSFdPIP5CH2zYKV/ZkxkGTg6w67LyFLGAc
M8gGrVvxV2tZjXWYIYyrpB15U1oDRF7nFTi2dyhX7kOvnukxt4crOOlr4mmGJK0iyX//QdS5xwUN
IOSH3i8sIf8a5KEmOFcyckuPpf4BJv1WXciiZv0WJ43d1oanf4m9jm8WEm8t25XC9tH/r4QQrwbz
Xy/r+tmdXkS3sc4/WmswCtDQbjg56c1jILLlFG88cXEYj5OEPJtkUaLoJkYO+nRzKNVs94hRk1xY
5Im45hX/xOMs+AjKOIHTF9Zi4GblDKlXmwx4rWHmpNpNU13ctm184XS4243NCyUieNuHkwI/DMVh
kwX6d+v9/eX2M27w64qh5MER6a7iQDvnfdzmFbNjGjc+hUJHZY51Ud+1vo+vlqhCAvsTUxidkaSh
ZHA45Z2rM8RU1P21Uqts902ukF0xPeDPqnPzaBQEc4FejySpO7OJsu1kJnEDSZsnE69tGl4CdYq4
qX138ssIzJBjWPG7Ck/rxn2fhjncA9o1WOs3iqhNIiDDBZbpYqE8+YcfU9jANXg0UjH3YragVZ8A
DLso6rZRHBqDsqYGot4A/gNjcGk8oR8gyb80/KA/XAF3ALkIifhk1Y65SR03BG+T/7SvNhMhR9sl
ORPCCVHYJYdCnLOY3r/KLqpvrFoS1OToxLCo+zYEeJcSpGBWjL4RgK7mbrwvEaB3B6CTopp4upOw
mdLlPdCCmCgf0hfqeACkagZYCvdFXF9kc+YK4Z5+E3r8xGkGLkKpkANCJkFUl99NH9pcXH3brlrz
d2nwwo52mdtVuZ9iT8B5cfjq0ka4I5krUTRT4Cm7ECPUmjCxS6iChkolbqNZ5V1YZ+RVjeWnFNTe
7aqtC5unNJxCwKGYKot9Q/5CKylaeBgw9lqeTAaUxyZh2X+DGrmDekpfen6MiCfhJfk5V7clTxem
p702uinKwTNajhDWw8Q+Iae1iB23GtO/Lg2V6nbxXZe+NlIInDIx5GwvhX/a51gWempiaDfTq7kE
4VehB2KkQjhPsNY66e1N4JI6GHq0KTpavlt6uwWlWWFdnVg034lLilYL1BaT7Sf14gLf2U13NIoS
2Q8MQVnl8GQvx0MSHdMLCgruuzk6Zkl/w0hJzBVFX4A9bfWhA8OtJqQoAFHG1WjGRBGk+x24MtqZ
Hdbs5YWBJactr9OeT+u7exXOZZD/pdPWYRCKJ7TWPUbRCARfDzjWSogKHQHXXSwW5S0oSwe9hI++
SLkYtTLnkDLZrN3TPGeHew8Vc6zfMq4YyW9H5J5tCqRhQogKTvY5XVPxm0ApGhsU2TX7+KPSqhDY
8jS6AousxiqXPDxz/xgRKU+aIY9fiulkNz87smGzywNpwVE8RS+CMGZ6fiPhEosjKLnheSghrXWQ
FWTU2tvw34rE5CsCbjfY2eq+SeZa+cpCqQos5FZVMnuQrlq7GGuRvXvZn0lM7xdBYwFUeIsS2N4a
61yHmWISvw/tUgmLiBpdtgLDdkXQjFu+qtHWIDGOg7GCWkMN/vtMqPqDBjcHPWWeG2JhhVVVeBeo
EIrZqbzXI9my0o1RH/94z+8y553MVVyBfCxEQrb9Mdm8jeJhK3de9YXg+o3rlrrI88yh9S5mvTDG
rBORGZfLz36k+zyI8s6MKWV+9IUb5iXDcQGLssG4rTzjqMFsffPdAEBQ0WFJsWPIVZIzVRLpocjY
FGQ7cLDrrEP9kpWrPD4r+U1Jq0nfmxGsmkGwC1YgfH3izYy3t4xUE0GALms3lFSngxeblQ0LP/Rm
WqencdrW4W8o04r+1/GO+rs/MHjeqmBvOKnv8+K94lnQ05tXas3FG8WaEFLnAUo2wYrN+MoF5YEI
NhZjU62dhsuG54SbtghsPASVshZ26NmgTIIcbdPY+pCeC69SnuR1iGhT4+c8eaWDvgFkf9iXjrza
zEONrYq5696mU12Ra8FmCo2DTSvMUqkN9l1+hXGg/G984fV5nsaAxFp88zQ0IkIdcNUPXIuAKAzS
tCmouZjhZAAQL8fidX7OuTCaOAqXCu140efkzwKhuJ/3Et0eCgUk7HSiHgJg+aGWfMuD9ThPjtJG
TP1wo3OcBIQkUB78Ggy7E+2LbBamVhyjhV53OOmf538g3cEBIe5T+vtvpJT4M9wS4sL2+exR61UU
/KMDP3jHpbRkAB4MY1E35VbX+WobfkRecFwvbMfh663uaViira87rtl07WQMpuCQfqhIg52P7U3t
cN6WECw8E/RKpDjujlLCD7Af/HMQFxUQiOUP7ykKxz6OTLIJ6pXkqijszyuNtVI80YKxM54uMjQX
4WqRZv9sONOarB1OjSOKgz8qrNH7rP/4PhH3B5PYPX3kog9KliYSF21TNXu6c0+rugtEHpJYQk/Z
f1rPsyEcvmCp0l8VS2r/U02ZIkZ6pd4VvfsaLyLLkuJmq90TZ50tAcI9vTlnFwq3ZSUITIpxPau9
EEWiqwcgJ6trLOZGUphD3a7L2O3214s5KPyB6iAMisNcXZRqleGFhodkUotJSSB83/AhijVt7TuZ
be2T5S04jQmx2nLNSLUskRdxCBuoImjdLp6fuxDUQErMf4UXRr2bFHsGCoNj6YVC38kk0Qg5xVh4
NWxKJQORLSv1AqaTctnryFkzu4Bqe0MvCGQLKMWc/2/E/neZfsPDMwCAv6U8IXY7vMjpOl/yyYLl
bbDGZPNbKxwKEjDJa8b59VyndXVyG5AQfiA5mWPo6RBH86S24GlNRhntH4Q3JfVY9G9EXOAewSLo
9u/RgnHD+vNXinsx2DNHzo/c7YXEnEl1nu9mqKrpj6pcCOxwSLkG8mx8n8dTnfsdsnREP4ScMIRR
IhKAh37kuCl2CvXiiGdJKDAobfF0u2BDIEeuLjWOX80b8Bz0VrUDXV9HoQbApVaYzV2vrAQyZvB8
Fa/LDhXYDLrJlWgO1svsoA7JWM5XpR1okQNHI+5B8NregMX44HSFXNn5KFkiMV1veD2Lt1G7H06q
3pbXY8i9cd259ZTlbOjK83mJREhAlwrPS/e59a6WrQ9hYc+bzm9Gbf4B+9dMKZM5MhLvbePOwT8q
so/UPEJlVxwOYGjYdKk0m87SAn+qYLVPdUYfeIH1M4dmAHnGL/tgrsqjZ4VJjdSbOBeJo3nffxaz
v4Dl4OpT6ZA3xEnC7FkHNctPmamxVTOP/fvOnDecKHuVWBO54XNWaYV2nZmVGEmAXAobK4Ru/T5V
xEC9kCHMXeBNCC59MaeecJgMv7iyjL0rsVYyYL1mvITPH+zO+EjZMy4yYY2ZFbpV1GctC/QWiOj2
GcMvLNjFn4WNLapwTKTEIlZyg0nmsMeAW8oOtPAR89qTags82xGjv3T74Om9OFVrs6wNDPLwGkQw
UYQQhWmflgHIkbqW5lom+hQvAYlrn/bkH0owRc9O+WBnrDjuiKpRby0QegpjsLx9991u+Zn+QL0B
0iwv5p69vutQzkogFwwe00UzxFHfr3DBXbUhFYuiEhp+Db7iqjllzxPiF4v6V7vMpmNjjuywf6cq
n14GpE8EOxNazjDfgKlZx0m9GKhQ7pLRA7Cqfk4U1sgV0MUkEl1yEDesQNTGfTQ+7QpY7TznQW/B
zmED4JnC+Y3bNGFFCE1NzDGP6G0pyMuCAi8otNp0KPB6W+JN+psRQZDBp7HbYx/26VRG8j95h7ZT
EdqN6hdOYwu4mC8WawxZrmlFNKzQHlG7ypsf43QUoRvjWPLowaRwnDMsEN4otw2bqEUTePiPJ3GU
ASlaSKzyNNReRwzeEiAxY2+MRIlAjLMsY9U5eeNYVCh5IMzjpal9DmICT/AlLFBE3yWRorFiBMS8
O9TcfzJRMXDYTJBa7baWeV4wm9RCXwlGRMqbmQXBKawrYh38g9jKvy0FINFnC0OcvjjqyQzP4mty
PAi+G9c8UIuG6x8trx3hLYJ4dGDIv9obucvz1NvvRla8wPOBG9aGEOVc7e2IAH1Jpoukb+2Mwy9Q
hVyToggxyOdy1J2wU5R5bBR7EFog8fDxAOM/lVwp4QqVbc+w7mosrIxY4Z0he+0553J5slL6XJhH
HRT6ZpTSt7+4QjQF1fM8GpzFrgKBpMzL6/ujs1QiFszuqcLeoFt9A8smvULuyT03kxdYkJqjdxaq
DsLHwvcK35f9S0VjPclO0EIcCvQ7U9CMNP//IXeVS8EPHuGu6+WlS/VGcxg9jdBhBtTlbGY8+Hzq
fkHwgJS1w3xotLw6jq8NhEN1TRdL1dL5kWOH22nYdcXspbMLpXBU3IDaE1YpMF4g4BsvOu9CD65T
KNJd/wxGMb/NtG1YXYRzUQNFbtrgdhM4+Pk9F0MqmuUVycE/ewI3yLN+5Jmm7myhH7gFpfuKs3Am
2rvpdMJ7VIqlea7rgLK8uh4r6o3Kb8VB2R6qosLskvZTsj/UGsufPC7eZE7B95lkVlFWH0NCeRF/
9yJmMbbIjvM5I6NkUffAdHXgBWOMpYGK4AD1zl7N0amvpN16QU0FACNNMSSAHHl9aUeq24JQAUdv
6vP7Jn7/oawLWP+Wzm1nVLzizciLa++ghvQC8Jo6fWLf9HnfO2HSFkzRgXVpSkMUZcFE2LQKu/Ej
qLJmylNoY5gYjcE2+eC45iO1TKr4qGioR6QauyDfDFgYjhMQKdMdvWy6oqg/4H7QMNs1CYLGCWT0
tSYzFoQ2J4KNrN4BljP23vCYS7RTqPdDcEwZLRsGjNPh4vjh7YGXTHaJC8sxclYiGh1C7lq+xkq+
caikajTXJPlvOsMwbB5WRYotoujAnHn0+LXMsE6sTDnifC0YwpqhLJP8n4dXrycVdrbuJqWeeV+J
DI+wkyl5EjEaLy6lBK9a8QC2t/1bYAIVIgLk/8O52mISHOA7O7xxBYRh3XuSvIrOCW5moPLzGJ2X
1osJkz7jx0RjgLa4mEBonGWdFfTGI7KtMX8E/1R7kd0UDEbgYtMVsYFhogscVaaKMQRj9z8mXJhJ
Y19aHk/2pvbrjZee34iC77DeCKyKi6TIhcaL5mNvU7o8Xfe1ah4V4p1XMZq2mgLuzGd/gb2kguf4
4oYlaJWgE4zVQE7Vz5CJTnT1z+o2F6+M7F311//cyCHn9IMyUk8bsvaWuwyZoTvBUx8ciqY150tK
zANzjpPc4zkABppXe/x2J3b0rnvVYt9t1Db7Z9octjNYt9F2Qb2ylqd6WDpGfOdIvEP2u2WK0ZaD
3lk0tiQAG8xd8sNDPEfw0BXlQ3WmBe7/XnXYlU8BxNMaQ3QiELrAmSv2SPwwLno0WcNyMjl4p82l
GpODrSFRLTXc/MEKjpamiVzJfioIY1pBS8QFTvOYATOEpqr7XryzInezghcM+zoMLmaN1GqQbCQ7
ZZv7YzRV4i0UcnmW9WKUmcZ5CRrwnj5DuT0/o/fyJcPI7DhAu9D6Tz2LeDHDk62G4CvW4oMDXYqj
7ffFtv/XjeltIFo7k3x/fF49OL/4AbXp44xEoE3DLftkPGEQ9g3kUSrTGzG9n4JL3fr7biIHb3zM
TAdn32k3lxCxd/jnKeR2WdwkeDulqN6Xf6IqFMbzGmq96EwXAqc1eCm+149ruHc1eMdLuA5Q34+v
NbcRvi4bmwz+IylsItbwqCkDwQYo6pjdQErlrNu5d1HL1g9GdeQ40WMoJPKKJQgO7tWqCJyzDFy9
MIpzl2DoVKSnc54Jxp+O5hgacuKn9JXZIURPpFesb1G2RFU6NWZO4QEJly/s5bt2JYeq1LfEh1OA
topUO2eNKH2eh6kjxhGUBr1g49f54XwT+V1GJL+t95ZxPxcJUyUDfDQpYnw2naG9TFvaDMgbuGcd
1SNTIkuHt0ogyR5pFCjuGi3oN0KXHl4F9gngNqt4uC+JcotpmMZ7Vf4EN23aVsgtFofvLjPLKhjJ
isg53s3ebm/nbmNZV57Jl2Wty7byN6MjbHFsSgxqkJfO1znjEIjQNf6+NOGIyFSMUZImHBQ9sdrR
wPq6G/cmb1KsCb1osyAabRzHZ3glHu4AO6wKW/4MCoIp1x1yrf+OPHxEyG4tL+Q/LhkF5ovQ+ne/
J3Gt6oXNLVdhVgxmOVSrqjqYk1p7j5Ws82vcCla3Ik1Ub0BhjIM94jNeK1TpoJFQEsgDJ8QMI1gs
mKBHRutVjGHr/X7slm1GKF/1TJIpj/i10sYE9DxG4LqTFd4ANSL/N3I4joPrVn25z6Wo+sea8gnG
jKHbJdKU/AgEMEhD7maEKM+MdKTNP2Hpu/zf8kNayZBKDoGyVAX9ijNI7ohmBg0+118UubAdUA7d
++p9DrdQzYfWSRWH4tXfZnnRgo1Gp+jamx8wRi1vmmP0rBA+0W1yOGfiM24qGERamliPm918R2Q6
A3r9MgYi3bXDBNRPrVk5EKtjDUkgqoyp7q3LI+JVzioI8yfA5Xfk2OuJdwDcRHYYprstyNiR8kgd
L5xJWvyQBXZdluQVSlqjVrYGN8PR8x/F52EbIRe3o3V1ECksE5r1uQUvbvh5LrxfJ3cJnPPFqGrn
b2XxqNVQsNfEjYovoO5pIpzxr03bQzEHAt5ktnwKCG18u6MiyWJyL1u3T9xzWvzNnmCT7CYYAGlf
296MWWVG/vo7uzQm5ERko9IBcY6cmXucf9fAyiekr3awu18Fd4dAeb/P6RNa9x9Jg/yxisp5MK91
r25/5j+QjB0k+UrBppKScTD6fXsLTO5da/qCyifd5h47hUT13fM5FE2YOeiuNWfQ+bPqvrT9p10m
RHOgXSso865sDgNzW8UHvvtrtnyvkUaRuAHiFvIUtLuymfsHAMFpm/BdpiAKwaP8syFphnMS0nj4
fWAK7xuPn+lNUECvLww/ayo6KM+kj4K4V+2oh7eiQw7HRkkYFUS5RDArTXuxcKkqrmRyrtrWZGQ/
47Rn4yX4zcVJTlJ4oLiafdQCPOaexqecy3SHBUfBotEuCRix6NaCZc7oJ670qoYH64TcaD2Ribpj
MHFHOdnuCkMBZlbymdE7kWqivBQOUY0GTJpiZgof6IpTQzX+YVTKntijBO3c7P/9KqfBY5gR8LhG
KhQcny1HHJ5krWjlrWZoJTvIPQQWjI3G7vAO+z6EeB8520S0cmkN716JAwEMlkmUDB9VNDjptgY3
7b8/S8IU6TAqLg/FFMc0cv0i3RFm6aAK434ObQK6Uh6es/Wy2/jE66g+x4taWBC8dwijA6epSiES
J9VzOwt23G2eFjFYkG3TEZLPIMvdBQtQ/dWzPPNScekhHLLOrhg9U4X8tgyB5PBe/q8XisT+fG57
TP8RNAX0ON/zLtyNC9VSnR8HwyYvm0y2gdRNd7sq9+/xpWpq+tynvFNm0W3fkFDiFkFz8KLiZ/dI
u/fR+Wbutsh5Y7bRq1S0IrPe0LHj60aBbnemaXxJmi9+N48KApfPkh67f6bVXIRhCMbkfmpIjekd
mQIuLGABf5LUfKtCJbgTICemF4t/q+3pu0bKMu6CEbLl5Bv0URdLSz3cWhWVivT/JUEa8OfuSOWY
dh0TO36tDopXg3+KqxUi7I49r6ov/QhwptFKZfcyaBvNhLkiSF2aG/AGsj91vnFhzS4blc2x6wvp
ZVgtXYh7GUwx9aOTM36s7swm/HbdpSzP4H2pE1shLj9egtbNs1/Rqm6jwf1XCwWhLDkp/gv9Sc83
fCEPgxZoUc/33T8K7JpevI3UGL9vqRWtUQabdPBq1FZyLz8T1RaDVAr/OceouAbEXW6F7jCIiO2E
YlzTdnLcixpoflLNrpXjzRIstWsjgxyy39wnuDgFmCStIRzrUKhSxYMF62urqce6UlfDYyGjKabh
Yyb/A9H0cGDQ/5RtqwS6dQsNVmtRksi2XrJEPhj59Q6VFvrHkYOyuunzI8YceEBhsmysH8MpoyRC
nAMUSEGQ6vLKbg7IujYYSvv8Zw+9rMdiZJpj0KLTBFsfzKXgGhQeL0B+V/oIceNHA3yJnxzgNHNz
+3Bd40yls8lOtaVgrGYWgIkbffUMmAfmY7qlmT3FfChuIwOVlXYDZmr+pwvinbRxCJ5YMDdy3LwB
FBDjtrQaksH0wHtg1cPU+ocaQ2I43aAjazTgiNVZAIzzEfBy53DLAPJt8giRK7RoGZe+ZY7EnCIG
G4Bylcqj/bVBvX1pkl7kdMRn3ZqLXOEbJTpaEhn/6H1S+7X03mGMOhsG3bDRi8vLz567wKqmSYNZ
zR3EgJNtVafHjMpzN7RNkPbFyy5k2a2w1pL2go/DS3ACDkrvLvU5Zvl5bTagSXKTOlbKHWIz3ERQ
gbAFo/Mqzz0UXD3LaHLtBTG4Znm571f84+nG2SrAb1YgXlXUTPGjQp1w/XnpENT/7MGUm10vbGGT
Xmrg5ui05sLjBQq65P01pjcdDhgP8djfVIqujXteJ/0dvZ3AbLlfN/shbqeWXEQub0v2WYD1SFUY
b2txS+z1VN0U5H4AX2BjbIoMOcyx7UjMG9lgLkrHgn1XAlrbNX/Wf3B37o5b4OTqVo+hBXLZOfCB
xDPejjUljCGJRNmcPKRFLadBgQXxsqa7+GmfaCgbIuK1i+qoOlWyUwh1eqITbQmGcGyjuzYjzmC0
OdvQycgMABPpsbganzgqo0jpJcgKd24tgF+XfKWAR32DKIGTMjfoYb8loK3GaptKdea0svIDnpDJ
DRmnK0Vfk6yJ6TRpwaQLUQEdn12xxiFYEDn7gA6hygDxqzuA61zm1ItmW1MEdzBA2xJVWmQzmPQK
YkRDp8N5MmLGZCZzePCCJET6C0TAXkbDK9KR1vYtYjO68QTF3/l175bNXiS+YQP2EsZVV1UMgXJ4
hF1Xx0R5dHr1WT2eirwTFzRcZIf7tILEdZLFwVcE6ak8+vSvjR2ZxoAATN3x0LYNNTWQ4zbRpwdk
xl1T7nVJ7oCZbdU4Y0hRvY0x3LLRvGJCdmUQhsp6mI8HfF/Vi0sUxTFpORfjmMtyW3toNyqBPjkn
oIjhp0WZtSBvxiEWtXOgt9rmu2zYHy3X8atpJh8/bvUHz09xo2FoWGi+uS0reJRzZ7OF8QkzfoTa
uhxkNCewCPVmghEq2tV7elulGRqqfA6aYOybKlH4LRSzn3D0VHJyL+1vstysr1wEryr9EA50/8qI
DuMGSiPnvYOrCLUADBctWUEiSb91RUS7ioW9agd3hcjijvsB/zhaHkjya/laNAsTkrP/ebr/Pd0x
uK3KTaHRHhJuY92m1fisIuFXbdfbh7T3gG6HZDtRKjESOV3tuOWZ0SN80S0DFsJ/s2bo7JBgKmsE
IbRZH/ZYjyi/LCmZ1v0p4dOPvuuRPWRZeistMhHqHDleY+IQNRKUDyIi1vU9T9tJ0E9sJREAMCOY
pTXJUPhQH45qIPKu1dUYq0B24YJQWfPzsvD1dUyzUdBQYm885E9Rtfz7AiTK+cA0S31pg9paGJbc
S9n/mvPbE91TQfVBNP0Ts1R21OC1Z0OUjOY38TTJ80Y5oCrjeh8W3RWlX1vuYWMZoKgNi1m/lj2j
6DqCzX/cGJ5Q3GAi8iI0tDmW78e2JZewH4O4t7Hk0CowTrRSVqRGF/sZuMFg65XK8ahRHIFNnIwf
NADO3vcnL+eb0PNFsVrC0+da4j5twWHaCiW3Bmy0D7M4A2Ox5g8FyNPQecZUK7gEBgV3QtKhwy7E
z5z5g6IxznA8YQdmTeouS6ltwI7rw7coxi3jTT/vchRgksBPPOyiIBgVjhLphF5wPZNtIkEtsbgg
DVdiCTLxU38QBIGvncb+6GXttwRHby1ZgCkp02r+tTCS0DtRw4Wi3g0T6TcLWIwM2MzFe89MjS0Z
urFTkEn4zmyuAbwcILUT1gHhfoAIa5uvAO/+pbz/MWb51uZBpkadEHgzdFRGXnJ8D8ycvALSGx6Y
T3d1aPDQHdbXyPEcBGwEZ0dHxAwCFKy1zEcldYCRLxfn3oBJFLBxyVuH0cPyTY/pgzQbv4qvVywj
Qs4VIjYNsebwobZfLwbeE6+WJ7eYPn0aSojGpejmQ304I4mNYeelORCHNQ3miIyLztmSChRDx56J
aZBiYMTBM6HexkQatkGSR5Sv/OdTuKl3Ow9zUU3BUyOjRB4S36RnMChcBqibEYCPKcb7Pyfd+ixt
JLPAQZ40FCfjogPkBOvubRi03zZfYnNq4HI/g5x81/jKSLJdvKiqR4voPFCE/SFIhQ74Kas81kOH
7a2eXEE4MVloBtCABPX1cY3K5pwYXp8VJPbtkEy1kHgKQ1/PloitHKkgjg3+wRMaFQxLd62BHeqx
TjF+rz0pkhX6+EK8/dbx5SdH7sk1ph6gmDSIzH25jhFDb715/XIGiUD0XpMTDF/vRwnDqI0B2Bym
SqCiwzQYOa9OB04Ah9o4az+p80CpWRTNLDmbE3s71avmepArZUT/XoJVkpE6d/H3GKFvKGOSnXMd
CncHzkc8wNVZ5x5wRMgBZ2X1L+oWKgzlMKObtzDFsplaTKCfNbhAwa8mFoODH710cnMtFmUqEdCo
nQeDxqppZP/B4hcUI9m+Ikxk4LWeUbK1nWkVgsRjrZFsfDU19dfSyynkEbrGn9dDN8vWPxYJHgai
xf44BeCYR+C+M3SEgHc1PAFJrz2M3oZGGtiLNr76pmOL23q9ni+o6q+NkHEdwoQL6uo4Xn5BwRzP
q7RAib06RPN3xJ5ojL3M2kAVUuJiVNjbOulB1gVGEha4U7211EMelBLwOlAJmxOnXva6WWmeRiWW
zzPMlXaNQ43CKnX1ujW7g+pe6CWS4ApPYAG8MOnENVlejzDXSXRohWVR1I0vZDlEnC6xiVoiRVoe
IvErnAC6pTG0+LF4JBgl1GaZPIA3gDq5psdgl1StK2Yk41dQ9HT5OM/Ieffpd/Df3CaCfMjRK8rg
LdKYNft+aG61+Yg/NXvriVKCjYDVgdEOy04jNozJZoYZfteYfWqxd+e+qjUhQ9IsgTq20GGRBtSS
TRpFptjorhKlEcFWw7AdEtaMWcLIrX4cJA/DSsQSLW4dLfTRnZxy/ll2WiTdBAnIFS6FYqkMshuW
Q5Ocp1MvH8wfHRSOKAe1wSkadpIKgdnw0ZLA/qjCcapqe2Vfyapfi/RTFkAeqLOHEpKglA8W4Nve
4U+I2I4SzBL8UI/bmGwuMzu7BRhXa+j1Au7g/n+kiD6sSLOFZNIdyE3nfRN4tm5VqenHtUGYNuBy
LSy925gDpHMzzt2I6Ut6sSw0VauDdGQzCjYT2feVIP41R5oPlftlb0CtV9QIGcTTJcmZCPQ529VM
Pcqm5lYATCV1Qt41K4N8v0Tr2NmTAyAlP+ns+FOKWzAghLIVV/Rg/awvTNJzs8aOcol1eSNP2eCk
XCFJHpGQpncYsbdEaCUFaP/9BCnEJEgMxRYePyIkWDs4guUYmwJb25XiXHatjFv2975lYboviouL
zQmNa8mfA9V/k6hiumHWrJQxYBCuYS25I4Hm2OJimBN2gB65P9SnDu3WK+gSSN3B6+YKr0G/aAki
JxspmxG+m2odoFbpxRQ9toEzKLo25ep/x+ZlI8vXpVfq9BnHAy2AyqrL3TScgiDFYAJ/hpOt+kr2
dLN8biAt0bKck/lu3JTHN/izIolZqGExeEPzQmuKYZ25Okk9MqbVdpI2NvYYKfUcZy5cdPJyVChK
zn3nVo+D5s4U1KE6mOQd/+CpE09ohor/cKPoHpqSYSzZJmJXrxm352l3JGbQ8HvN5JbEtsYfZApQ
wudjzV+qcCFULNwig8Qpkm9cqPDduRQgG/3SIsiftqwC8n2+IT8D82BrNgWqbFjJaKAtNL4f5P8W
19Ru5sv/f5n9a5KNsj77xn3H5VQEQU8hCvbNtNEMr9yR6xHqCivCT2ywzQCGZGF534a08eB1EsZk
08TtWR/1a5U1lBdljnO/7MvHPY805hlpPjfzXrBC0wrowSi6tGvAYNRVUtoal+Mxh4KZ4r2/7anl
E2rYf2aX1Y4+X4pYpI5rZ8vSSOIlEjtaL/6SZGgk0U0XmfpKajcV0zzD9BjsLCIp9RB2rSN/O4zr
tPsJmGP2LN9z4I+Ce94kMwTaKTwdAg3MpBxKeEhU5CpU7HfIvDwjZB2y+ZC/QRzoCBxLfI+M6ind
d85kE69asasb6a0g1zjGYj0YeLs9IeyXcucTERsyvyP807TKxeU2sEpHC38nFa4iMXxpCq9GrwSu
U93L7KdvBLtGOpg96DZtnrG4iYbDTJhNLm0q9Yfc9kLDCO8cX63GcilqQnbH0muBlaJ3VzIAFDT8
kQGvrTtz07dL+zDNulDd+hHegTmJt+pY9n9F96UuyZd89zzdl7EkpxliYNqCAb0OCx56x0pYe43K
0O3OksYoboaT8V9LNHplAfeo1CquYbw9Ued1SNComd9rVH+WcwpvxJ9GOOMwwntpOYam3RBiEZw9
xRkZT/cX15YUrcQH5W/hTDFW7mbUdkXMvlqSXGvoS1sk76m2DbgK0fpBieuyTIPI26QBmfsaVqKI
E8IOOsXKOLeLIMvjFR+btr2ej+RQvnSmLzcTDqw3g76xcgIaSFdYuMavi4AaFwDb2wpoT/C3q/l2
RmJ6Peqs9xg6t6wgX0TiKVsApuWJuPAR1kc0qReNyPkG+7FROzrBNDEgCn+G1dMr7m9jtpVu715n
bL9QMi9UQsO+vesrYFgoqxX3wdeLSRQN+rsv/iwha86QDYnfCZ7oee4X/LjWuNeeRfJf3rDzfpe0
QkxXir8ooQgk7td/XkTqDrxb1iMYptGyOdQ2zmWJ3i6qGodrg4yAb+YHb3b5fcOIsBJriLwIWzvy
DK7+LIZdcTtkAmHDFTwboopZknFeazi3NgXJcDW7cQn4r4LF3Z/t905qo7AVk4bN75HwJSQMJPNT
LOsprkOHXF3OVY8swBoi9i1m6DvYb/McZTfKzZZEdBLpprnD8+Oel1Oe1W0ZV3n+pFuAaeWbSNm0
ca9AGGj25Y+4lllebCDWptId1Xw0yhxmhb9FGj+Uvg4JVU7cyNdEKlXpx5Zi0lCxCp84tFA2uMuD
JzMyaaiF9PqArOrUGKU/1ppSPTE1K2VWyiSrFxZ/f3ografoSGEd2Qs8JMKTORfomF+UyN9M75dy
Jqm9g+nSn0EUGPRCyYe60onJ+NYWOiXPtZHUwwCXPoQfqoSjnAMFrTO+x6OE2OMNSKr5faSIm+H7
hdPlvYcMiSM3+y3nmTgeUHMjhkQtLWEsy5rpY4ijJbs6poK1mRCg/KY9xygYY0LkBQGxSoUQnW5H
OXpzo+8FNhhF+HDKEDVsDh5hnBaXESxj33cTFjufmOiC43or5FPvx8SLeb855jwov7sBl28TqPWr
XVakemMmoWq/HPwBfF1RnKFC2UkqWIrZogkPgDPyzj/nOOJfIPuUs4laFP9N3jVjS6oYpf6/93zd
OoLZcfL+dvCuYng8FsqRomXnoCEkGiaKjRIn8wZupWViCn4ASNeESoib97/gq2Ujn9wlV/yiWpyY
uZrtejIAVB+SKTYEG6HfD1HK44Z1qd5dMTvEAIdHZ3NNnqix+1VjMT9SxgnX758R9tTO9/QMhlfn
U7cCeeac45+d37SIxD7iW2NhFB4BIuoly6VbqCgvSfJAWdaKB/wuxK9P/1NdRaTFM/YhPcDRym9V
z9WPMOrh8jJuMuQzI7IlkWK/qa6I5Wnc/kOgyYP3HrhJwwHrt4gVQV7Kdr+RK//xRaVbJyUSRnx/
9E3xULP5nT+KEBVppagMBMRr3EL+lMC7cghZGdzECI+C1SBQEzgYo01RV75ooIN20KN7t9gvdUbi
jBPDcR6KEPcMi6uYlMfxKnl7wYcMkB2Pds6rwPpa/GtPcJT/1rbFWLQ7l+7IJunJJdeXrR/dAK4S
lSFnfbwHpJQYm/nEDt7HldPFa12vm9VkS59eYFOZ3/iThym9mQXFLygBXzLgfUd11y1ZPx4yOI8F
R2I+aWPZH/rAHO/k+kd9sQUZpSyDhUneOAELkrc7mAyvxvcah/h1D29fL/yNTjy51fbE41zI39Qk
6kMdfbhppNJp2LKmzFaRbJe22TwzTeDc8ZE2EF1ew/4oquqYj4crasEbGdkzPsCtqR1X1JYuqX9c
Jr50IM5LyhjI8CVerFl5nh9vTuvNr/DDnd8OGbdbH1rvJu1RbpBwi8WhO0xM2o2MBNpE2rt5CbHe
CtH6y2YtFvUi+w9YoWiA6BumCL4fdAoLaIKHX2oH4EQYUhR7Ls7heW4kDAOvaFYBjNCr8v0MUAYp
+tRzN6HEESrjUabQZYHzFMeQ6oKvYz9gLKVU34u0L0W7MAGbL0aTs/QGGOznJyqkj8OFlbazoQ+q
BICxw6c3I+s60kzqQ0Ka5+anxoUYzb9fFZPtyIX4JPI2vKMxqUn2xK/eSlLR3B+YGseZN1JqCSLQ
vI6Pf5nJPwtLcHPJzEYKYt7JANW8eVzQvdk8Yx4xkBDkUhlASwnKreVrfOBhos7OqGO80rlDWqkF
dvxyhxSaxtxA/pBaABuninr+j5zUMjDQIHkEpU/P8r4pS029ppxZKywdnHnaqqBpkHXce0lUw/he
q6oN0o0yvKVwlQdP8lSenFk9n4l8SiTnZ5EtD9oTpQeFRK9z2gmCThjiYJDvW8I06R9Swoq9QNq7
3owxgGTxoEhPVoInE1gWsJOkfnUN+ErAy/LiArE93syIC2tJP+Wk95Fr/eJiOkzjJVzlOFlCfINW
VVgAIVPdcAJD9uPttFeEWIyTBlXq+g03moZ5oNqsSCe7uqBbjQzgDy8btraNFvzlYvHaNXKF7AC+
v11FM7aLCycyi0KvlsMqGMFRfKV/27VwS/05QeDQPRwpY1IWWWfF6Yx68kpBWl9Y9J6E86EH3Bbd
jNU2IEiZM0oITkPFG8meht+ODoUBcrwL4jmxXGscmDrSotZReS96/QiyPeBAWYGASE2Nw/doQIxj
+yPwem6UAOIMbhboch3lEYhmELg/x4cnCIB/paYPlEKAMiESj1cbjRwqE8y9ldl7oDVTEZLG3vcw
deX27Gw5qHJt844+ymDQ8Lw6ELatIQkuDB2TtwVCtwfwD5s2/A1f9t0qIPSJRfssV6lVwNt26lUn
u3SD6bX1Lyx8FZsR1TIyIQxJbPgszGM1v7fPJuaFepNybGhuis61/Y0T7c3A5v8lHdjtH1YpN3lV
rVeu5Z2bij+bagFVXQgS9dPp059fNbPIG4xdw9L0BqkwfHLaAC0Vupr9VZgncaNxGejpYx1ycsbz
kZ4zgpWffSppBlcRBryyhde3YOTe0AtERfxG2lDDVz2R4uhKlUTt0mDLGxrE7JJbk/UeLHVWMzU0
x9bCEkW+6+rue03KtITrJggh0jzIzjzuqKgP0d3MgZc0iHjJefFCQpbSfw1zfw2J0GjxTCM0Z0Dk
EhCpgSC0w2WWGb0jtRRbl1XbuwCFUciVdvn6tKgfa7OmoAZsniPSiZu96DBbgp50nVmj0WciJju/
0U69IFLtTODWKKN/qAbXfL18BHuTvKI+2YYIZl3f0x1EJAc9qVHCXpdLiLlZWaHimzIpCZjXFuB1
Ske5ZE0Bh3HaisQS4EMscNHfn0OwH4un4kW09z3En4deV8YqjFG0JJMsDP7AApRv9vCbkVX5jKQ8
PJ5+nPUenNI94jboVUjTeHTAGP7o45nXTXFJz13h1FX9//boBFMirzwz66yh2o14VL1v1zm3qvNx
z0HFVdxt6oJKUaiMds5JjYDyWwjr4UsrWlInCzj21388hY8G5GoJZtolcP8TC4NZYPf00IJcbyfE
5eP2Ghklk+e79FnW68SeTEVHdeRU3Og0aBAtO5H4FC74EW+B0NcI+KnTg+oMIHmRl4QLP/TY5Wku
jskUR2LeYx7JTjGIeaOR94yTVelVlAvs9Ke5HLbbLBXnzV0QV63RC0Uuh6TVCPy4XB3geKmB34T6
u0vBvILUheAOH+ZV20YGcZfZreZqwsVg1gkHMxAzK5JlIYzfrBAiMqkB83qPOobcgnFR9StYrQ7N
ztDOkIQ9XvXPMziqwmN254o2wFE1SynzITMiFTTDWYcWXc1/RYL41MoX3DmwpcQhfyFkZSroG9eu
n3eWG+3vhaQ28Q5f6HwgrmZUUs2x3mjKKy8G75iQAOhQRP2tCeyY03jBrKVc/Juyt+f291eoi1Az
aktb5UxmXsSbTuqDdyNWM50QJYwCZiXN22WWksqhCMeDH91bimbc+DdWW8oLAmqXLeA4rj4XVBBU
eGGezWd40XEFjv4uSd7aWi9dk9wH7PwjhB+rAxW458bnyioNM9fKVscRAZCny1eBJh+WShag1liz
XD+pfco5d7dxaAPGEyE20uFqPKb+jDvpqvRK6Gsa/eXbKZCt6xodGJjeoMOWR9fXrcIXT2iOZ1jL
Iul8IGVmBOzmurrV2oAsboYNktrjuYiEO/SXlD0UyhVoUzyC83938geacxFe51nT4Juv+/mJezSL
uNGKJw3tAD7sVL2QK7Pz8PxnKN99cfuJWZ6tORwgDuLxqJB7KI9fTs5m4Y8rqv/Eq03PrdxRwUZC
QAfw9M3bpGb9bjKn+4AyZqDRk3BO5WjyCtqTxVNF3azvySQcmx4ATj+UPWVB8WxyoSqNrDLbWOXM
jH3M2J3nhna0+juzqI7n8dj4onP1X+T3/SzeOdkUNeUgC1LCrtIL6cl+rskDJBozKPZdCwimmG9w
xrOe7OhJlnnggY+dFJrFFcggGpLD/bAWqKQps/LLePp2rPIAi8+XWzK8QY5pSk8qJb6Dt4PLwRwL
bQXJdmbwA5nnx48cyxlBeb9//GH2ukPoC0FUktz+Yb9s9aC5OVu9R0YyEGlaSal3coPgN6rGxxle
U9FUXrCUFYmMI8+l3+LJopFUrZ+/RKLtvBg6AgQUGXvLR+J1NGrDCKJ/bQxMmHbhxBHRMVHdmEpb
IMYrviEjfO2uvJFnFQiS0naepLiy5t5W8IBJaSBq/uGYVyrdDDAIHIeNnjMS/3Z2V3UCT8lSidIG
ARr0m6H2DIZxZxsEaguwvfNGPPUw8iYl8aE62bQgP37/G6iQ0+PPtW6MbrP0U3Xm7Qs3OnoZQf8O
ThDK4iY09RkWS4OHdp8bC7SK15VGNJZG+HGJaP35K7J8INNEaXanogjoTFgZYw2TOWSqn1L9hhSX
UkiWQFvO8HgkhqesOORyoT0U1zawd0xWaKuKzjhIFlbX1BvAV17Bx884OFf5h5qo1gGMpTiwJL2w
erATa+Sf8NGgmy6sX5gLoYVXjZLD4Rd2v5hreQZURofPTvve4PCrHUsjgzz9dEK5P7A9xGaF3fgS
ygK2cldKB7t6iM8v8nSZbjUFSys4Q8tOrRUq9dIU4V8L0bEif6KHDPPJX2ulLXCJYGVh+QPmKo/h
JoiN0f9oleykJvlsruCPjGyfiNiDhfI/VJYCw7zz/OT2RLicK33skpD85ClVYnl7yKDgeVjr/6Ui
dlgBK9qw8Tn25ZPMk10IWHO8jFlwOjuTn1utACU5Aj0JPKOAC43BtAmAgZZ1C0jnEiRVJHOJr6kS
sgpqj5WHVPH3yyY5Sw/h4UN1KEUlrKIggYXqmyHiHAUan6tc0juo4WhIBlczMlAhbRQsuJOAn+uT
yI72rUEkl7SWFBGovDN+tDVB4WjIz2GtlZ3FXdvpCPafc5L7tW9dcbMq5XeB1z6n7yV5Eq+lZx1L
9TfJDsitstrTfJ3EQaIXXyKTBi+81dBKrwYRW3jYNgh+qr8CkeQonl/2kcb9lvLC1xegN+c4KFdo
cj0ODipVBxDhlQAPIcbBPzSW9kg1SNvaGFszdnJmO95OXpxWhyscrcaT4lCNgauvZwgful5wsbK4
dWdUQT2mVKx81dr63b+LzL7Y9Igkw9iVbUNoVDlovNaduOFeM6+HvLrAOSEz0SF976oUvSzrEUqe
z/Q/d1jTOY/ZIH0cD+PgkprXRi2iOyiHMHxb8qjn+qPUdAdL4gqOJgDanq1W559rVx0SOrt7G9bu
h4XcNWYnPK/EcxZ36opBDweSwNlykzD7KC2DGYvin4qmmD9g3vZulpt4vzxe5lDhanQSLKwa9a5y
LsgCXaUEu8ib8boyawvEp6K6hPyIdHCRucVWY4uwHf8RFlNQs3cs3L4tsWCDShF4a/XXSTUhPhEB
bw7kcdg/hKNOdgRfoeS5S+JoXN+gSuOrsnRQnYo2+W0bm0st6tz/C0jm7p4U5J/fnItUgDI6OKDL
wVgPS94Duqw0AENf6qU633fVpUMuzuj9eLkcESgFUH2rGiNjs3SWfrbWHlMhY5cjTgxmBmP4mUM5
5DKgdKdV7nxuBwfX5uI4/Ud7o8gaqmv52JH9b0cP+1jRL+PgK//4iB3sXfEDdMfiRUxbQQ4qlHsf
/LmYY0r2oOcvwaUL09BUh2yAQvmLS600OHophlYTmGApaGVv5Bh7lLhLtugkmhGa+jeWP2pIpcb3
2QookYFeaV2EFf3lA/r1qXsdvEGDP3vkiZcJpQErADVvS6QlR3u+jn060Bl1MrcR2A3kslVLY0iz
9rsZ3eCwzTHfILWM/EkkJBRfr7vzGN5WJk2QcQRzlXaY3OyO+hURMcrNpV6kOhEqNgellxfImG7o
TxrEKK90ZLFVy8ocIH1EIZnLBWJtGIv7gIY3e3ALNnMSOGsBb/tC4G6KWOXpVKQCNHjbYmZ/9PYG
V+BWBkG7ccj9+vuBQMHaz5PUS66kd/g/mW5KVl53BEri27JWbqeOMaB1Gq3WUeFsXZA1eTm2khkw
M9szP7bCPrnnH2RM2WjncYgw325klBNF/4R+KBP2o7+bjGyKsNP/uRBjTI8NfzlIYNCnayvd37ex
DIeDP92bBCHvCJyhhhW74nBWKoqj354+HxL3xsGBNgqQTXTEC9w8wE+oqCtoCL5F070s48/nSMaH
1BhAXxyqtdn17hHkEcVQkSyb6heYPVI9Ts9g6MM8n62dCeJzrTnUjCjnOeaqdci2bYqDFdyxzJLF
18hLUgfn+3lalDKopP/lFyrmlO4I60R2dPlss5nl3RVBeK+LS8/5pjNB57ElS5h1gW5mD1ekcE1P
ze1TZ98aWIvEPw0M7g6+ADbBaf3LKVCYIcoJxN/YvCaeH8FmkGbzNeELrOuUHW22pCAmv11Zn/2K
2IkuvzyZiTTLVF9kJgoF1ZVUZvP5afE9Bz1EfPhvD+1laHDfDioqCdNL0bD8VZnJPmzAUbEzQApa
sPmC9/EFR20Bk9MVID4folcf3zhTVpCgOesRJaAQBEo+Hlb0BPJyZCzuzR2rrH8TS2IBmDa1tmsU
doOpyshVSbyGlHq6Co7F/Au7O3QEe1M/dPTHUDn18vE81IQQriXMcTp42I31JAAfakiwHb/dkbVm
EQAtgmHRJVZ8sJ6tiNRgLR806nmnCgVeziM5JKp9arTW81EinKrQpT8JKht1caWcM+4y9F8Utx8P
wKppzAZDagDIYoNSlSMDxVhkZU2kIrT5jID41p/V5RgWPWYU8Y0bVcw6YgtlZTkTwW35YfHib+AT
oBPN751pmbNZw8Z1DDS6kCebac+9eGaKYNF1W6lYGvFgzPvadbKXfiN+jLFTLzu/nzxuQJ7KtZ6k
ZJiWYxxkMNgBRQKu3hfsx/0AWbE5KE1VVCK1pcfJn+yAxCfN35CI5QgJs8MD+xUZ7kY9FOZuau8T
wbyiJ4fzqZ2egIVOnwiYI6K+QPsgoHrug0WysppUoOxEuud2ePG2J1pl0eK6GGWNPIbOau1TjGsH
jpB5o7D61Qzw6hM8zpJx7kne0gkeoHU3RV+sXqsB9uFtFn35UA20RwaXBy8DRFOSopp7mAhFQQUo
OtHBjQd0p2hd2zKAjBhA96adZVTlE6XCN6JxQPwudw1hVwrl6VqD00b2OsViUO0Xvg5LMYWaKz85
e7uc/9v6ZIKIzaZFXVwsPN3ysJLn5nJCcQ8amwSKz+Fqm+kTd4viDHGeeWArOYgrw62yVcbIlTVh
eZI4hXpRqozCzHehrvL6ZnM17229rZM5kOBT9QmzT7qF/H11odx9PCmwf+qS3Szs1AO5J7yNozGA
xKpTjGDfofn8CKpKlPqAjUbq/a9VjfjFqrsWjoOk1yPnWD62JWKmIc8rDk8Iox7wW02o9rlR+m/a
+rWgKunYXXedbfVTTiGUNoSpnjvD3wjoBD/3hzJDULED8FamyOTlSQkSW0lJZejsaG0NtPTo9DyM
IQ3qJNK0sP0bcc/8AFsP4W6jRzx/zH40uxO1M6T3gEheRBPOtB9kY7VL6IAZc4qRe2oRFu86ixZg
xLxGWEurUTJfrDeDGwZp73bPzr+kiSn9bBcNmVuJo8a47GrDyWBLoniwgjwS+Dszltx74m7IlZmT
WXVZf9Lju+Z4B6+WQzsgTcyPD0DLNULE/hLb1qCG/BdulAgpDWFfcF6e0y2pjSSvgdy2FCzV4wps
l/ZVw68hKTEOCO2E9g3JQCp7kwSjI4dRtfk75H9V8oits+Cb0MhrarW3yfSL3sxFAtn3n3NpGlm5
/S+m6lKwIQIpJuUTS0WCYaXT47LNaNwkW1+Tmym3OvMQ6+m1yX2jKxAUXQwUIvBen2/eD7TadgMS
t4VnXZVmK01FaZQly1yfbxyXgiuwvEWtvipqKywb8eA7MC1CxXUu3v4ENiLTuBsl0IUD81Yd7xmx
BIUhWy3DDW6qbRQTPW03xHs3uOAXbxAwDrM7yBnIoBgK/K5TmonVD5HChaKBxhNUxlNJC8Nru5sv
AvE0rSjOvZqducMpzOgWBwE42WR4/yvr9983TpZxG/8v+gkKYj3mA2j+nQn9F5Wmzu+6pdYF7nn7
cf4kV288z+Tl/pDwijuKQ+TR+B5HpvEf1sQf1GBC51OWVB9LTjtm3gvisXkcZs9XvMNLqkr18Z5g
74RzQ8YzVqb+H2llB+sMyRNWHp1w8gmbskrLVqGzi2jU/usC/wbC+zDuuF/SgtG6/1RHZr074X6Q
vujzEquFVkx/E+FWGLByqK6Z7n1XQkH3/9no8W+8+eFj5sg39fYo4n7vd7NAjYdSPGv5TZqbvGg0
354UnjzQ4EmgKR6Tgg3R1o0Jiggk2ENZVueGhGDMKLJeSivdNt8MoWaUfvOZQ0pQTsutV12xwt5a
aX+iIc93GSf77VYnJkDqEtZkYugw11XCfr88bnjKa8nV8CrbvtTfCa2geTOdtGQ5f3Diy9S0gZZX
zWTPjznF4PF4/wnlr011PHvBfWRtGs5BK9LG8QnAFgE/ccJl0ORv0TBfMyLM3lG2LI+ulr2d9Ib/
mzbsM/BUcdyD0fTwiWAicADAk/O3k48IHFHAfkI3EELl6+qTbAwIx4H5Nd8vKY1Fd+Nd6FcreOuz
N5BQBpp45lC2PDorZtqrtVA78hC/GaMi9N7tKoWV/BtLzRVfXb8f1iKmi7pi5scBclSWcyQRlxJs
9gHZiYOolVE7VMBCan0G/zvT84fxJ495M2EEvNjf7ogPi/sfN56QpncuyZjl2Dtb9Yg5E5pVivH7
/WG+BEcjTvOaI+TGwmBlgC744sHx4xoazHrB7imFmrSJIAUG4tRwICLD0RshmlNUPCC4FNQjajln
D4eeIfiGn/WeXp1ep68Tgcl+fi1Pu2yCNOG848RHbVI7q/zFK5/WzwvR8dwLcfFG0PIAookX/fMP
IbcgOgJ66hHMxLQ7C38XQqQvgsQiMo2A/EAVIN4PRRXLtuUwqs/Qm6BATJFZLSpmx5WllP8ISTv4
Ag1HQZZTNVdWB6th4vMuBJSN1H/lRN/iXmm1xz+CeTyOk2HeXd+0jGPXV7FgrOz868iZnbSt+mN/
4N2BSbfKC6BZ8HhrMmVKQEQWWZgjoYVDl+/aLLXLA44qjmtCugub8STgmn7lu63KVcwWjkIpY+4r
SV5382AojCpHYaMMnkbb+iZBB/1UhOm/I+5VTPbSzbnt3hWEin0BHm/+mK9rTSJBNfbv7sL9uDsl
zhXzOLvOgvkFPGJQ9/bT442+goLDcY7K0T3T7pc5QXhY8D2hCBhMGp4+9cLkPNzsqF1JOInBpcM3
FtGP076OhrWsE1ohLw9RFzEf3oK5HwOlhlJnbGtesU3d1PNb/xIYxG49NAqnClluD4xVPjbtvDmH
uXFOF+cFQE7G3cn3MngnHzVCEc9vFnDg07Jkvz2gL7XeTzUaFlYB3p4nJATflGdNp874cB9M7zoP
S48GyIKdbz+q/qfLws//2ShUU+3LaGwmjU8FlH0zfpEX+lMFBrYFU+p9KCnNWMFOZWP2vxCT70eI
MAltmjI/TbV64GZjM6cDPJSvREyXAaKmOhBoIXC3dEdfkR2zJMANEyWNCABZW+kRh4VOGXoq6ag9
jxSUPadgQeCmRSln+j/eN35pvu44kL5eOPGI8q8EcKhsQBZUy+hpPhZKtGwJPahx3a49EAx1Vy41
2e9b2XFhH17naa4HXbZeXV8A4p3dBReRxv6VFIejgjIvJFzw9phWjfwBPgJ9+RrQkHlHD6fD5/nz
hh/8vduI267WDIMPZd/jOumLgIJTWl8KqI0cEJDRj+V+JaM36aC5hq9ac/TImpJY68JGgW2JjK3I
zT98VakK0KT+JhUFUIjhN2a34ZQmose/65BOJx8qtLNq7T39UQlanFJuVAYz0yZbrTSd9HfRLRZ3
470S9v8O3Fd5MipNXC65x7khrVPzzEFaZyJRlPk2tQ+i3JcgS1hZmhAJzfdz3biYuloes3Vx5j/8
6NelR6Z4IgYtpoinG5cp1GpwHsF+/GA8wNdMikXdy69uQ2nq19jzoOTyJaT5m1VLM7JPVsLmEmob
Iy220gFkW+k2UqBJVLms6Q5nwOb2zclI1Cx7kRK1ePijxFq/sB3F2HHPQz9ULQ/TSu3KnXPWglpM
ms+wFcTXtPGwdlgHnXPuD3QFbzVfnKkiTeOgUN0qsXHb8ZcM6IA5/T7Xm5z0uXYjmXT0XC/oOuih
r+IWSNhSO/8Gk9SByet6Nfx82Dd0Wt0GaUVDd8UnckiuevMcJ3iyb2Acg41kt8EbqoZrALzqAUG2
Xt1S56I06FPbf/DPPXdaRTxuIXPpwjXPhVxCRGZFfU4NGtJf5TELwyRl6v6GSxiixSip8tsoDgQA
S4z44OnXRyz16h7fKZzuL09W6vnOIH3gBwM2Q3HAUkVkgGXhoXJ8eMDOxG+HAPRc1tuPTVP1rv0q
8ujDRfMTrV0jvqeu7FzObFMkz1kaguMgyacY4K7ikDtT5f5G8YAuMaM305cWoHRSPOyPdRxor25Z
t9x9LHw4zMFAogmFKDNZGnuoCUu4zrEw4v33tqCtnRFiTIzJHWpkIWr8YU42s2sGbgsMhilayijB
k8A72YCJmD3MD27HlAKCi7+JrBGLin6tEu26Co0MTK9ElEvWyXO4JJlHfl8sS72MTcgLo923IWvB
ZEaeM7cRPPRcyf8r2s8cZWUnYcSpfHd/gvlws78BmXEwChzr/tkjeFZnOHSyaP11biBLWO6k9mpl
5XzGlnf1TKbY9WtLHlDyQUEIZrMA6H5Lyo0Bpzq8pSZEGB+Tm8sufGkZvZoqQleg8H+Fhxchmsoz
BkqqptjKBq9diQ3sfFwTQqcg2+uIYU3F/vDWxOht6egKt8zDRM4aqOuRn9kwV08r13YRyMRNR5Je
UEy/a1XmBm4qu+9Dm9WysGTdrvy2IPI7V7RteIjKna95hCwCnCkCW6w2ysT8opXYDG0gBMXjqydA
wSl30ImuIHCl/ThiGu5tPX1cz57OX5kMtI/P0Cdeq0tgguzpsyDvl/eZJyXjj/JzuYeAoom0FK1r
CNX1JbvOSuKjIi/9DQWR9jsXq7kq/8B5HU5d+HA+6v+Lt69xBwyjh8euJ/lmvfvLCkW40X2+mZFu
19JvS8OxvlFXVqe1gUxtvRupGH3dpwvHqkxdlBrVX6D+E/9eOtoA/CXLa7FpoNuag5drhINGe4ar
XvwtfROubAllSGfwKA5zoZUqqVLl6wYqYmO5PEmU7TP9YejLOhz4BnpM4XCWnO6xt/Q4akr/wIXp
Ury+ZHf0yWxAWFUBhqlK+S2JPvELJXOEzeaFN2VmykP1UTtzRYYzeRlNrfu7c4oz8X2D0wSsZ9rv
0GrA+55QCZegNOHwbXIh2CiIrxHTliwFIOPZH4Hzr8ZMG8itGF8LGTMnUowCI/RIBBy4H/dXSikb
ma+xXr3myQDMi9lis3iMSmzqJiGN5xb5UyQFo7GqFGUOkUxU4O9dyEKGxb+O+oEpdfK8UD1DX+Ie
K4GXxwEPyQENsnGobBGxsPNq1MXZQ1gTtpLf25vO6XNpDtdZH5+C6Qya/ePJHC+PxFQ6PlW+QY+d
9Rm1Sg8Bt/fVKHF7FDLAdEid3pT9S0jLCAH/+Pwxlyy4zhcb8WXoacVhINY6bNBRh4PyQ8KLzVeM
G5uSvpbXWTuR70gD65SOsUm7Aq+/vmkP/mWja3qgohBCkAXvKPd0PMIjGI9lEOBGBnfh8Ec7SOKp
E0hhFHVo+DRdDxmXWyssHVdPpTJvztyHpDgV1vpipQ3ey70yYpikoUk5mrD4undVPsp9qFAWXj7A
Cm8peybC6Vqo0e9JW6q50AEkqZ+ftQEJJRHz+R1yhZeA9mf+NibLVbHLbNB9DwQ4GZNOKMbxhvv5
BSFVgUczY47S+AaO0tg0JlYT/ax/QFoI2/HN+iOwjjZklEUW8Nbscnl+qKlNVvncotI0TvhVQZLk
oL9IhiY+iT6gmsKLyHYKYGD18GNFhsMe2Z3VikZhSIRjQgAnL/M5HK7y4dx6waZWcM0aYFvStflZ
7c+wWNR9DvVIZDPbX0zsFTbAh2OH7ZabQKI8M6anZcHbvNLBzaRzNmxwthDTfwlf5aDjxn/G6B9P
SwhZKYpZj71hKGzDDMFyKvJLsr/ASSJCL5xHJfGy86lDV9D2P6S15bFD6nGHvFCplC15FVfYJDfU
X5PpBYcIT2tOYz/Y97pSWi/cem8ylSMdILyHhxE+JL7MCY4wwk9DOH2bPlzVqwjPGoFmJbNKCo/4
4OirxooD4nPKag5PfZYETtfB5+eMcdpYuLODpDN2by8sY7HkRxPahYeP9ucsRZ5UrBACNWPjFmb0
K2MA8uG957eOdqk8IOohiSU0PJr6A7dWZYu7QiYbeMRGL1avWKjAdM2TQlDe+PRnvo/99Pysbcam
8y1kwJcc1rG7x81QSvQ5IcVdVmhFTuPfRI8/mNdCJlFH4avH96KThT3PYX1/RaZTUiSz4l74YlZb
EZY9dcy2F1/PMF9xM+4IjBUKiC489hE7xUWoyKAn8HK53Yi/+Da7qfFlOdDwDtRbBMw8Hq3Ru1uQ
HdLyrQZKed/D1432AZegrFfbEMZjCqkzLldNvn+WY4gIUYO/3BnGd4h6Bo3KsEi/NvvxyYwPBsEW
F+faKvDg6qNWMBF7kkafKwGkTKOpiZNNXXIyR9GaCe3T3oMzwj0gXr7xb21YH6YyIehM6lnD6nd1
sXLScgb8L2eff2fsgCh8SrVAOi3NomA2uK6tgnXQyPCm+JuQEkE7A04Q6C8o7R9CES2sQnd9oCNO
2kdITyZoNUjO6k/aQ9ioKE/GOxnBsKlJVYCUe1dwu8rTq5ad63uuCSglI5OLb5qy/F7uZhUAutXl
AjvdSwOYiHFcKhWL5fuK1bbrwZ8bfdWydJFViTwd5vn2npW8EBydhpx37lGBuO+t1mrFBm/4Ro+i
o3ElALJe+SMEhhOIwxt6FbyiAvdzXsnIKp5vKAp49c6CV7kY31ynB+37Oeg65YExYDloV4Ddxnzn
NsINgk04D0qLo/dAvEgeQLD+DmZH622JTh7Yr7/ZmKEOG6NQIZJATHLKfUkC/nBYNgRYc1Qvc++q
GvkgUb2Z84uQCpzOMO9nJmu/nFjgTXZZvuVbgMJvkLM1IzSm0R6+bajnx/gsQZg9EdegpVGhzIyM
m9gFTsuqD02+TxSMO8UN46kwr/X1FvzW60sqtbZib+MM1bzlqshNftoo5NVk+QfiJCDGkGdKq3Rb
EFT6djJcCMi9HUYcY7HfxcbYsAt1GEAF9ZA1BiUZkVSEwFt509rHbNoC/0Pzj5bz6ltyQRsBo/Ql
HGdKL8olyXb6+QRxR56KH9EQ9NMOz11qsMTywAyU3mal8lGbm6fdeq8AVFzdKoPHftmtoGn4e+CV
v/AVrKMlIaTTgannDNVdbu+uZGRJiHPWVAsTQMKu2zRgz3QPtoX4uJ7rCpWcL2bsbs8bdm6sV77F
SPyXEbE7z2y7S6T+HK6kAtuXmOdWwVqyN/10cPpwuGVD9YFtPSEIhJ+OS/jN0AAgprEDysdCRpqX
AGg6qPSckJ/YNuT8WpSAU7EuHGba9jaLbd33bRGCWF08TMo2gTHYfXottVKO6P+hKdKsk5b2lmYO
zOigov8sq1YZiYCfz7nN0ydNoei6sgAXV9kryE+eimz5zt28qKAtsvBUjmRcZ3NuqgsM+59+XoBN
txt6DWj+gDFx3nHMrzd8dAX7hn3LJHnxwi1qxL41/vo/tqIE2ExpUSbiZuLCki2HdiXwOfAElbnH
A75SdlU+gzOcGjEGfnsBwHj4AgQ7TAF9SqThRLTA4EEtCDdszcqRyGeQuwwkYLvSJmBKp8ko8y3f
2VBs4wjo7vIceq7cp8ZVdtrrLOEKZe9U8Cizs2DH9I/J1FQyz2QjA7Jqee0VrrlpehrL/h0IKmW0
1IGnQkXA1eFahLbhQrw2BaEHcQfSYi1v0uJg+AwogXJGvbkhYAwJI30PTz4J17ocXJssC7oLmUSd
3j6dch+2HXu9ikSUixihBZmf4sT3pNGgHmo3eFvt4XXovj8islM6M2B2m0Wn74TWosxdwIoSYzO9
rPtmYPzQx6C+IvtMJ8P70S9U2zMPAbULs5i4ijJMbd2QfQLCtHB5hPuDcrm1jd/mAJMmG26BtooI
lOU+XfCIgeCR8LBSNp+VHqzJfD8my/7fY2rAiuXJVD2iR8/khWunGj4/CTzP0srzm6cRQCHk9k6+
PDc8IpJai7I2rwR6qHd4V3AXrm7sEu2AxitwWf1LwfbTq5agIfbjpam7hf8YGaLJaylVdpRm280t
JsZmII6A9v3xhBrcwWJ2o6NwU06goI/+IrvQWldIrIgs/WnPaq8Gif6Ur9nVl8bNazEsMC8v9VyC
wm/kQVYcc8fteVU41pdNfE8vkHwhLoWqWzQVac/a+Hx+Qg1Mc3p3X9BfzLs9wZlWEaVATGVguI22
yVaIiKr88cblUwNBbqYjUBkYyfZRmfTgtykoOU+SIumT8CQFns2G/SRUiVKxgEOKkwYJKhLzanWl
O+rFH02UuavzmSCkQZWSPXECHWYmyuP/I4jtmlMAD8F0CRCHNi9HrQYAN+kzUioy0Drbdhw7OZfH
mJMWoXZGC81+Rm7GIMlKK294R7OFQ3v1wT+NPT0dLtt5N3BMca27vOeo62HJ9wOf8ADR0zZZMiu0
6A/JDPmKOH2XdBxzh/eC/W/shkDuV+8WkhQbCqe2xR1aJy08hwGqlpSMM96geZz7/8xWtxYjLADn
WQ6mHXX858ARTpYEZDCAgWryAhx5pAtZgc6joDsdfZAqBCtLT+Kzoytvx5X38mOftTLOu0qR9Fy/
uKEHHJOBMYTZGTLwQqww99GuDget4R9wv9NDpvln82+MvM61rUMqdGi2CbLfTHCe5O9CjIE6oWRg
LZXNCVhnIWYRomkCHD1LZHnhsrRu7bM1A3nXilMhUa+sUoZwblVqOhF5KrxoPXAauOe9JvPAZ0Ee
rfOSt5AZnHa85iZXEzim/3CNziidQkB2DR0xw3lBm0+5R+U2Qbikch75yWmFdbmrkufp4sDPlFwd
Miz6/RRsdQzBfaUPB/gxtly+k1QYOz3R8T7mMSOzO2P2x45zeKwR1rR0aUPZseIEXMEcuUfZW/zV
a1/Esayz5u2KnPMu3E9MvP7gyep+c3tntkQ3qZxV9YDUgZ6nuvETXz5OYqxjdJeov5rGXwosbkro
geaUGxeav2ee6yp9x95v5Ws59Q/axLoG+MXoVQecc1/qg76cjW/lN1Ehg1IrMUHQqWd5rKp9UB52
Yc/SIZmXYwvqtZjg2gEoCTzZOfEHRQzRwAJ6SzlzFgveUAO3NnmBXfGBR+r9clCSKy4g78s4voPF
v19B/JOByRkbB/gPt2Xnxt8w6m+dQQPM+gEwsEQ+6O0ATnm1MAGB20I5Vqld94aKjMuMCDgwirqo
uiwzBx1BtO/yM4SSu1uUltQtcxjYnBcVS95r8ZbcUSz4LRZdyPSWJnCiNbXLdDKVGSGEdGoVASJh
5btrx/u7kDDJZtu2TRoHdlvXudy8s0EDEmW/b2ymUFO5vvSBIDT/o6atL10SsK8kv+83oibIOpH8
kSOqNEsHR8snMc5TD3GG87EHllAVmxuJbX3TzuNpeKidEXMRhssVL39TTRFY2VGmdYXnEGfU1KVL
Ah0xqsiIx73aNxWfCV6EAGtkjMKEMJJacE/DgMf+y6VtGN/5SbAtxscYauKbx5EyekClo3vug/TM
y1PfUT5F8Bt6WFj/Ofo822bns7ZB8e5kQBryhY+tKtqsY3jZUMEHZw0RzMA6N4ZrijBPkFE/EDix
rK+p1wIIMwn3PBbACh5qvMOQINyo01Tnklb5K39fnW9JkOjM3kS+gGr//guqyaWRSFn/RAUPsBPF
VUhfyF/yV5vKp0Tohe2evJOYY26nMLhdgzMAHvrIFh//cjOq6zupRe66wPD4g3Hw3yl1ajUV+/3/
wUaCOqb2V4RBTWShFNPScSRWoAgTzMpkTm9B3kWtnnrNq0m0lFx+6tTjNSicwMoG8yNppgMpIpVu
aGmdqMkX8J7984u5/ScgjJ/l4KInw6nxd35v4kDyunSB5zHa7WYO+UZu9WwgKE/tLag3LhuzBGEi
83LRM1T552OK+Mw6HyYTpkx2BU0+pbiseWZ9jDEW8uPAKx5JdVVVKuBM1sXIm2lddIcO/j2Wvh4A
LeqMWHK1Z/+d3v80ZAWo2aFHrEYxBss6JpW5OeM1prhtnELdzC3JSBcaCn1KjEn3Iy5FxTT+BbEK
ihLmarn+35H47j/Wno57X07kglTbhNKNjuV/hBcPLWHXvgLMNqL/nHQJW2XtW+DCsxQY7Xsn2/rn
H+lrX3d8BvNgj8TNxWqBb4EAAbb08qXnEMO6BDvvT0CDw4hUjIUq17R7e9+TmzbFdWc4k/iRPhUH
APqgWItsZpE+BWoVfsKZRtBtQjRlH9HH2nS0CuD9QACmM+isq5ChwpSt2NpK05nc7RNE9KUOm8JB
nyz3a+yaMrgbK7CuIsbQMrae8qD/l6QHTiOWZba+KrpiD5az2C41IDHLlvIVeydLvy902MMdL4qD
WaBIKJowjSK6tFTNj+7wAV1w4n5ePlYvtnE9cqJfnncaMDgM4iMgQOTN8sHPnlr7u1dGsNP/468B
UTVtT2tkDU4omu2dKaM3NSoQo2V8+2pX329VReOK/2lc+Za4qr2EB+MR7tI6bPzvzsAAgOiA86hG
n2WN8Jgzgr0d6BU3a5aNATnI39+WnjUCU0EjUaZjMxHiAGRmY8h5AeTWs+ZHW1nSrELyRd0EI5Wg
QTQp1+EycmsX+fVBfxqAConPQjRazOQLiRWKN+Ss0xPLrh2PcqvOuvfp53Lf/afHpBX+ocAL5yDW
tG9au8jLQtmsl6GPhaY1Y5RrT9e8WLYtsulMuskri/edRyUGLHaW4Z9bJHEwjBJw4lDWM/3yj5UM
WUe7Djl7JJL5ajql4rwE5MBcM7gku3NhgwvGAljWUsiJR+wpgFcYmGxrNW0V/KKVbVkMypucNBVu
cEkBj9/FiwsZJEw1I3rXeLvLX0cOf0nWPrmUIoJnr6m2XxpCUQ6YyS+jTIPMeiF57JHpH2ksTiyA
oNgwAiMWq/E6k5hBjNHsfPAP/LB6lJLjjy0MceMp5bboC8fktrAEFswJruQ/aOBni3ToUaeaR+vr
szxR0zDXzqiugioVbYExFIkG8iOz+6JMvMA3FLlWGRGiFwNox6tX3H7w4u7pnPTphRwsexzsrh8a
2EP0yzeMfMGYj2RFRFcScNLKW2Z4B3rrLqkBPw+Nlu6A6KSyetR3fdlkTwT4WkitIUPkgvx0olOP
xnKWLLd+mMq/GT/Re+VE1xTblFhd/mXjk1lD/RiJDqrvdZ0rhvp7pRDjCoiqkP/NVdK/FgIftMOL
i6esrFMlVMseueo37rfK7Gv4grizANW/pSFd8LIFfiin/NqwIYpJJPHYlGBFtVCD6ngKIGXVycfx
3efu9c28x80Hk1gYL0UUWuDjnRkukg4g0DpWbYMvxyPZSZAwtY+MVE4BswI9L+Ckrj+IFqLgoNOL
Lc/SoQSwAY+vEp4H95qH24zddoPc5c8rWFQD6t0BLI1BTnrH2E6d8gQk7qo6QfoiWH8hTxk4XV2x
skhIt6/EsWO72uDDXJ+n4j0FKOQeDmbW375jro/9n6V9N84MlBszDWCBA4e4rUgPbwInmtVgfgwW
8RKWHjEB1+G+JgFy9ZQO3h36r8I2XRNS4A2kwPYgMJT9nbd40ze5knEtsV0dyqaLE493E5s95tzg
fQL+zyD3PqYCVHQxknpnCRNalWPM2HNWODH2f6rB2o33isiVgXG0/gS+0OiL1p94OKSvbIkEXJQ9
BiyM36+34+eCCp8XiZx5kkNB/fPMJ9NFXEPKUtM8pKaINjar8BYb6zvFwA+WGnFH8fQyHZFmi0VM
OhK5wnOaY2VxLZpFOAw4jdlqHmbcRI65FyUdLlGT8/1y3K/xSOX0T1LksoiNJxPyfmspqlTmU7mJ
6l68RK/B8WVqWnK27av+fkPCmXaiC5G5HCeZWkoCc/F4n7xs9avnlVe/f/3jRHp6OFFkfZ928Oi+
26G6kmvB4b3JtouzMF0M4fkbmrdegxBOl94vjMg79cTOKf2jWmZ3JkTz8JtR4TgEd4w8Ae3csvL4
6IGc+i3NC72W+bAq8jexwvboK4wiFIH/P0j79XjIsRkLcfJE59MeCTM0HAaRgBMQKKnerxLShEGJ
PZQnXtRkVgV+9w2MhqBTWAYKY3/dRDKb4mmYXKYgqMDHuvAm9w8gOFw8/EsDBo9GBLVFk+Uhxcd6
OBfq7pbRrQ/khHKWx7IvhDUc7MyVPobCwkqlk9s5J9W5qbOaigUU6DBlE9F2NTdtPgdaYfmfKt1m
TLjlDAAsDJ31BSg03XDcvFPAMpYMYL9bXIoXKoK+qsCmfa/jYJUPwiGhvFFN93Ke1VV9mtsqGZGO
ah+s5UAauV6olHP3J/myKC+MJxmLrqdx5wLBJ8pAmBjab4k1NvPyFomusEpN6QxVeKPoDbzetY+e
rf5H7Aw38PjX533p5Cu2My5FhmhcFDilLFwQ1W+uTjlCXWMlxox4IADeSEfiDRcovImscQEZ/tmI
FsBEvhu82VyLfKxFetpCsA388qfEooCbFB07/zgYS644wPhHfNrCqNeo8j4r/ewBCG+TlhmsagAF
EZapM5IVK/kLu/SJW8G556h0q92dLEneQEIdxVD7HeMRvL7daQUWdWacvScjnyLGuAnaR/QWPikJ
6u219tJ3clJJALcCbiijVd5Xptpn+QJeYFiGsHeyWpdDk8RU0CxrOBrdDN3PlEqQPUc+NYhc1oUg
FAb8uD8nnbcaV5SVXP3fNsLdG+dGlfzM014sLC65C9VikeX4lKJo1com+bNVUHn57ckb3UDVjevP
iKOwGeJkyVuv8neJDyo3GUk5bBqNFB0mDKcFRIN7bwnOnTF4wWoI6KFh0GZGJlM+iAXZGxk/JHK6
bGvb3bNhLV6LL1UiOa42KuChKJWrYz72CpOTat+5u4RilNPb4gnFL9I4f8Fr+6Q9UYTN0nuY7CCX
q+VTaM4U6DNWQY959OmASgQeRluPWOQpunUylS6K7x0zNeJlqjfYtldo9R/bklPqrCfOkzlySPV9
0CjzsbbiIhP07KoyFVq53UkT5Lcmjb3uxKOOFUrkh2fzoPvXi4tMlVN9gGScWhWwTl0aMHQ2Rsp8
EJOgEPSbub7Lq/QnH4INfWrv0lfUBWVuFMdwLNYFootEXwLvitxdRNxzh84X9CxwRvrKR+U5tM+L
37JfTHxv2zGOxsuPfkxYs0dWpZgE9iNMgBQOci111gFLzpCPkV4wggFDLUoTXvXyCN9Hv6hYEZlr
vLvyeLRPUWjg4EJbwHENwuO2xH41Zrd7SMmP3FKXZDUmFwc5dQ1yredmf63+LgR9+WebiUOLgh4d
Y4w81uFhQM6bfkGVZXCQrylOWZFg8/rgEZ6OjkrOhnvZTg1ihbwmtRidOJlvyj7yOvsWDO1643vv
r0qUaZeqCc7pe8BfuPV4WhMiSQaWiR/RJlIyJABavvx6Q4yHglPVNus3rIFKr0trrPkGg3PAWYQy
KiVOvqkJesQJ69uXXfJfJBwLeOmtRZsCLahf9otdnhpG7RNpz9BTiN6kDgtUmhZ/nTDpr+pNhBeQ
hZfitl6d2++4cgdzJl4QtDethVOZ9OYEqlnf+q25rDMwT8FfzsoVTxf1hxozDzSPsWycMZgwjgO2
tZOfQIrNSHCdwb+h2zqqmTFfisVZFEXuZakuvw/4DaegFvBwtVPlYjxHbk9CrlSX2ZxA2d1nZqHO
GWNI8st7q/xHzbswVjLLLr7yDKxaEIGUvlq3sLSq4u6Aqa3wCXH78gZqtMFQAIo34ebcJYo0tdu5
uSdwMuwFRdNf1NvgMp8Ukwfbj3EmbY3HcvGFwGEx+8GjvhRUXwxEf1sCZn/YzmOQhDu9UPdSU92A
Gw32f0RCe8bqDtxbcD6zHOGxf7MVc818FUqigEi7Eb0iuxV7uUTXSuGA/dlSaXRFiqrQDAeNOywf
s+pCFXVb5g/Id33B0gl7lHdK79wglZr7DB0dGXGlT1DXtNbgSsofHnmo/ObxgHTonM7s63d5VeaG
8cMJZvvDOck8OEIa1zJ5KR0qrqL0B3APqWnVqelZ+kzTms7KfcCstETzvHofw771d+DmuQuy060i
GKuR+c033gahe61LutA2N8SJo/EO9mE1Feh4TGPAv2/OqdQdbQpoN3K0cRsFx49/LBBwn1DbI9BP
iWwnUfLQSTC9bsGGwl5HWm9YmtX+PhtRaPk4O52TcI2XE8auMUABqoho09UYtuq7xKpMcpXOgWXz
uaVLD43wUnK+UiRX9vKxs6r2HBvot8ZT9yWeykctUX8Kbh1xbXkXhUYbAHe4JRBLRNE6ZdbZW5dn
cD1sZVtlVT53odkgqD91hptrzgqTTlno8NVL7cHCfZWDPQyUJaKAxW36jcR+Iao9wDraZj3+YlHN
jbjdUsUVUnn3yfZRi2YtnTdnaE9tmO4XojA3I/+k38Pgi7xhWdAtBChyr0zHdd3aiYwef69N9mvL
oSgFiIvPNU1AJyG/1w4K08cUIqFtk/I5y0OV6VPtOCAIBVOPZz+62t2u3/g55AZsWFlcZcyMzQLD
XfTK6yoFIkRlx9boolHcEi0T/zll6XoSmaIbGqA1DSEpSvAToh743QyLzvrQCZgd8g60QEhTd38h
xb6V4ZW12XSCgE0553ZjJepiIf4DR5jI//Pm58LIHBqCeR1xf0DoniaVaPYluqkxD0wcvBMp0yd7
1SApwOx0WV7RUj1if2i1+pW7WAV/zkLmXUnHL9xL8hpPrR4H5O77hkzbaWUKzjKkQJYD03wMJtxS
XPQQwGy06sCEM+MIWWRObo9wu48LkHtI4uBblrt+xJ1rLx6NebWrgpgXq8jv9JKcrwdCztn8bo+/
LJV4yY+bMO/UweBZFZERt+MC6EhM5kjr1BKdQwGQvwYh4O2XR+ehQkPV34aAs3/8aDa03dUIGTAH
NE335LdOPRBmYaekNbIO7NpMffh/RzvgTLL+K2BbsK8TyRDDXC2qiijoHaOFq3vJMcY4wWgVYpXa
dXKnC/s7zbZVgIqGfaqFb2fc++ZFImDr/fm7PjSmaWJPp/58G89g08jgF4wSqZiH0fU9yEmRgQ5G
ohZ1rV41FQ/ySZk5sCLSFLXh8BL8Smw3iDFTIxElhrlyapiB4bNGS4XsKu/mfqng6E/603B8QR7f
illcOqg59MzUDQH31zsWAqgDIkW0L1d3A6pm0lyEwEzoUQ5YJgfnHmdoYgcoDw267tmxKcc3xdl6
oF6XPRQiNdbQQj4SIfAVpLYXgwxSb1XKrWcVg67KTlJukbunx7kjx0NH25hqtvBOSNJWcwtxow8A
PHPrZQlYwM+CPVwnYDxQzqp6vcCAvD6frh5XSvWqjexwW4XK5624v+zA63dwR6LhVdwzKDT4PAMO
+JSti13IkzEJmUHVV7UDLJ89uI5pASQLGThDJO7ii1K0dU55Vzh0AKpqru2Zowb2IYUWT45r2VRu
n7sExR/PHGRU0pAnthmO8eZhKuONX/MVz1MuodorZoYEryx04v+vxPLKh7JrLlF/pp2NkaTHHyE1
eIL6vh+9K5QrXFbBrD0aw6djIH1Ct4O+fxqvT/wzcoMeiLff01lgzpFG9xLOq+ZjCyo26MYkjLnL
EIH8bM6Rinf3ad36s+EqBwC9mYAs1jP0qmaCsP3N5I0o9gKXVxR7fUAMo/eOq5b2j6yx9T7LX1dl
tNpvToweyMh1kupgoQ5LW4MQe/iTHUT3xEi8vbBjSklci37ng8Lz6DDUz+D9r/Z6uxpoogP4OMfi
wwiCSteBctd9ONnTOF9sN2ygIIHjxPQ/pA8j1lMRsZX+Z5bkIjV5qji2g4+OkJJqIdX7h/Qw80xH
OBudc1kp+USnvg29U7Zf2tz7Yr5Ik8v9CH4YUdqBBjEfAg4muaPmc1PDE/0LmEY2FItKx0XTHQST
A58FDeUl8UAqhgkICXzrEXBw1q9ix7cuIWsP62XvLbknvnUo7M//12NVxazxbWAvx5vvtTLnXLaV
R3Jnsf3OLZ1C82bDZ3tQMh6mRp9JGHL3yKaMxacjeN8MPJxSe7fLW74m51IIjleHfa2R1G2a7eQ6
4ldrHyUglzG0LEx5lF0lB8H1ObcFBWK9RCKln4MrwbXAVaLpQC/ReduPhvXivc/H67kvfzvvWfLF
S2CnLgWga/Mafw1mMnc9S1ULJBLOKwjQm1h8uQWpE4Sqov/cUhVCeptYPNkNFtwWVOB57cgONtaI
Ewd7EmOmuLrKEW2Sp3bP7PXlqrtH/2lWsrCz1XeZdC0fYPSxTNu2GM3g6ClV1ezjnVfqit+CvGBw
+suk6GmDnA7X12J8aCIciYsf4N0YwmbGjc3n4cjE+u4sdXpm5eH5izYbyhn7zlgUGtZSwZPfcgqu
juZRRJ0XFZn+372snRTR+hVJcZzXl/ymcVW+2FRYfUEAw+onjqNu6aam4Cgbk3BIwz4IKDObMNZy
RDD/XG0XJJTUltbalO0FqqYwulV4aFhuxNrqna71IouVhQ4rQUOJamCMN3yGEbvcEaab5IKJZDmm
LltGq9AaYVsOqyZY2z59xjrd2hzfJ7yt+kKq0A3MD9htLKF1CrSZhEYC54OwKYaRMPrOxPSrf4NS
D1Vrh0Ov1NaUj1RHqjJ3pneX9xKjNJj7H/rbroArbdsg3wWxLRQeGmtD28sxKrJnhROEVa4IFJrg
ppKppNxqRvEuJVp/+gqvyF+VMorjHSf4wDQY3CWgngS24DMPEAIQDWEGB3fsc66kF7rdClh51uWG
raJctxD64PIaXe/MwU2Gw0FZRGl/o5Oc3DZz+YU1EINTwpVqt9UOGnB0QAXVap+XYa10i/z0qQ+8
H+Mk8qGzumeCTHhm/AV2FD0Q4Hwv6N1Y1ENv0UZyRGLgX49ccgmHiyrgXw98dPd3TDxSu6pb/QTP
15NXK5b/VPLwOAR3GBYsP4MK12cSgQiQkcqRoJ904IY0JfR5A6JMROke/rPEisAtHYjLjLxHA2Sj
OtvgRcw5hBgkImdO0y7g0yGa3KUZ8XQ99+9qhLO7/Oi0T047l4fz9vhfvYL014Yg/qbj3lHOWQoW
c3VTc0iAeHX5OYy+MVGFjctbtvCqn9r8Hd02tiyYe+iDeVSKz5t/+XpCm1oweBXE155rN5yRvuz+
TvkvClw2XfChH+kxC/wSwN9HAJVXTyEXz8dKNQRxP2xnCyr2CpGSq+xtg9q1SWXzvN2SnrsNiokk
HGmUCcQNRkrqe4Ue+GrXIjN08bV41JSS+hV42lQ5VkpegeIJaP8XqOcHi9lIU12paMQ3auy++aJu
164VK6QgclxHKj8KTzDoolriH6wHzWF0/SNlcunyLq/sVinHbdqV7Ka2aw2hWasL5BAWo0M/5cMb
cNXwmF6IhZx9PIAgjXcS/CLmBgx09bubVXJapVcVri0Cyc40z+rA6xI1uqTnlHPvrgWUkP2rEupU
WvNWADjA4f5LthoNnh5fi3sEOlZIEayiaX0gUIc6ooT8P6OrsRbR2+XbJXA8wfJ/DMIoqUMZED/V
wNZ+jQjoBa0NSBDquq2OLVZhtv4WR5D3n7b3aVO4UBtF52nDLWb6+1C43IJg/DpC0bxLGNsugXWP
fuHZ+bmLoP+SR/Ad1WLEpwZJIej1QqMM1HitUkGAWabkCi6jDBO7NuVITLvJvNLziClMZdIhbftL
NC/k+eR14UBsr9nO1NpJp4N2JBMTyI1ewSp3iACRMUaO5eLmo65KVfjG/HV+ue4tpcZ+demMURBj
OXzMEWIuR2/nchGNJqxHRbnxGqftlSQznUSwVT8vbH31W0TzcvnoVB+TdFzHHkv7VEYt1xaK+PnL
QQ/g9ru7I9Y1nkOJU/Q2b2n4osoaFicprJ/2PTFUC3u/VgghMsOQtVastMSQaA7EbnLouf8FP6O+
GtH4WKtb8uxhAeF0Up4sPACCKmtS/qyZKicUMwBy4QmaZAFu3PL8mNcR0QF3bitcrBMGoab+iZFx
QHS9YWdg7kHkWjp/9lw+yDPDqUArxQ3unX0btP5jMMjh/7ke4dyguQPJI5CllZIwc+hGeQFymM7e
Q6DlmasuKjzCIxbGt+LmNrvj4XClOyM8KHZq91/nM8OgarGJnE6781JW7A8jxvQXdpSIxQCU2re4
VmDo9UVeYamcCVitw7GqojUmn55oXkxLqpJX2AnGuLLb1/867b7jGV7Xf5uQA2Hn2hAzIDUMeHuq
JN7z+rLcxdR3w/mHec0nbautm3gfjbrsWVCOoyNeafaqaWY6tu/iQGVgKmJqSqutWzQj5WZy3MaY
5ZgpI49FRjCT/sBznoHNM8Gjiuk7ApIoOduuCZFAufWqHsWp9UJleAGPS6t9sWPtZP9P0yy8jxDB
o/JvbsJmKDcnYpixAx6dp2XOvnacltJsLSQjrgu45BwQPHB1nAeIu4y5AteqmaaZQPzN/O3mCh2c
f3tF1vfwhfpNigRv5o8bN065etxoUeuPXZ96WUqe+fpcCEgMpfcEP1nDQ6Pb+9TDgHLRdGihJDQy
FcWBmJU5SCNXw0swv1x94iYJI6Kf4KFtGgEfEYwzi6A2cnWxJUDJwkcXKCQBKzYGL4EyrHizA8bR
27o6okeVYZm8Y+hrt6xn9G/O5TEgXhuDtUUbD60thWA90653mm849FZP/r4RbkhqcXVCoVC8uxI3
WesZxf/oJQp5PSA2TRRu2qpCZrPjadAe03NUcUKXvFB3FpbWrNdnkHDBaFIrb7mg9SMEYLfUw+Ps
HTqjy0WM8KNlLn9eZ0pFUQmibZpBGrsE2j6ssoJMR4e2dB6V1eDqLFXvIx38IkH6xVw2fXs8d/Zz
JWq2cW18zZKNodHI1tR2fNcfZX6M6O6mNaQDoV0/ocEAVID3PiPnbn6OfnmZqVTZKZ3WYi+xL+5i
m0qPnp0KwjSZ4n/qpfJbqsXvi9YQvIbwhHGnwqFsVoKGP5kKm1vXhNZvfiB0p6fO3juXO9JGI2F1
CdMfMNAeRsU5wGxyG2Opor5yqLGqbatytuYIfCfDRGCsQQbniW3/Eh+QNlhOJq4OUEh5Q08FwvqA
1xepqn4bbisuZBysZs+fBDGlxMmwnyC0rwKngln7JC0QWSHV9D9E6bsRhBlGAqTE1uetCsRGS2Yy
dLcEDyMMF154EN80zj8STxjYAsr/6k3u5hEihw2u+rgmWweZBK4f3Wwq1uEho10HWQ8QE7aNPVzT
4DIifHShLN/YM0tGZRGNxmsZOHH7/bua9NSKaYj4l3a4YP/OQlc9NqVvXq0p8r/vPb6wJZrp5VNs
y26ymjd14piizwVxSyEbZkgMqvG4Xm9+FDIHyDqtT9H+XHx7kFQ/2U36f7RSdjKrtNerx14tVXsQ
geP+XkMymH2vRWOofPkPiCB99/jiD8+dOoNzwOKQJSNhTN7YuTQ+D5OPTN1o8khYgxy4u8eGvH5w
AYgGk0OVP1JQSyM14ihvwPs2HsAhcB+80+y4QEQE+44GD5VsU/UkLfp4hbjdxDNE5BiD9ZEKb//h
g2U+4h5e007mUtz4mkGsN03hdcUkFy7qOOdtVGUqxwdG8TsbnZa5sQ9TXeliGxwquZ9ksQM/45QV
mZrWyRkpoTDbVz2JmmLfQt4DQbY74ovjl0brSYRV37eDpC98if6K71qM7q5xwQVZEUBD7YIn8PeR
1QG4kC5idnQSw9UTqbKln9QRLB3CBMVLI5SHfXPn/DtTC0IVNFgyUaJgcWOIPglhElr3Qf3SPRrW
/DyEx/ZdXAIR1xHGXeIuvTyCd0ZS7iL40PmsQ38FVvaxTVxYeVjAte8dOXC36OmrJWbA+JPkwwLE
JWWcWfkq5Xv3kycWMXoiIM0PesItvTP4Zf50aQzJiFaEdgVLDC172OjhGB/zugyPXw9yQzUdQKky
eth6srhJilqpdg1fvpvJm5tkCFjcne5AdVR2y8B+/FqsV2LHpweZMJ2xSytSvwKwUPyW6d4sTLro
j4enQ+sgmp9T446rKsP6cn91346Pvl/Fpz0kAveXOyu3iCiknss2rMFW/IX3AoUGPIDzDG1fUlxR
d9FQiJ0nP+zk05UqbkJtKqN9n6dRNIoke68Cml8HeBP5j9+r7P+mT4RqTMnp/OmWPXwq3huCFsQi
ZFpjbW8jPBzzhZET9XOKAIgAZlUTLB4bGoQ9TbOmpVu34rc6sWb22xBRwjX6qv8xdmQ5bvqxtw32
FBP4J+5J+OeGPSipUAiAnGxL2agioapWGkw3OiZRn6U71dxeaRCLZPzH+qclUpwhgfX9+XSPGhgN
N4rvXtOGXba8wAwgBtDQ4bVIKjcbZ/Tgh3r6qEW8nZq17hHKD/R3LDfcnB0NxwgfKCSgve5kZMMn
mC4OcyOh4MoWz83uY5uiDTDNaR6E2TS2jZVKxo7HNX/8EdUElXvMLMNskA6mGuaRucoCD7FA988S
UnbJoYirwuqvTADr8ryz8PrxjqzFtDiwuvea+tlujNcHOvr01/5mhwJlopQEB9dwSRrKFqelgHpb
WqQkbTJY7YSCGJHC8jrqKlBWHNyANdCbnw3M9wsY94Vrlk6ZnQQA/r+xK2TiAzXmJuue5pZKlQ8w
WrvlE9RQlrf41ab1di+Gj1ukCpDG/U7I6Kek6rSEF4hjOl5bm3a1AA4LuvqZ5Z23udJEsyVUslX0
/BbvYiORp41qaPz0L/ArXzjUksiCuB7J599Xk6Jc4Jh7MTDSohnax5ZW2KaQYZmdiMYOe1F+vdaq
aGBazRpLiWCzIb/T3ovD7oo8nWK/luiO8Saec27E39FA6DdHwUSPHGB0PTFkfWib+LgAgYh5s4ki
uQOS97CJc1Z2O5cOvl1TK3o6rqCJF5ZIs0yr7OF0XqATQ/Og8JsrjAdbIUKXN+3ewfX5pg1jZMHt
1vUYDzpEmRJCDQs/MZX9MgUCsbxDtwOVx8p+g0mZ0SVHnXtkcadbA5SCq2hKdPjtmmIabagsh9k4
WRCiCHCmoPEVvlVzoMq9JiCL6tzuZJczwqyLtVh0RBNC1SteDqDZ1GSJ+8dccGDQm79cuLdtYmvC
kkjYLj2Yr6cMSxKdDwYHJ+tKutnRFrgtwP8t3iHVFqxJ3cWUvCBX8OC2NahohCqHtM/I/5R+ilhs
de/R4QqqGHbTzGdzcLGRVHlkhHtbkBBsN1MmDALgeVvl2SO1qFHJ+TJm6X0iGjMka4sbr9txclxP
aCIBoszJ2JDDmTLEAlSkNBAftuGdJ8jXXRtHCnMYyFr8xn6s1vEADYUKXw/x7r0zeq0U6KVjOqi2
xq98BMEAJvRMw+/baXX+nfkBlzYQxELF/ok0881aUftzY1rjOneRbonhvsQZotIm1aOJeWUzYDuJ
pSXdzD6cZOcU+/DekHuLySPsX2PBcXHbrBNXLd1rQPMRUHW9sReWYOjNm69Fu/j0MIHLuakzmclK
zRbzUp+CmscIT1wLrU5tJM9AcqVRvabHYAabno1j+IGxIR09Akltb9SCi8HP17KFeYtPyMLzsivz
2Nv/LXhrAujsmDdsoy7oJO5P3BRf7duadEw6wgpceNdZ1beFPmj3u18SPqsCZOkaZ2QcarORrCXe
CJWsPnNPmhv3kmsNLjUHUQBus5OyaiOx6uXDj2P6O7KFEWh98FlQgFTz9HHfzRSvLrbbOWsjsk+/
vyLV9jhM/DGa5VkNsNZiBRrET/JsDkENXuTCBAa5Uc9i68Cm6WS+ood49Gsq28y0LZHcDf1xW1Je
O/Gl1GTDKyEVrAOA2XTktNG0LffjkMmNOj4FyECwVK+RA6dt4R9t5CnIwNZ87YK1ctujJ8alvtjV
krKGf11AdK1WnvOckqDyuW+kOBJZWTQlQRCwz89nHzrXUEk6CjU3RtHFYEmCFRorUfs20X3wVIjF
7LRllDbQIyh4MlqEnwwl9zu9ziqXY5yo62ZzR98t7KojvQrd0UbimkwoC9DoFXjbaYJnLpweNrwk
Yrrp8sYueeBphv0R8BCNrC6VgX91b3+boalYluR0q6jLfYyew9zLxybokrzO4AYdYtGXi6g8lnbY
w8NXP13fM7yyuCAQUWm5Yt+rFBk//8VYoO276FttDkSo+C/kTXlibpnAz0sKB9DNm7O/5PKi9w3T
I6scjnTcrlpzCxFuMuLy+6WLYc0wNeUUGzkB+p9aCUyjcu33811oGklueILGw/c8Z9l+AkkXfBZC
5pY5UU73UbsL7MuyiJZEGIz8VaAh26xtdHYo6PpzPpApWmMnZotcV0NIh8VX5iZ4VQdiLqPW95Im
N5wdrNZU0yeTy9VUlEX4hW+HyKozwIsy9bmi44PXHgiWg0Upq0rSbKaMB6oGVr0HV4jA/boRXQ9j
CLfD0qiTvvQEqm6FHBh0Fc9V2W4IDZ61P4DpA5dgyGdOc3/fF/HfBgH/DSAHOruYTAXYES0XGSGz
b37JH46qFHHa2f1uCRtD2XVpV5UUGtrOo5FGT4p5DBpvojHgelUvdsYrsNNTWo4SpQiK/HUbhhN3
um1l7R01pmp3HUryHdpQ+moru/tmz/xeZss/bqKe6vm4hE3u08AifSfncMsW8nFiubRQWMT5ruEU
zKBRuMAx4pH1prj60EWMaEuc021oH8KUp4ecDrXOjQ5iYH80d8HuxYAuyFQIiEyRUHRcEzyEQcmK
1DUwzB51F2sHF1sOz0EygDVQ92lU4RaYNFG+P9DFX9WZTb2HkvbVb1mDfHvH6qHsWoThG59HCCvH
QmP3yPyD2COOWwHBhxjhDYU4Egze1sVJ0pSZuJVOjnGPfHxt/fqeE1tXUELbwHiEnT+QIjrYAZ/1
yLRic4P2qzrCxY9L1z9PnVMGsIP/W0MdDv8cRz8nVVARB2mQibUeU2qCXR58W/qU7I1my2qqPfNf
JKTBCbWbe48gOKOqhXILq+vQkzu+miXgcTwawUGxFPDVXvQpYq5z2ampX4iw6/D66blhoBvRpkLL
0VMe9vsisr6ZCuxzJFI/J5xhguu/EOAdcyEZSyXYrhyonyuS1mIhpsklUjJh/6c2leHYT/nSfcDu
ifXPyRdawrjF+xGSwqAPzq1vpt/qhoyCB18sYcpl/RNtU08UjYZErxWdCdZo9hvVWp7G5fy7Dk9b
ilCVgbw0fURZfCTw5Csq4YursL+tirRMg3PCX3dUhFbRhBRJELv2XMNF/P5OIlT0l2Zp42YCzKFd
V6JPmmK15xUbQn4BBzFV3p2CG6qwmpZwrlIJsIzDNtIaQy/pOE7sPsAp3sTtYyPryAFyPQZZzdEE
fG1/wMSk6ZxL2+mJUXumq6bsCACRZ+pfUWciQQeeYDvHR/hIlRDWCO6zCZG+O756cJIaHLdykupu
ik4EZz8oJQJzHrBoEgFeh2UQxpPA+VCKHuC1GquWr3OtgDDHM9rLOoJqJXBetZkpd88RPd6A+gMA
ITrsz6RJamgi6aepwWjnSqi5Xwwo65+L5dbSP7hWmSdzMbW1pfP9uYvdTdzfPWNStUVdKMYGeduV
tNwS7llDFIgW57+y+XOiYDlfuC+NP0SiaPXD81tStl5dhYCN0ICjgDbM5Hm0+c8yrAu/0QWRKW0j
sctfmR1XKWcxxoe/0ADroxtQf8YZjqGM2a15Jcb7J3zAVw5B6ZEEc5p5GU6QCH38bwQQUC+iuJd9
zf9zEp2D9F8TC6AhPSAeaBfSa2p7KVrF9Vb1BPAJatkNy+TwwHZJWHL6ZX4ZjrLcKbgRz8HH1PT5
HgE18Mv7Tq99UrqFWsbrDpeb6xYpsx2u98GeHZwm8J1J5U0Wcw5b8JLSNwsj71aniM7FoZMx9bUQ
1O3DE3KPl+OwIjNga4JIotToALipldi3LS2AzZ+xQIN7/YMyqL3BX24l8+3uN/KVV64aZIkaX1Jr
BCq9Yy6eUM1nqXebp2uPvfqhQz5IKeN94ohLJsCTXg5awtFTiY6JGFp+8qmSBh+ZaQDo2fDr6NN6
TOey+anM5YF0a9wmkeZL7/G9eNzcMPrCZX0Tat6JSPJB/+wvcmYyMLhe1A1/p0N3NoASkx1rd/lh
PVJ9QraHhN3lczlBVbI1p+Hq5wotgTAXhuqJlXQ9yOaHGoXhPk8cNTIw0VfIca4qMAAf/liZ8ZjY
lEQC3LNuFBTkzw3BcNeJZI0vaYkWv5eBp72acZ+NIKgkjglgBrHqe7CXOEhAQl8tvrXqHQzsY6tx
Eu92c3oS0x4XCTWXzRLVie9ED0KSY8ZJ8R6qGf6F2p/A0Ci9/JZYYvjhKQOPbntHoMt4Eqg7ZaAv
EX8PCaZWgYTNTUUgb4r6tOH+NodIDkc8fe8mT8fhmaZ1rWWunUb3ipSZo2Xyc7NIyziHf1O0C/ul
yTfVuEEnO7V0xIrKfEPCGtRRGg6bXTBoni3BO5R/WjBrCBz68zrmp6Usyww7yLoGtMNwS17IrMdg
k732pWpuE5BpAYGHV7j6PM6kuCLLmC2jvCgGGizJAK9//7uMWg4sTCnHCHbD/Q9eXvYqWtPaMKCh
a2tNXk2Up0Om1PZJgFwSE+RsuvojLXOdtBbtbtDNh3CVEeNPiHcMTDwWbaCDq76c7aRr5rXG/PDc
9Ss1AJBZu0PFCZ8ljUxaoA1A4Y7nynnWUt6APQUlPIe57p4PBcKKNXm2vj+owvIiawA6f25WFk5G
H4jPmS+H999xxEM1XVoJdm6hgn1jy/iSkJyKfpQhcQhmyZtMumX2E2QwCMRYRwONAHZHVdX03e8W
uP7W8qIIJXAVu5X5UAAULUfCyhomK8QgB7dbXL0f0hTQe4hRfdtCY733n6ZZ/u21PKInJ+mnQ/AZ
in7ctqPbo+b8HgjiYsCgIsjlHy2UBq6P3k5X3Rt6sDwH6hhTAgKWe1k4PTqW2UnLWAhym+JvPRBY
IkoFEkntzXSFNeBSh0GIsWbGEZ2rRhZ3i3OjzpmLNyZ1o0pQ93kDKhxK3wpfnsnkVC6eZlapmBtx
MO7/khAwUbHms1o4HZq0C0WmN4m6jfYaZOVmUbF/h3gt/kFTSh00qBXLZuEMr/8TyQcPWI64eZxl
7anp+GTIAiqgOy5Q38gaEYdfRgp+sgmVY5PuecG67xM3MgVd2psUz4bqa3D3rMQMgMdbqYbJ9HoL
/a5GNO/HqdbQgeh/edHBSkJm5x3Hhmr/GAAt4XkdYiAj4OLoHiDCMQQ1+EbQTuwNnClNIvOQUteS
tf7PQOBOQ/GB6yEKybvpowsBmFlO42vs5p2G0RyeeUsLjXNzKz5rm+psTeNSE9UWdCNUwF27QxVL
AIx4YGx69jZPyD1QbBRTBZBh08F+5MEgXNjV4VW310m7lRNr3wckqmE8irTYCpWMse4MpBkfyMxu
OtodflHq9+Z8mnNpm9vZtMTPsLmx4tgumhihjnuBp1C9FKyOEtygd98w0CdILEix4jSy89IPApdE
pr5WYfx2oq6a3qSBfeqjPjhpeFSnD6/7rQ70nvY0x1AJKjHQwdpWnktt5DxP+pjoP1GuI3I6T7GA
UcS1bBDkfM0pqoCDWQW960oWoj7F3Tb1V9L3F0fa6gbyU7NdLmtvmPRwGTQ7NQ3LFNnALD9veY7A
jHjT+r3ZgUUUkHsM2Fvh0IoTYdu6yvZ867yw1/yVr+hJpkbAT4mlUZ1Icu3Q5EMwVTyRY6lZkgAP
ddeuWAZJ600eRU4HOXDI+o9R/YTJN6cX+1+iwA6/e3XwRU1ycdjrVR0EF8P6+rgyFYxrYSlfOPh0
MAIva81iM2DwmHbSXjSpjwRWutz18YmD9s//6zdjjtTtHFXVpyPj+apZ6UGXaQ2l4tND46QMReEi
1MUrOZCFBRWjMkJ7ALLXZ1vfaq8rhvkSuVuJ3ZOoMF6S7yeWWujHQc7/VYwj0ctAkwfAfijQfGhm
FuXblVac3DISKUfPxWeZAXq/VyUpymCObYYq05d8vrmkacBw07WmESoiFg7xC705W+Ahkszs+fuL
buU9+ZoaS9jT5dJ6G584Hsy4MQYdwCIa5Dd+XzDBsuB+Pup97ZfiVwvagaaNLvtYu7fDxijSBxdf
mwoFXMuCZJfdMeqSzMB8Th3a5WavlKRSdoawBj8jp7mgr4E3u5LXl+Ov58LcNwtkKGrYPUiPRa7f
7IpUAwHkpwtU46/qNNWiMoINxDn3IpJYojgvOhK2WbxcOV5xHbYWIzFlxPxPeQBE0Ig05f3NZYoO
feiVeJvEHBWzuWuLSJsGDHB5hdt5FD+C1FEwHwW2UbmO/t5/On/Q+Qv/0rg5ACMGDgUGOBSBFjl6
Q4HE12JPR1PhGBaXUvDOhv8qvt7kSzQ6J1yteYb1sVbU+aa8C6ypZZIGeCMe4WjiDePB5WffUV6d
s7+WG0LQw3iMVuaxKmJNhQrVCwqCWTZdo+mTUXw4NidvkBrFxD4OHDIbX2V34qj4mj+rmYWcLvgo
wmlYwwVrnN7TnFtEOvSuRTaFHuzbXkF0IA+LEnOIkJC8XmiIa/d/JU5QChd731Q4Lwe0lCNPcF2t
89lJ+53l/emtQAhnkN7v9zCe9EJ7WQXhU0Gc2gZyVhlkakGJLs9uTMufUhsKFxEDS2RLbDTJzT81
O9JqRf7cUt85ZkbC+MBhMWlE0xCCn12+BLvYiYmo9VVUckL2fBboIkOH4sd1iSfkVkb6gwphi242
vR69pb0dnZE/m+HJrGch2w0rf4XB5OnfCGRuXN/xCtDwOd7u67MEm85OteDUBzhJsthCk+tFHClr
+tD7tXxxSquvI8BZ8M13Fj3jdFsq7QQ7nNvA4ZiiNHu53waemltwAIDZXsjusE1MqgZbYYNpD9h1
BuDbvcK6/g/9nkjIxqPX354Ty8LBp773/TyVBKkZlWmlrMsYgiaQeR92IrcMehV/a/b7D2Bi+VWo
fT5lLfrm5CYwfkzPpti+ubZsMPpQbHf/U9O2LTK0N1nkp8ujbFHSPoKa3bK5Ae/sP0IU/QqbJaTb
azmkD0TiylMzSa/e8TXgpiUlKqa3TkrVIa/Wa8E102nYKaKbT4MUZsVaz9znB/V6XyHicPVZdxVX
p9n0WNFUxQogYpLqVP8vTXpX2CFoIo0ZsmNN96XcPWUilim4a9Gg/nx7hwZm26YtFeRBQh1zJgqz
iEJn4bFLkmiqxR0eBiAATThDeue30YfgrQ+BLdtPdl+QFGBuNb3TB0NsyfkSBFpclwDqAGGGKree
G7xso6olGwJMmGNhNJMR6FJtEXfkX7ImYxrpZMnbwH/qCM7yY2QoBEcLaShncCgjHbrroyVdJztu
93aOaWjJDQAJBTPAaSwkXtFFQ1wLzmDh9yS7wfk8lE2XSJ0R9kp9BzJwWfItfw5Ur1noZwCW3Wjn
HbZ2RYHrgQQhQbtf0wqDsFNU99Fg90WXtzmJ1CKgIuuZ3+RvmZaeCjPa/23iH819IarYbyUobihH
HTRMgCK9Kt9Vyox1E5P/TL0WCBVQVEKSykh8Y2sOl5O5Z7Mp2N7cxGy7dvHkmJKg58CNC4N9dUgy
oqRfcGfYJuKGCLCEV/yT734++1GJVzeDL8VLbaoNYCyZ43RVa4G0YP0b0OEy6l76J3fq88YQcHMy
oyNgmukv2Ow9HILF0ai096C1CLgV3bl/wTjVooFgLqmORB9uU1BAlAYS+K/wtcXwvu8iKacuqdAk
M7sP4D1cPfeaxBRbnme9KEYMqT6MOXBHfoD+2u9z8GFkjbJ1gkQqujumJ/CELE0/b4ArHoieXH8M
ubkKPEWuLTWh7pHEP0/2Guq6Y750V3HmPjAMxyczct5YUbwZO7s5rVEPZ8udco1fY8O5g+gwmxZJ
ESz6J/PDxj7x0XP0QM17URo/D6PyYHqq+wA+rCK9gISmRNTLEZja1jz2zHO9Via0PmPjjQt0oofC
hzKvpHZyheidBt/XDU1scTtWH/CtIHMZe3DB2DxMicEZwue59us6WTmhf9WmBqcPKbMHPJ+IylTY
CJ09u04WhgZKkf+DxP8hptcbefFlFVSYQrLnrHGL4xShdhbytOk4xjCRqBwn7+uar0NyoNP/Si7N
6l3kVOxAPMRQlFvXCGkhTsXGib+QLip8XhqqFfYSmhpE/vIV9DWAYCoAEG2claFqn/6d8TneS8Jk
pznX4YGDn16ZGMyaq1W+Mbozqc6j2i7o+rVDiHqhcrromRR0a6dGVN5G9nPEpXwo9lHeKrwT60B7
WvwCGnekmVccOvPpkmGnUGSlT/gQ2hzA6alPx0Z1DRqW6IfFtCtkdIHwZ0A/6vuH3fcWn3+AypTf
fEGvtDo7GlcB+0bPOJXrGlF1rdsvnh+0U8lohxJJ0PJR0t1Ip63XkMRF3dFpp1JA0c+r+Vaxg5i3
8sw785U3OBnVK+mTeHdx9i1PFxvvX9yB3RNarLNvkkwmXOiSIR5WtFyVoch3EfetJEN9/K3UBADQ
RWUFJwpeiTwOan2eyirXPNpl+nCINoc6w5OTjT57KcAGLfLlX42z13ZVAz6uytAR1TvDq0jpNUF5
+p7da2oT+vMtwWDr4DcErI7+FDZBSkmaoFNI507bYP8Egff7GsgOlX80Us2ZV9qApGsoKphAPDtZ
gOHVrQHCh/uNbW+C0zL5wMQZuXdSsmMTuHuS01+US9JGuLM0aNpvI98p/e0TM2wGUG9RShDrGlOG
D5v6PPFSK1UCKfXTVpmAIFIr7tgV0ROHNl/DCghLI0hkePW39CnI0kAJzdmYCIXXwkyipQL110+y
eHQAQFsULtW0Yeek3/8EivjMYnr5lC6LomjLSEXw+qM8y/selQ06SwMTosV39eyJX7ZU53zSzwT7
gtPCSto8eX0+hHSMTGQgvqBtyhmIvvQqW+oaw+I0DzrjAVQ2JkO6bEIH1UWWdkcVQfegdii+bB5j
wNJEy28nuK+KEzzvb4xGT1ATNs1HyBQhqNr+M3b99uW5D7GEy51bHT3Khyx0l8yR6LRayqYzpRB3
ewB+B7kL3rmAchDn3qjWPIe8rcrV/KYCkJv3uMvhZYJbbQ11eJ8hphuE2ZufFWzXjR6oEJJrIBlu
aa+HVtNS8CepoiSUHhVT9Gq5QplfAs04ibxKU1anbzYFW8RVBDkJ3F2grl/rJTP1hdjfKjdTcHHL
EZv5bvp5WxayQ13fDP5jZrMwBqY0XMHo0FlAX5mq0LHRXniwdMW2Eh9Y4cVhjcDu2wge9UntIuAz
CZABC/tRKYAouvHjEBpsuVklcpQRb6mZfWJd+ItTOzN5pip/pVzLlcnORxkbEVRErTQ7LZkMhGZr
FlV94H+6Q6FrYdhcfCxRjGaXzW0VwwskS643F2L+IzUI5vRZhs8fW2zkKV7+313ehLk854rN+gus
CRdo9tsSy/aEVEsnuTPtGmisoV+zRa2EIuxKALnS2HATU40W8PfaVHEwVs4rDhC+sNUHw7cyQEIM
hzT9IHEQSAXusmL3XmahloyiDlUk9uEuUQFmzLQ5L+wA1UKcX7NRUCnFtPlUtjM9BnU3VCAvXa0A
FtBwjJjQeo7D6f2K/c6kIS+dfP98SIjJPlbZXk6IQUjBf3K+Ym1h8wojN39OlO41VsXQtQLS+Imf
A7VwRHStpMS/IsIrNzdeaOkQZMfwn2SSpF6bzBtjGxIcAk8zN43H7l/rdrU1b6hiklqHtldJZdm8
3ugbSSqjvnXUiLRZsccHVOX1Kco7BC913MZmsBQffBuB3zr4b/E2fM1YReWeZiq5jKgyA6T0SjRZ
3FGaoipwapJiA5G9adwTqJET4HN7u7bjD6BKWL02zprWEAj+/o2kUNomiA5/o5cqclIlBVFkpd28
l9zadCR5p5VXUvjQ+sDVyYWiogsqf2IyQ5QAzkQcygFKWO5/nPo7V1uYjjwGJ4xrMkjv8RftJiTY
9aADL2eOXgvAKg21RH6lk+YMiNCT16bz7N3UHLFt68I9SchNlorQ2phHSTW+KITGpyBXHy5N3Imk
Sojhywdm3JdAE+kYn0XuzRt89xY9Tv2QtRY7IHhdDX5zKS1sZYJPljS0SyqwkLAz/mgIOCAYl7OV
KCQG+BsKYnc0vpEhcxptoIm8Yxj72zKsDdWUHJNXWeaS8BD5cJqgFKJEVb7ODn/clGkhVFYyf19J
QqNypW/JfSJQJaxQsmwZMChbIdpCRfhh7p6YnMLDnuqonx+u/OuUo2QJg6TTRQtrIacBQ4RvMtXU
uVTkiowzkVsYplCq0CWXDU1az7ndfX6rnsnzz2NOXDBlc8kRqGIs+FVTEOvpMLbpMxS7jvIQvV/h
r/zHD0uwmncTIga2ZbFve2M59LZ9xkwLOisqfGPAnBQPQAP2lPzpJpb6Zedp2Gt+SA8sBNY3Vkyx
oUkpJrn54uiUAikdnqfoD6vhKA9ZkaYCd+QdHsFq0mxnjW4exYhunxNhRapA+GHAiaeKWXolhnYh
M0hguU8oB2HlJbHDrJKQbaAsyXMV/1WuaCwceceO1fu4FqP8hNjX+ULgB1HVKQiugFNSjPCHTr6f
DPpqbxGs2M2CS5+KA8xzyNC0QyBfaacjbMesfUe28blQCupWaJWu2EGw790ICsBqJ/y8j9EvDtlo
gbqS/kU04xiEWdRe3zaxe4dYb51ofnVG65pwoD18sdowq3Q6OsICsZ66NvVObO/j5+4kpcLaIc1a
5uXVFtdArJRZzYMOZTqImWtlNyYcR6EgMdCfqgdBawix5AuCVUCV7ZC83E6NqVoofuJpNlRXLuhP
MBVNDknI2g4R/BXqupj/6DWUHbGLLryoi0rqMndR+eaHsih/hf12iyR3tSwQBljDMlq+yXp8F9sG
bzv+7F7Cm35jJ/eTFePs0v1HL6N58Sb6mNsTvAcVz9OuC16Hg2XWvpqcfnatfhUwgVB+QZ1fpPv/
N1a69foMoTxJACbGiNt26FsHQ4yKHUqc23n9jQT7n/jynaD78OWcFH9HljZmGweo4VxDrpHlVusK
wCAjq9JUEIJC2KugbqtAmW43pKlInxcTfbpS1rldzZ2pZXHKCVZrjtJYXZLBhlMpA34BbHdp+AYb
K4ll6PzWhqDIifP+0T4/+BSHnJzxOzQ9Foo9s0dOSmkF9YZD61U63UKMMfWwjjW1nSGiL42WSmih
rnXqyDE33fxwESzhXyximQOqhiL+/TYWLo01w6h0iX4MW13FPNhdunbXUVRE4nYKFYlfCLOawoxp
55Dj4H954S7lW+lEdYYsCJHzdgdZ4xCCeW1JUTE2wjiz5dGIPZp4tKDeeNA3sjr3iwGH9FNRj5E/
SFRgmW436q0nMATVAaLFYrPtTBJhT1cxHe9BVfXKoNAWuDrh51XHZ3EAM69wadmvgUyazHmIzP6e
MREOTFUQauCoir8mo3iaCWe+duPAC93npuVK/PB6rx7wfJxisR1GsOPGUx+tNy419I5WMVCZbmIM
Ph+/BGTYtZ8fh6WVKEuQdARXns6VKcXB+WT2JZHnFTAjFm5O4d6kZp0jZXixlIXuWekNeXdIIrA4
l8gD3tyMEuz/o9O2brKddtBCWLJCKaiqTHmE53JnsrFZgEs1lyOurKtfHxuWHvwKpM/+OZU55/09
mc+8QwbBpTQdUukOJOduvONB/suun3i79jM0rEC3goW0buc1MOMfZJVW60hrAQjdTIUo3qtOv7Wb
TQw6qXKlskNHZC7XLnpay+8VgfGZPKsu5Cgy1aTiEG2QzYcHWnZc8DKjhr4J6FzpslQH/i1DJhYn
Ge3s96Enhmg5TA+8clvNJAuCpJhdntFfY2YfZKv1xwOjvnbw4EgRRsQbWgAecN0u/qS8DHAZ1xP5
8BPAy8FdUiJUQMqFyb9oUuUpuW6x07uUv5/HKTasQRKYBKIlLSBZf4s0bnvekw6aPgwPznrznzGW
qDzG4t54FNz5d9n9Xw0JtsH8OeT9EOJyfrOP8t8VVvOtpbC89YLjealA0AUaQmSP4aQj5LNiyIdT
uUXnVH3zeQR4ORfptD7yvlsryzWhIj2ACkbsjBTLC91wMMQ4skv9ptFDxlAjFutfdcDbKvQEL/BU
a1XIrZ87H8zD4/LTjfOcyhUdzwFJYVP+w2Nnw+trFtn0oqyQPjCknqCfXBovGXs6bpVDbSDegs+g
rKY1iaGAl6gnEEPDUKJQUX2Vedj5hHUJGN1IOXvoWuNuwRQ3Xy5KKaR6UBHoEqDRyBVnb63HV3NI
C5BeG6br4R4ScPKfiWKw/huJEpzNrtwdgzuU5VkRtj5wxD5wNzXTbVoyQ21RIKVvjIcrU3Rcm3E6
te1XAlLfkeSYcSv+1jouNvxTaJxAwcwD4QfI8Yv2rUAj7t6oXgCryCOy80RbHTwYX8aOExmw1V+y
XssPIiT/3yhaF+QUecw3dsxYY+4sgTBEWlXUCq23PS1jjcW9eIjeSaFSYv9VQ2AmZT/F3vy68iCB
BpINL4FW0Q90mcteZtYuWKq89x+EGWOmOMa7rOZaz29Em+UuCYVvEhgenz7WYVff1wU5CzYd963P
Bcdnov07Pf1xW84xd9jikkLO/Ad3v2rP6wwvcFRNcogipbON3iUW8P2ITie076CtS6QbMUwJ62vq
6+0yYpFGoT3wVgnGXLAbz/LbX5BIDLebsSQkfvejbMR8dXlhqHM/bYk8RKrwTorO8LsqN7KHMga+
SvnvG6TzR6g+9+PnwQv/fRdlLAbLXFl8H4jXIyom3xusPsGa7/4CgWIM9kjCxNseIINMFAjxTFBv
MD/n09x9xlhRVGvS9/dvLdZtQMhLFc7nbw8hpop6aZJru+a6HW5+Z4vPgy+cgbgz58LrJghckOid
Cw5CEcbTH6Cb5cIJwiBIr5OpOf+Tz9xvZQv8VsjSRNIxlGV+YexNV99YC72zu5/MNT5gsZ4pGVI0
bf9vye0AsLeoPWozlwQ0XetB5NBYO9xB3LnnjYfqdWiK8IXKXZpBNelg8egrc9LQ1XwOtCdWi9+f
PV30SyVgL/bx0yReG0vmc/zq+iJYqY0wLX8lJkAwZuCJJkjXoEwwMXcDeA0l3VPG8uG2sM0pNRYA
EabUrO9XqkZ1+n3LLql2RDzYBxd8aUqrM5/PaHtIWndvns6+w90fJ8jSqU8+bRZfNAXGcYGTLaMd
Ofwg3KVh3QCalyAUVNPU5ZxXuPJbQhfcXsxR2QhXLjxk2xZZPaBGB8i2qBQg88LWpQUax6g1+lG1
ncsKxErSn2Og6NVSkQ7p3pE7jiO/V0UlDYoscGJ06Y/EF6UWEDVV+2l4b8BKfX+WFS6cp/P4VdCJ
tODHhiYQDbCRXD1YH9oyD2WOQJZqudvWMKyePSm0nAPamPWDb/MDcxvnPoNiV0RHt/fhCnLcFPZs
NLK/v6CFIhW6M0h/o7udC1RHTJaTSNZozNb6o219Kcpo9afIuITOpUXs1KR/Kgyh6ABdpWbDsXyL
KsTzu2a3FGxQH+D+6s2lyDLwUMBxbpLee1ceBL+S4w6IjMUCswXGAORgrsGO6eiQgXFBfNSc1A+c
wrjOE5JAs4odNsF5qRo58x8OE6x8pV3Sm7OIHGPMVW2IUVBPEQDmKSVNOal1P12f1OBpXMbBndwV
9ByE73Yef40kU5j5IUy8uLDHeEKOYJDnqfiV4XyVCOx1PXih7Wp8YPor7OUcCTbwFZO4TuURoU6/
WCLDi6qd257R3DxRA/TfwmbN6rGTpsJWmN0rV8MviDNcK9iLHIOMAs3vm6QIfLXI35FdDst6Yjl/
80GD5OsLXDyvZw9qocW5CqwJYNwivpeHtYfaTCsA/k5KqCJgjjDtYnRdmvX3AYB0NOt/F49jclps
OXNLeZPyPcaoHw44BKHUtTMwsYt/2MhKvYNjd8VVgeOZ7wup//Kdb2DA+C0uvJ3vJMiQMymSorAw
PKMwXQHCWZ6WJtgP2PWd3N2eWZQP5ayjSium6HkG5MvzspuThbTuJoPKuQHG390LBzBr8EL9S6Dr
qOctJV93S8zrzjAhkCdUe9Llfv09l63LTZf3wjSnWDSnXZnH84nv/n5m+gzBXZCq0xbMHRFH7nZy
jq/IxO84kQhPJqX4gchOgqgT/ec96hRWK2n5s4ZNBnWhqFVMIlSTC25L7yYPFls5poD7WiOKsg8V
JtPiGbPG6DfW4xNu3RLWUyfm3u25EOBEf9tBD4nFUII1TLAMTUEyZQJVH6qEr2zhYiHIAaNcWOxU
TImv6RP6tyGJ3TnmEtX5kOSTy92ShS7xPdrFTS2tf4jkHv5u/5+BBKKgRBgOWJLe2dCDHio2psCR
2KrQJ8j76MgTriSd9wsUL2CER+PtrfFH72AKNgCXCc8/1MFnjBsjdBkNMlt/F+14Q6SywY40xba9
2aNp++qBDxU9G+wVI1Fe8sUtz8feews4NI1irqjVtz/S6OGXY9kznG4Ic4OJPC7A3fHcwHxKVDZv
/Ajkns+lk6UZ4YH0f+zR14EjaGpa3+8v3JQQVb5PS+rAR0i9Ig/H0FPTyCBrVhAOehtNrpL5kCQE
1/nMTS+PVbNUbA/DJtkVTd5EtOSjWNQEIGRI+6ZprtfyfGVZJX1Vfkc2fLevZFq/AODOEIKbXQ9X
NVQ5evQDEMh4omjWmoSIObkCvdWcRWrG4wmP6JJSZyawaWgzgktYyQnuxmmFuy2ngt+JN54GF2QO
kT5SKZIAd/xgiD7wU/gqHz6aueh+hZRVDixgm/5ZO5YYc72N9Mnz73Z0/yIuE1VnqrrQlycp1fgO
f3SJNaP5SdKZx/JdmdaqQXXZ1E3uREhGyas75HRkkURSwG/IqjHg3Ew/QsNouLyVVO7kaEcUyuwg
XFJTY0p/QbTMnXF7DceH1r/3Z8yELMYzdm6VQGS2MXEtwwvQMNX0/dSli1KfwOaTiLr8a46mYfAK
INSmSJOBwMiGYnGqIf86lKMZ3cxDKuUChbMLam3IIcNFEu0UuHQ4HIfyQQI9rap0GYVRzifQ+xaF
flrlnjSeC08e+zyHlSr0Omyy4s75Fxm7rOVXqyA6HFAtkSPxBU/NDmFQWzL8c6kb2s2LK8Q3Kr7g
zrLtq4DEO6eEzC0gaJ1Dd7kEvu/5/SbbCnu5WQIBVaSge27hiMVFLKNUOTKnUvlGs56kb8rBTklh
wTa5+h17AkmYowqZ1k9r52RdHDd3epl1i1fHkcVFFiK4YIjmE9hzi6sgfwu7ayZWGtA1pC1jUdY1
R5CcC6ZeE1pvL8RD/m6gXiaxEd7PM4uoWxs2sjKkddNczIksybzmcTLE8lkM7olFUgw6dkdvMvSY
5Pu4rpo1E09ZA+kjZuXeAJC8UrwTuqWAYKjVFzyPQPZxyUPxxPlwpOvOtD7zTx3gQ/FT8F89zoff
Hs6dqqpeYmLfns8QmBbitqIZYeiiSouzewmVJ3BkJqlSTmjwZNz+ksuBirN/EglkX8J/423sUAT8
4qPWPd1PQ12Cq8t0WZjHI9qVYLMfKs7gVSZD/nzuEXMgRj1c21+srxjxsgX3F6ml14oYNpgp3kvQ
QVr/ZAqURwlDuwYyxddQOdK3ciKYqlkThYpJC9C+H4gqG49ZOH2fppAb9mtvVbvNam4MP4J194ZW
RmcIogA7kBVujOv3eTGk5R/hAD0rt+EZmKc7Es3shGNClIjuhyFlo1lH4eF46fh27IpaS1bNsLau
bcJXcLo4Otm3VYQjbKsDbLSWPyOhVMlhK7YRxTKOLJsLTUxTpicg2UviTeWa4YeKN6Gqq4BE36an
97MjSCZeqNq5EkBjVfbAhs081Z1PRtnSW/z1m5iclMdOkGX0kqCQbTUV5U+TWRiosjkqt14K9Tjq
qYz8i7jxM+Bj1Xd1i0tF3pNSmVcPzrvJYxcGvsLzWweRzmBCEry9EAkOrEo3/KfjvMlloU9w0nY1
2sLIAczQxYJB9iPY3kz/MRGU0wUQn+wVYHWKKs+mO9fX6RBkS35H2g8Jmw1zN8PXFRMT94gg33ks
upn2nJUHe1mOBZBUyVymTOEqOaspwodA1eY6rdhYl8ucfJYgVc3jn7NXDEPBQkj85uCIlQpx0fL+
doQb8nqr5rmKSghNt0/meIzGzkCbOMI5T3JAydMagReNytL//Trxvm0KOE6/hc0OSETo6vBrlJgJ
0lxl0EpUKYpUxl701GE8hQ20m4Pnm2eO+M7tl3WIUaxYcLhWsyztwS6mqOJQkgpDEj4nV9CE4yyi
iSii27YRCvJr7K0VniGyZOOtcoeK2+/+Lyngzf7KEw+sxiYr2+xRIexltedUPY32Wsd0jEtNXG0G
+Ltx7v42GiG3HJKiglVmN4qQWXRqWJ5DwudJsM2dtg2uDD62lqc1U26E3hGItzaoxU2nhkFBpZUj
DmpmxwUcJqNoWexSGH4Yko6Q0Lx2cU5U7y+gt/sqE44cqoO7LxobSHvd6hF13+nktJeiN42lVdQS
5q6bBF+rPzcMiHt/DIAMwqjNPV4jAooAeb6eorZDOD29AohTScCvfYA9kSSkIPL31EtoJunsdw67
SVzj6icetxPzMCe/J0wplPITEIJMkwQGL3iC4x+wO5p7PofokZL5BIEqj7ZrCp3FS46FKp0+YRdi
FgAJ052FPvplRPWAAJpN6htkUptFhjiFk0I+QTl0AdZUscO+4I+Ghh7ujBWFE62jpgR4AkSaO6Ho
R5TSitTr4DgKZfuOA4m2N0Xa5r4TuGDqbiLAzW5YxLrYNZtsgYV1j1MAuVltx2qxmyW17Tek+Gok
pD+M1Er2gc/HSM1zwJ/CjhrNqfqiCqG2JfD1yTDahzdF+ZA0JoDlSbbngwTc/DeD+VDOW4FdKRuF
+VGfnnh58+9e3CZmfWMY40xkaNF8BnuGQIXPPeEQ3aY6E36rRetaLJd/UcyPQyqVwn4dPvffR3TK
0xtsgSqzqbZKJljejUftKGze5CKo2RcBFUTV6yr82mwo2Kvi1KM6hlk3N+CsX5EYJs/ZCI+URwoJ
KdziI+5oD5z/CLbO/0R/nNBW4F73WJyubIWLm9Gs6/csAShvhOEyaC4B/ZqRMuZKDamKCCuTpqBu
Xvy5VKfaMIhPFSpeT4YF7Wy2nR6UCvGT88YuHL96FGqs+YBTrX0Vc3PcTNQe51u7PItbH2S4mH28
5ZmiR1FM1x5PWGjbV71bzIcmUs/qqv/4RsdMdQCFPz+RUn/7wB77QGMccRtUe0H+MQdgTGHvGErH
h/M4OnZNrvaVfZCtjB7V3s6jZ+zkbBHD8UNsKJcajIIYrl3T55UIx1jCdT020zMSqQvYOv7PnXZk
WbxFS56em1x4YQ/+HMY6DR4bqYy//p3NspCrKCRgmV9nHDQ3TPh/azbvlCnlK9fpmx+GJ7fPPIAG
hVEqF/g5fl+dS355S+w2lNtf2P2pHLdiqbaqn3wkEwlaA/gHMkEDGn6GrwXy7L1cV+wTCW9s36WU
pbfqdnBIWCBV1gSQeCs0Sf8WXAVpMjYjMOD03Stx3lq9uDPNzinUNTqGq4xO9RbJUXCAOEnoybU0
21hbVRgXrwhzBTBgWXKo5NrwQLcYOWrknZL+BEBb2eAZhZaRlcAP8WiEByy/WScKSaSmuT1fO0Vn
SnWJz0pIleWONpLsp8omi9h8VDZZG9aBqLl4SIl7PCkxNIjTDFdP/+ni+LPe+rAkoJlgY1QFxqjt
qh5sMFLf4Iivarh6S1caIkI/UxnOQ/rVxN3Sv6rEyJlSrIGo2u0ruwCfOdLH2ReEM3rjIC9ZrRXZ
M+HtM5A1s0Q2+3LLD3TaWsslo+or9cuaPWqPasREoL3TxbYtifwID9rh/QLWEELS7pSSZZ9HKJqF
9GeFg/+quDWRq9stoG1Oe34wcUWyWTHUjgNYnnYGz+9rf50mQiiiGbT6RNojXwIu0fRBk9koOR0L
gZ7zrYCj6Ke4S45zGlOK4M9czqbWiYNdsBEbGPhA8yu/BnV2W8M2m9kK7lj9BY2xj3K6tvS7IBid
dGLYEwRne15EjDl+gaBFTR1r3GBwlpmKmd7dDq+ZZ257zNRdVXm9Ln07pcBhi0FIhyzq7pwJtYD5
B1leQp7RK3YSOSDxvMyoTe3OuDVmDeIoz3nQ3osE7TUS2K2+B+g8gb1vGZzv82XvfSjlRPBczFcp
c/Y4nwRQM/la+g75nlQEnDQoe1M4p5I+XJ9maOaujCyOvkZafsr/FwVQ7NH20iIuMO/QfzD9k+Yz
usNmeMXxk4umvDC8uw4nqu/msjc8EUCDp55U8UqPGO8LirpDG95OqZu7e6vcgPuvMuc826T9rEhF
xmnQHVBEBulnJjBc8JRY6Hn1ewWIpemM9728Vkhc+nuJ2Gp0jHGa+82Fy+jif6ug8wbAK/OzyH7P
hSA7uBMTO0rDA718jpKR2ZZT0W0DDaKzaLuuO9kPSX/DiGI56GUKDUE8gO7vGWVXE9h9Zm11Yims
iWUlmNTyCp+ZoMzhUVP4iEfam7ezMI6sDJ/7lE2AyuEG+95Q74GCX6P3qkO/f46oZyj5RQwGkABZ
GYjxN16WW9IWGDec7M0A9Zra64wpoj3Ot3nudNdwyC/8KKGE62ZMk5l2fYysdcblMCzpcANXGUqv
r3pzLZQM7OM9ToTJHAlLUhfT4QAfVSF/HwenBKFJR12/AY89eW7xZOx01hRR8mym3miDau7t/DV4
/Mr97X9h2IWXtwOE0HV14pLlNuqcZsrAbM9aFl+wAT+VXA8CU7toUCo630B3sUJFmMPlfHbOqK4B
LI8BPpTJuq9NHB6JMw3x6tUKEHzoJ7pThPVUbjY+g8eBf29PyvDQVH81dQrvx1nn6x8H0fyGfXl0
klVHqMgNyl4zaK3R+3J2NXptbI4nlYGSsJ537BR0nXf5DQXCwwbsCUuP6RtT2nKnDr/0qqQoRbbH
lP/mowt8H12erbAZ2o5l7AyKGV43kC+eqVjllRTD4+PBRsCA1N+6nzbU1EUEEbNZ2VX/zsc/7HfJ
D7Tjd0n9VGbl2PucDxcETkM2x0tILQ3F83cHPUJYDsuWE9mQDxGx762VEXXDHR+bfBYy5/NBvR24
0YizDYW8ffxgSUK/U3N0VEhKBA1NzgxJEfyuObHZdQNE0q3QoOC77oKorXQblYlI+YqkAA5U9Vlm
WxbFNykfcADZzRdJfTjl8Vo16XQ8Wz6Inoc4G7aqDFAB8YQPvY1+TBJFl0iG605BiZSgW75LIpNL
/NFFCW1Yexz4xxLlSr5Q/VWe9YGDBCingGzo6kPYicXcy0WdfgzvGYPkPkcNYKTUE5Y8Sl/qPyLl
8m6Yek9T8mr/ibjzoz8YSpWvhbAQe16hIoccQzoYU9C6H7xzEr385QhE6rTnjF0lVr45zJwFFg5I
38LR43tiz2HX6XdjbwSTZo860dHS/oc+1GSPYJkUgGOv7a5T5EA/fu78xCiae2JT8xEDQVrpKrs2
fDwzLOFkxXFs/y3tnZVhgMcLeSkImb0zWsWNW/uuvVxCYbuMGjQFsxhEq5XfS70FCXBKkg7VExyA
pl2TtEZEtsuUaaLLQqu2VT359FK4ItlvJ4Z//L0hv2v3NmPv8lUhOadbBB7lva/2E7OSqYakCQWv
ENyQwtiYzKlAnZGadwlJ83mUgFBa5zqX1TAwEKR48ks1sGRLMT0HsMnLl/MZ4dZ8M9bz1fYsP/d+
WAgLCG2Zu58cSnN4YgctIEjstTZUtWterDAGaYMCYuXxaBgxv8qtgDJqx+1DtUDQ/jy6RE4ET5Qr
FB/P0/EIwzIjTdBPXWLT6oJGc2fdrqc6e3Ed9H1cqQt5IokAChOY//q64Ozn/2Po8GdZuI35d2e2
iPh3FR/pru5rMJAnTsGXi2YWdDq9yXH0YZrYBd7hRjhqEnMk7l6B4nbCg0tab2hYX3QhUTTAHJ0G
qG00d229mo6LKhqP8Iq5rPg5kRe3/LnUAMWENnEMuoPMfd7J+ASlNtBuFePn1QMrIIbKjxHxSCQL
M4X8I4Q9hmSx7olA0sCsen7z64Pu6sflRgPv5onYrT+DGfHmApXT203QQCJ6zp+pMgXWsL5XzpIe
IPgPqpJLxgRxBiE+wS+kJblWyP/U8ygv/N3of//EDhncXJFfbfOUe6WWuZvQ4uJlxzvg4CqdPrrS
6oqA8ER5aRzOOvXtibWPBXEKC517CFRg03Gi6Z44n8VYsIwUQ/fOQ5LCpxKN9WY7V/WAkyc5wXrf
CB7+ZWB5toOw47yws3WrA08h8x5tgm+ZM4B6YfFJHg6d5B29gAaD4HGX8MkjVioDG6f42IdTyQgl
zKMKJhrYLlRhonES6roPyJNRssknscZNTgTPY7FTjwHy7IqcyvX+1eTT06J4gPXOcFCey4WAtUtw
3yMA4VagU0WUgynjT905gf1hA4cycBwLVGan895RXFFy48X+FRe5FH3SQiEeU1aao3pY8/BNFekf
FN190Ix7iUaLbtzN6BzyeJKZhNfG1Fj+19zvql4xwXYAPa8Gvhi6B4TMX3BnndbZ2JJM20pbrmgc
3uK8t05WZJT8TXZiS4JsCHazT7i1Rnd3pItZDvyKo1QME8NAHu9YwajtqbkYeBlaZvUpe+jAFzQ4
a6elbTU11pjQUs9/jwwh5PZmS6j6z/PUU/NcL+bFLQ0QiOw3JTQIlselL84Lo8BUeX2oJZtzYa1u
tdF18egDNsUIFnHBqk1u7iaYeEefg/gJW1+1+ScHh1wkOhitf43XIAdyRWHElY6t8bti1jX+VZr4
ydnpdZU6z1jvldoYpC6PEs7sJU5hwyDoQPhd21xQWHYGeASjUNAvHPil5YXA+DqaDwdZqgiljlJN
sIDoyALyLijyuontZYe0EYafyPd0TsEQLY7kQf6Z5s1IyC4eUSIlhYrjkJvG+tbapG7sc5Idb8Z4
Sqy3TdX+x5rlfuzjvm1n0p03/VscKVVAx6MCPS87oOAWra9iLHeLC1hNyOco++y2FZaMJA/bdbLd
taPDixkmOkpdUDIwQAHXLMZHM16PIp8GqHeQge+gzBNbRZEzI5qbHoxFJtBKP8VvuIRRujFIFFGd
+9EtaOktYjKWzohDYy2XUb47EJXngXWlk3m41BY0rilHYbugFUcA2kBM1hbtTBqK2x26Ghi5fsZy
oWyiFTvHXj0ZZnbzL9gyZqIZLsX1XXStSUvZE1mChD2AAdkTTPOtegmJusA8HIQY0iUKnAS0EpeV
uipa8w0Jq85ABLxXTURSAXziAE86ZAejfLNqRQrxYMQ4dfRgg4RWW7sK8hSBAjlSnUUnpbps+jc6
d+M6i6fgjrJYtWtFwcnyE79JE/sJUsd6j/25AZVS+DUBu6Ok65V7MgAKno00hTwq9a4a9tlZ3xp+
iKBW1t2BdX/gi4vM/QCBN9VaKw/AU8UsSe/mmehWMwnavw618v4bHVghtclMJ6J/Zs4oLlLQtWAD
1pLk2V/vQOSWGLb0OYqF72RnGs25nkdbAVt1kDFf6Hz2O7MUODBsIi+PyVP0QUC0WbMFkHPg7TAZ
7qBYN1Bi8gs7hzthRVsvw2EdLPl5Ifm5YyGra+zlOh8UgylfEVFOjPNj0E/58wndS/NZt9ZTyH6I
MEX0s1T9l8lNQ013UJn8znAjm/koL4nkZfIMvlIl/pDTcubq8rnGg6qTRWhI8E71HUSdM1+9Km5f
h6pzbb/KC39/bxzCY5Z75cU67YDeuIkMVktVwc07oqBoLUO7FOOycYT3rRi1DsL2I3MsWQW1fzwd
E+Ubp/ca8BxpiWyFXp+10OyuxPrwKIuXIN0vceQaTiUOGa5t2QHuAhq+yOBa9M27sI4OTRu++x2M
MMhNeYAV0+3oz4b4jroHocOWNT6CoG/SqCSbjdWLUpGnHDCzIGHUrQF9UyI1Oncn3Sv44b7Ts2Xw
cgHwnNsj3FvjG91HxWE0zu580Db6BgBL47WABVz/OBEmS3KpYx9T/P6NzKp7Yc6KAt8WQFugyQn/
HJ3XUehp/UjJ9uSd5VjnFHmZIPamv1aVZrROWLzJLcmwts2AKOyN5Mr70tTuPlyQNEwsyyyUsQFa
tJvftXvH+JqsikpTmLczUz/BPRkTVXhxDbcOfCovP0lM1IYksDxWdkiEYowozoIFOESJ/mzkGcEB
UIUkLXgbDwNSnii3QU9kOIiCRA9yJzio/z0hpndd/jakKUUjJ7FkcnT5vuF9xcVB5m9cvQf5+SJ5
vJkZn4krCrUM4Z6eBZE9MgOpFiYEw4GSHECwz8OD/ETBmkOgkNPR2FD2xi7rFAjpw0K4Vub5YsEp
XmvUKfSJGqc2FApV+9Z4ll5IFJLvsb5zxuYWu8YSUHQfhCNEBG/6P+sksINckoM6xlYDPjADkMjG
f61A9t8cx00Kin2ym0UAytaXeA8XA64lTAT/3jOI/L7p1gBkE/47XL4t8PtgtMiaJojo8u6GMzyL
P6IE7q1bX5QPq3y16oIZ5SuAE0EQiN7en0nEu85hnYcWKsYS5wefquGHwDh/Pu88m6+MJbo1tOXm
XiuzfA99bkcAz+KtrsHxRK90/1sgsS27ICka3sxc0NEeNJAiSjBykhCA4qPV7gSSZyQ8CmJORBcb
1evvaQPPmJ6sopgrrpKZHTdgb/ETQBnHfUyty9xavkU5J9EflD0GONF4M9faLhccAZfPnnJyzeWn
5oveQ4U4WXU7j2ZjjTClNByf4BuvJ9znh3UHKIcJxgX+EePmtnKKVQrwSQQ5ymBt3nEUFyVFTUCp
M6kM0T6SUAdB2CWY1PRFiDDIB48GLA+MpYkOMXrfR5G8oEMXNH0n4FOf2yUS6eW989odkv08JqqF
ffuIKo1igAjIx/mhpGUZVXwY0jKdxLp5YZ+qUWJMYUnghOKH+wqvyuY1QM/Tx/z4yqng5oZQqlaM
E23VOWaFUeKCgmveWPC7EtZza+knlquopsd9J0aXKvH7I9lwOOVbe6moJ+6tmBuAXvhnxkvyTsMv
cLIgGmAu6QiQWN4nYfPMtwWaffndUjYGvNq81mK++PwnM7cD89R3K/IwnaFC8JguQi0MgjZ5EXUz
Q31KffyQwkLGEWtHoF4gqrtlV37sBXv3auq4ueiJKyBj0P0XfGDQQO+iRXTQnRb9/8RLnuZZrzsx
NhSQRW0Xuv02p0WD2IxWLCRMqVi6dDeNzrBgJUWiaYPDdov3tq+ittNH2DVZTIosBnH8ZRAbEPcD
bRqLZ88FhimXFIjmXc16584wSw8TguQJ2mHW061Bu9AAUAAoUB1gSvSq25pPbY201SJvwAzxl4dR
2Fl+QTKnI34aTcDWvpBHrpy59WwIjAgrDc53swRscLWuL3UoNjL9x6tXyWsttJEdwUy8CXLdZpmF
iiyazL0CsOvD74iHFs5s2PEJaM3WNXeQYKz6IYfCQLhw+9sGrnjPd7hza8IahJpK4UZU9B7kG6uy
u4BdZGbcu5waXqnKFT+6x1Qj0SU07uNs0s8X1K+JPXSX+WhdePdPIe58eHc5eg64As5dz8UwT305
nxHioJelxqjeSmqxxxONMwvVy8mlq87cO9crAAL7fFqXGy8MbQ1hKrvGAHqtV9KoGELAsWVCvFh9
eVSUrLmWHX7QMh8vjlBE2A2ULcKrl1SIAgPFhp3HTZHvz2hmeGSPC2TOtho4h2cLS+UVve1HETV2
NQcx3A+0V0uKDnfeMF++kDLBUx/41HTy0TeGchz8KuxEbvo3THmGPQYZOaSHG1/dPG4l1iC0zzZ3
V+zH+EAUKba1UZjIP2yc2mOjWIh+jjQjpnoUeLYx+KsOOHNrfE645DVL0jiryvSlPrSJ1rIhmhfN
5cOlGB5rCA1LcTRUavXeBTz6sEOQpmz82ex0K7urPz+t7ydPrn+Bz0ZLjGTvf1Mx+PwVrKEUNw4X
XRzlYHN6pkitzq6t4pPs9EnSqN5NFWOSm5CdV6aoicFBR8Mal0xDgNcF1jGNNtlJip+Dp87Wo4uo
TLlNQnntmADPPah5H99ZuJciOblk/hRHdfWd811/PYiSCk3tdMa60lUz6uDqKl1Ey/gmfDQxdC6B
ZZRZ8XKhV2jKTIYCTwI8IeyRvAkUO34SNBm2LGHAnV/Z7MnF1KnX3ufcIOY6JOetTz5CvQQYAkaq
QIdBbIw5wxYOl4eLXqkaal/YsHOMnaKw1hjgL+zqSJegPRIUIYwtpGc0wh0vOsl8HkchEvHbXZS1
ugp09aEeYk6zE/FIqzAJxqdeXFU4zbvrEQeJYFAiUYbiwac/0IKzMVT4zIdTUKRQXut0e7lFF8yQ
mfxNZJFYCRFBGEHKEm1lX6Du+u7LGuZMIccVPnjGa7Vxo9NcKr7RPfLlcqg4lHxnOmK1kFzy0nom
bp5fyEhVxoZ7vX2vn/D7s/38QopNZlKk9gA/KKS0jPSZEp9z8/j8xisKb5BElXK/J3Yeu9FxboCs
slmvnmAgJIRbKorZhhugZWSr2yqxo/66anoN1RopO/XM915SHkcSxnEjHEoqKRSEdsAVYSeWILb0
JnH7A5EhdfomEbcqVuJjkvTZ+rFaJDQUG6ZrhhBAukMp+Za14dCU6JCfsFu+iFUpMw63fBZQe31I
DT1KvQaPIPdapj95Iei4onsRx7VADDHEeW5DbYHT2P0Nd1WjHZNH9fr6Ou9FxUWJ995EkiyOOCNI
Ta3QFI5J9Do/AhGGLQ1koHPOK8CcLVDjBWlVpyrfY8n8Ry4mVLGb0c61okusCAZGg5rvxricyuQu
gt11f7D+3YlyuunI9QQAIv2JAQh5FrUUyOvwiNs/fXQPmayHEvMxvXyqq8MDwboa1NVVR3YpjrlT
Gpc0UAhywPC0tDqooY8CeuFPLGMbzv+0GRftMDq6cM+O40kSKWBnR46FkP7/KMTLjTPA/22iKE3l
E7oUPvSV6558hW7Xqte+Q0N1D4LOQNLDwVUJrB9rZJPsh18Z8Adeqp8EXqNmN63NcRpO/dF+bFo9
OJpxP56oUxzYrHVP/Uj10oRLj3jWCm57xNzN684b17t59UVvcF1RK+TBJO+bni6RWyroW/STScya
xidAwIyxFqmh0hS1mAomH9oECylrTRQHXstVWb5+bJHqELl9y9SkIcyrYi4gLCA2MXzLl9ob6saj
MlfI4yVdpPiHfrIsvMt2UNSaLkIypWRnb75AVcNO5QKXv6xkcBUGGY2wpyXFUy3ehj425tFbgJeA
vhp42zht8tyA5TfJRaEQwGHl+3Mo3fozWvIGeXKLBxYbXkNuHstPwRki2DYTsjbto/l/6w4iUTxn
nAQ5GAL3/gM7U3uDCbzWczzng+LB+8suxRGr/2aK1VYf2wWjwOqtZEpa8CySDjdmyedlsZi0D50d
UfmSD8TxfwRwL/HRC01u1qzuE//mAZbFQZwjl0smQ7DxYEtJEoXFEYVv7DGM4KpIrZeN5EliXqQg
uDES+bd1xKIbLgsJqO7zDImksCLRCYgc4BMenVijIBjuQlsKOTmXRZrisT7tH05BDUMIRt6gyWFI
IhBK83fH6Jh6pcuPnxf02XPEPSr+rsHIy6SWbP3I3MBKxrz78emJvoZyBxaNWTFRRO6b93O+B8B9
mOJtWdRIGIyqtJDTDPQ8ATkvrp8Ati4ziXGae765WV4U9BGBkpSfPIBxVt1mUQ2ESdIxGzz1s1fx
3xfqN8k2eeLV3gUOeLpbstEGzCCZeDyYwHKzHh45YZKoUmhmihD4U6YfddMxzy0qv7vsm/VB1zfQ
gsbRiym/ZB21rci0cPuLBmE4HwF6NXsZ9amMGJ+95DOjgofV4U28EnLzd6vtFBQhrHd//dZQPudb
ByfEmkcZQ2mV94y8SD9+8AYBlhd7d4JJSEU3tXCKlCyt18xSIBXuC8YpuNAcIzCcCVn4AXLMQkaF
8Tw1sApoOZYNp33VOrMoaAWvlqFOVN20XL+jLmVBVTcTlAfo+C4xcOPsulXjVpiN/hHQMq6qHSje
ywGPd5Airey02yfZ9Gtz9qBIIktYlGaVImJSNUczd3DPLHHkt3sfJOlg91f9CivsMo/tUPNSV6Ob
zDr+r4kVMgNXgsDZ9Blm+iRRpxWO7+Fqw6CzMOvc2czHCpoPim+8KiYxgnhWiswvRwoVUnmxTyNs
nTTm4to8AcGeyT4FlI3T681JO0wygJAVCSHz4pQ17TEtmzPDnaNUndmP815m3Q/K/JwzLAtWfhb6
TTUNoqm7GmPfESfaZrr/2yZnVc/E3belv3Xzpsl/NOMVjtAVq0xQ6RFN1HwBmz1mSMUcz+koDpli
dgro0XLmjJe6vUa57gf2EI5j7bIbEmNWya4DHRE/8k/kso6EE2+Jpgk3otiPbpSpYCtMSBMvA27q
tQBACmdHN0GhIGfXrXFuyBOPtEiC7JnydlAhOjGCdNy+UV1QofmUktPOu6jPjbdncxbqGwezqftf
LXWhk7nxNM6bGuAZDrXE6wbi3NXaRwEcdbGLs6N0gY9Hdms2SxxUApT7WscquKwg9sS3z9rlRAlc
LCb7vRtlOopXbmeuNLaFB3b4vTaeMpCkAjIHtxG/SakoNqrjK/5XIjh6lbV3TGHFl3y8OWGFtVuF
g/XjHSCDP2yvm2G87H4XOnOazesFm/J22xvlZTOZxlXZEgaOylY+6SH1Sjgl/hHTpKZ6DgVvAR+o
+KJpk0o9KRTrNHIdKN0f8ztnoEo52jr8lFwmTSodclMil2qZhweTSqTdk35PeUKmVd2rbcAX4wX9
vBRfl/e8o9dTxbPE02/LJtiYMr5Eo0WwRgutR+6qWV99NUSTpBn5VtYCgeG05lZFPa26z5QEBWMt
9X9VnyCxCFVYUw79PVUieaBc+JVNtDcLgjFAi7YomO1eB4l7V5dJ7VeErbeFGmAjVJx/nWmCqYCX
03G9Vf6zKeBKrvnixphCK3wU5cwJzimo1JxPKy1FjA9uZOa+ZXaFafmY0xf9d5nqWRiOzH8guS5i
Ks22Utow6ZeR+1ud7BT+4jovl3idM6glfUcuFA0wGEX8pkh/xQLFVGMvGuDrUNez3gCSYgQraTCb
utKhe8AP7XjqSbLq/OFr1Ot+wP14P3Z5wtXZcqL7X/U7K9jKyIlWKSZ/OJ/cRmUjLecoTnLHiyxW
0kZb8nTY9ZBxUrp8fvNELIawshDNj+rv+R/PU0IOF0U/68DgYjjC4L43iCZAKcz2FRie9D2jP8mF
/ETnRCHMwksNbVe6yWDrq9Mm4lzLs6bVrPwLOje/nU/cYJrEMGjEtcOWlRAnkcwOL3hEbVD7VO2E
XWHySjiEIt85LfDa3T0KXpOs68ThORfToN2MMHBe8WA1Nz3jfX70oF71HNjmmWDPoMxzGODPdxeM
6iJ3e8Qcrtvi/4PA3TNfKtKuRylABa27Hhxjq3f0+BJ6sLLDTjEj7VrQXIDNq0hWQXeproquyI+E
PE6jS0dP8WuDApv9zKQXcHmZgnSR4Xlk1kVvBMmRheDBMIpsJi6kIylDddgZqPfbXcvSKyat8GU/
UIVdPvPzcbWwpRzOqjVkPl+djkK3nMBDJb7J5Sk82Xjl0Vzs9F1tuvRrigBwmxAdtf/xh0MacC7G
/KctUU5a8MZ7s7vLfTbdQLEsSCKOpiXuqn8MHJRzxvCnvz1zueNM6RynxkMBYUqyA7l+8CyeJjF1
dZjDMgJ3SrTX7z7Ky4gosV0T0FE78aqpo8VdICTGXIB2U3XtP9A7A1cV8+n5R2f04ymegqgdw2bt
DE0WJZE4Th3Mq9mCxi64qDqLWPwhVo4FpAWLJJegJIxPjYDjU83NI9rRHjMxBjwJ6bWa3r8sjXF0
o219+r8nHNG4PIh30oIuMaJ5TM8WPgV8KXpX1XC6zpmk9E1pmMRtF/+vpkw3oz12gfQ8jLQIcgbm
sejwOSS4agVyQ6ACOxXVxNP7JJOr5XzbIGPxYYfLtUzsm19a6+0zU9a66vVy6M2tU0pwlbXS8ZGP
bGRLUzT8FCyrtlSs8A7q1aJDnetmy0yZ3ha3HgbMWga9dz0wU1YxFxtQoruciWF+QPFr906aYHvG
HFzfQrXG0602vluC8WBf2NW9sdQ05zeeSIEdni0xgAbwlYWRUVUI4KxMGAvcdvAjMYdWtdz0ND6r
0Tu+8x5oI57tPhspN9M6gXqtk7l50enXtA14ETzX0pL5f1eCH4ChCq4Zt0XvqZZLAu9PNnpwCsoP
yaatdVQfXanhaN1th3qWjg0Zw20Ytx44a3jZYqkXzGpg9T79De2rpK/nX/CyhlfKLrrSskjo/zSH
jrywWCRy8BCRXyINVYZc/ExruGbnQNq1WAKPyRH/9ew6kY+pO7z2z8kWYXsMYGFGuMdVk8u4CYDy
Jhhy9/3iBTVja4G87bDLXNmP6WGE44yUFH2RJyB6Dw3DzOswBm0IynXuqWLEDg2iDVNag4mSMCKl
1xjC9ffZHNoGXNc64wnFaZgWn+dUdrMUpjdHzT/rsov+sbPgzg7AtCSaZRcmUVwW2vmq9GgzEi9d
HoiqaXF1bJiC00cObxBZB2MzTx/Ott+1om00DDssZ+Twq2iz7+UArJkOkaz3viZ1WwCBRbiLkcWy
cyfxYCWJxWDmsOpCYBdkTnZouqngR53ZV/zCW8ME3B7/anh6n16lwBKlxTUH9BmP6YqOP/ckpHk7
Cfb926m0E6Uk1cOiNzspaOB+r82y53nboljc0gJOFxU+zJaMDXkavSXnc52b8pcoI1sE/b9klWVj
W3u8AcDzWQF6XBbzib3BTuLpZUc42vuixZFE9L+lCLa9TAjHbFtC9JcPTn7MoeAL8w2AD+MUg7rn
z3HmhDrFJlye5kL/Vf5xgzZcmv2AsZyd2sqqkFecIP3VwdXKlbDLf8so9V4wUIAuErK4RwDrVDoh
3TotdPiFTF1RQg9eFNE+aOvFpP+qTOAu+zQAeWr1JoGXI0HcLZwuwVXO66Q4J26KsZFDKA3j7BMs
SfctLLIDKckws9FlTmo/wYSB2e+vBHw1ODohP90yGXVt5nIlVo9GAG+oXwKBnNI8l5KCidtykpOO
AzqerY6J+EkGrC0TWOMXTUidUuuKCv0MNd/pajcccoiWc5sRDX03JSsL+pTRfour6cch1E8F0/kc
UEqucCqKvuj6IbCx1IcaPxDCxkwg+KiZXmDvBkht6JY3WI3rT3sKKJu2/vF+Ug02nXs5JBRy0A4Z
+FZKhoKbSd+ZgeMdOJ/mclohVVxatCrL5R9JQ1VNpzpg/15Wbjd6k1ck7ZHfbY81z70Pb8nyA7i1
i/DD5PBtdUkLN3hz5zGXVQ2I07PI7mk3iCCt/wsXS5pxycyC1rLOqy2fp1WHvpiRJ74vM9XcpTAL
aiktmmlt/WE+6pkobcp9xoWK2gEPYcMqjpufv8UM0FKoL7u0XG/90vQRm5g5kWMA5wVflP2Mmi5F
0A88ETHiH2U8qgdJEKtXmJbuVbBkkFpzD+H7oTEhzaBYZs20eka8/LyeXVH2VZ9nvcs+XpPA7NzF
DvHKP0v4gdA4tFrM+CmuW9agqdDZhCjo5A/HFvy5ESZ7CWHXEuOo3rReywHsuUxohCEAgXXT6eF4
ez/DBb3EeCgqEyacE8w23qJzM49ZsZ5WvLY+ijOkOeAjSxDSXqPVL88gyq3vgTH/Kbk9dQ6RqTjb
2iOMKBXUunoo2KYfE9FhSVcZOkcB+0vCv4roh1SDeWuogJR6vCYOShohUj4D7VDzhf2mOFwrrqRz
XvWfIw4z8TBv7UaD6U1HF4UZ3p/bzelwxjoyu0rBf5jGIISgmj19hvYxWhjhrPGgk04BLS5CwHgl
PerpiAH9xNu6NcyPnVc1GkoPlTJ6pUr0OALmdp2/ATH2aqSSwiMRRDTq8AeIEBFckNaB9KvKBJxg
uypwjfOQe4vDwBzjslwMm6ZG4tw6GzpfQCSvhfes+MAi5JRkrXjb9P4RvW4DrjEhbButWCYi7x2X
Np6zidXpEN1uBpsZ1CLBT9YUBVxcAFZItWPEJLIVlaZIbdb3Za5aMXX0w1JdmHhoge9LX6JSF0kJ
k2LtpPWTmAW314uxPa0qHt1Y/ff3oar2zrXttoLeuaQl3MZhnWsq8iJDYoz0K6W8CEj8Q5VD6TI4
lcSo1bmzvXREgCPwhKWB9V0QHwPpqKmD3PIR9KxTRUyHnM8k/yTGRKBUqrIrKfny6jPudEp4RZ0A
DMvQq35jQyCalp8/TFP+dRRU0W1Rj7u7IXJT1YU47QL1o/NYahG7THRnd3bK6dfuFx2sXAARA0Lu
KW95pj4vy3kdJ3bnvyVocj06w5NBAyRvxGZEslVqQh8fA2eh/32vXuRHmKL9A5V+JN8Ejitu2QAo
MhAmibXlDnmMWXhBW1r2p9hIxXx9JgNzvjLLchd9G0f4t2n5jmOSW0W1P6HAvH2yN5A/hvDFEipP
kQm6/20H0bxvtNWS+T7x/h5l99BfuZLJMzAIR2qRA7mn/LOveRp+eSohT2/JvhwugKjDuzMWUcbS
NRwVJSBUja8tdr9kaxLWd5rbTadyc+Dj0nPr7YKGrMf+FYDPkq0U7Re5ZNUzfl5gNDOkwTe1JIxf
xsdKf8bDR7ltPkZgEFra3ae+gPc/Vs5XXBpnSty+frCNkajncTJt9LjIaWOTDsjlDyohgeZPN47V
pIASNOM2PPO8EXOL/LOLLfY625A6vF2MAFk/Mg6KmMvN1J3yRe1nDe4X/jFIprRu5bax7LOncdLW
ME25h6Ay6geFSkLwMGhWiz0QU+CTpBEm3vVUDY1OPK7gPZwe3TSgxg8CmjXf+3p8bZqOqotsswMA
flDt1U4UnEdZZZ07XMq85KndCLnoiBfXmzZ0XJIpIAJ37LZ2o7obhO3esUh1jk27kO9HTHnz1oa0
oZv0ai4vn1OzFiJOQNuHAQ3gIQSZCuT1A8QSt+BUWl5ol9U3pn1Rjpu57tu+SJvT4hWOMz2JR6Xg
gKvM6v53gG3UiWCtzZJLbrQMMGlGskhjA8/Ezsi+6UI6NEe53AXcNnnbEdULQBhWYBB8mE5sDWH/
+/pr72p+cBTHewsJN8VlmXHCxQ1Zl/hkOlMsqbqnEboiQ1Qng2kbnulbOJuk7yqN+H2dx4YP4sce
cdH/JZfeaGUf6uo/W5fTrTtDjTVKKwraVdZY+RkPt1dVaUbtW8MQIMh/cOCq69QU9ufdwtzIG1TZ
Ecyx3171XFZFLWmgAIFbAEOW2zcq/FBPoij078vpRtwG7EYMdDg8trcTNh5cEBLcnZ68f8ipT8TQ
z+Jeh8y2SP3ILa6jrtBDkRkEP2PePA4YJGLluWnXorMYn6vGkD28rgH1U6XpkqfFOCUqxzV1rAkQ
VzVDT8/wm8tqjzIfgpO8Qq7OOmewMd6PGnd1Z8RMG1o5AdM5xxurl45tqpB+R0ef71BWzplo0LO8
5WwFaDkBtri0vDgL+Q0X13RSs35lpZRBPEcBnkEXEHQTu7Ja37kEJePSXjmZHBYnfdT6EmgHdfp2
YLijQWrpucV0AmP5Ljo63TbTytP3GfOufzm2n65U76ih13cUN68v/ILxl9NMBshLRN1BBNEnFX/M
PxdIDc6a+ERD7bluLVDNZScYyIGTnG/+7kwfVY4rJeGxeWmCyEYrEuI66tKeZ+n+P8929sXPo+Mg
TcYAP5y3KgeXIDdDYanPY4+xUi4TT1ro9zmMUtKudzv1F9DnTQqBLPAD9w1EbXlc39zj4h9jlJMM
X0R4uOnbXYhjj7YnRdFafa3NAjcUpI38x/90+9S+AMrSXza/OC6p1eNAWBznRGbMfxBv+787fynt
392VEb7d4kEAxSuKujpbHomvymD4pTnDKuluN84kpAKKBLVk9DZlapgv/fYySJCGHJBOqCUmudJm
6uAJbw2h5HB+rCU3m4Eip4KOJyNqZ4a+NX0eSCLwx/ImZm6Mjo5ICrerZphOGDV6jnP8XC91p00k
cgCVcO/oAJrD1KO+QDwg+AmxVu/GXNOnPQI/3/rUI8e4bJ62pjiPUf+zhT+Hccp9PrOIAKLcEV5f
qUymYCbzwqSRrgeTNnst7JfrpYZi0e8BK0dsv17ZTcfNiDriGYqRAriOuqtP0L/C3f9EeIUWyQGu
x+RAhkNsb7OJ0ayMD4+Jz4vLNfT76zFnEnZZDaap4ElXYgjEBqzy6ewknMHOugw+ktTxMyIx4vV4
PBp++kcXRarbbsTnWVgH41k0xqITCZoiKWbOiEmHeik+Ok3/fsLdE5jeISH2jghCniO32V1lapSR
XdvrYZ8yklQ/KfY9Vq3juzLbPN8Ghn/QRZxvxjEwTEcN9CRmFtm8EnIO2tRRmaJ+QlpoB6J02YwT
YZWFxboCSedAcDU5BYbkxfwaAGATU0i0iDrCNIjkRXlVsiQSah2MRgip2hajyxW0TJOWjCVbJe2l
5CBC1OF9+rrLo9K9pd7ROLoKaeTd8VA0yRVXj5M50mpTYd8lDUldGqkpZOYJM0FMxJX5tAaM3ItH
YtLXKcTFF01XTpVtP1gi7tJvAC4raDKwO6RNV8VNXLucSGeSUN3jmb0/tpIu9zvibkLr0tC2M3R6
axRzDRqjVDZyZdqQvvT4EMMZCkKD+/Hd69/NzL8BuWWn8bA7EQ4ESe6wGkMhPPFPDkjwq/S59vw8
0kxiZGQyzZLD/b6sB20Xp3YpTJrEMGEfcsmwQBfBEwR2HRGDbGFbwywE8K6lTfs0b768CCF234b6
uU0YQyAfTcU9UWTJEWJ4FqgMYbfSFpzzqa63Qpdb7gjAarn8XHdhV2KXF4OIT4k9VnzpoJGsLrcg
15tsMsu+y7ubdWX5dFN7UzM5cO+HtKwaUYosTbA96Cn3JZcxNmWe+lPtfMxGOMug9znyVGR9ZSJ3
Cm3qShvml298VnLHupAmUtFniGWIBJIcNkphGldfEYfBotlUGP6YYJ/Vc2n3LXpOypoHCbz4ZGbA
+Lprbd7N/3b2DxKme5UUxTfT2jTszoQz5mPEyoO/3sKXObIA4QUeJ4EylfDBHKUZusL9UV2wLC2y
lg80HEQYhb7IV03rPoyePAb2tBhvSRYp07VjqbvB05f0g/0se6M+B0zpBT5YcrDq3qs0JT3GqKoG
Mk5hcUxTWYLYe0w40vJpiE/N5KZbn+FNo8Hg6ViQTwrTSRPiHD9aVNEKcPNh2NoTsR6qoBw0mNnz
Z+bRgbduhxH/rchl1K7qVz/M7xL+qagi7K9s/LkLARh2UdDuY6YhT+ze4VsDZ9QEvpKCF2gtOBfx
8Onq/2A4ovcF/EMKS958N1i3xqCm+EVip+AWg4I8FhacaHO0DujIeIl/sJUd3Dm7zGy4nkxn/YhE
dt3MX+pp8N9epmotB7peQ+uYu8uCwsyfEeLXIiU3IqFg3tJa6JcmmN5u7M2J3wuOe/gjfzy6aQ0T
oAZfKz9zWsQvQCkwpFt8D6F42jjyDLO442JjzU+xJ+hbWrhTmKcz6Fg66C1KNblPfpEeKt+5Yi45
0WC5fBru6x0NCEYjnBc2OvVaD4stlriuK7U4B07Pr3AZHcQHLF8F2/Zapbztl2P2J/uTVf0Pu3xz
pQnb7ymr95uTb8b+5wJlg6uGXUITWY4gEQaQugM/YK51i6x02ccdAFyBFhUQAeuF3f3j1x3Fb6HM
A56YSCgsHP5dLyUpvheG5DrgMKXc/4+BamVFVcpqq/PvGVLj2Z5Jgb/4JyirJqRG+rYWwFWOoIPn
/nB7qoIUa0YOzBanehHhx0GQdOWikPWYh/PpHbnCguVUW+Sn42l2w1CppYGq56kK/cIHDqVABs8+
aBgUa2Tw60gR86dIz3/eNhhTFbyUNiDdOOsD7QogGT3ZlVp1HQLeNqj4MyzaZRsmlyvkeTjHhGuQ
RQ8QuOfDFpbyd0aFSj02nClOdN5B+aTZqCN1BdSa9p03VK/qTJntVJVlXj20vl+s2bK8SjtIRsTJ
21UwP7/2hnQ76fLaRij8Enlb3KY2H5rdYAFSM9BD66OWU9/nonFnLPpwzcOJjw8nbsU2qMWaDUeJ
UiUsByqgfQqzhux9k2xPcs75ql6gl+j+sxxmT3fqWal6tb67NWYlt6tDtM3TM0C9tr7rN1VdDmeP
GcJbWnpLPnlI6Q4kmBYduFHsNLHhyK8OyjW5flXvy1NZY/izeJqFQ8c+GJdDg69o7eCId/sum5ua
7sGX0L/BCHWWSh/hY1+6yVuoxGmG3GsMaFqDIkD7yNLES8UyrYZn75oxPoorHNxqZlf4v0o8m6Zv
u9an0T7c+T5pcuZRqSCV1rkTmqwE+EWtZJzEOtrAbNh/1J880Ght20VoHL+N9tSj4/N6/vdTGaqn
Pb+a3jmcR/LAkUQ7Bz1mvIO7zAE9kEeOIugYC0Fj7y5xQXu0Gdv9VtV0HofqM+QOTl5iN62zDvks
3fejD39YlxLJVOUAgL1Mn9upvJBYDpdhtyAaK9F8mZapS63vb6zcBx20i1KEfhNfyVEdRaY8LDDl
22q1LOw2TDhWqVb/UON/OzwImBW3frpYgXLKkLBUcCrQ8rl46xF2LPyX8vxzcovM49wf4F2pUjOK
xeev1yTayjAzET4Q0nqhsuLWKHcfism078LAmBIgEEc5YBq4UdjdT7cIvdwYrGaXl1ehbRnQm5s7
L/LeDW0OqDD34f+9YXkQVeLO+l34IwcnYCiqtYej1vuAdTu+P/9xZfqlr5nWoOc1I4j2Vt6jKtRB
eAzM954fscFhnos5kA1DHEvsGp2/X128gP7zA6Zl04NjcG01kEHb7clZq3QbZOeCztxddCQS0ZYF
wZFooHtIwz/3UsMYjlgnc1vIPlOWlKet7CtXzIubG4SPBxlSzdG6i7RlYk934t3s94HspC2qQVqB
R+hpFcA9mMvgw/pO/GClN3bM3Ar6zmIUVgWmZgqYpCfPGnE9L7vtcslUHt2FEXgN4vI7/hsuesd+
DOZM7YiU/VB0Cw8uxOIdkgkshW0X5MebVcP7/4hpVRpFFnUjmuSJDrAT2f6ehSngMAyaVsdS8/nM
lIjVPgw4XZg589zMZq7Cm2Ridc22y7JvZ5XeizuaxPaRvr9brQ+79Zz/0HrI0KcahbH68GWQDDdJ
tJIOnJx8Y6IWkLewcoDRckK5UhM4SkJMnJkRglRmwG7wE3P1sOtj3vcQgCPJGLHCB6GHQLip6Wex
SF7x84MTIMvQ4nkDa3BYMkEPIUkMcbcwVYofhEf3x6Ylj4V7rlqCK6kSpDtatXhwc4ru8EtqauNm
c4W6jJExcTeagx4bsBuN09UDJZg4SlNuA2SAwd7Jky1uRNj91X3cgWvRJK3ociaW2pbpxfh3y9Ah
bfQgSG4JrwCIZ0a9vp0k0wheTB3hGAN9HEroa/sTmKhcajLMVPfA1WuPrSXPYTOs/ihUlegCgwKj
eqdKBUfQJqQd7UHOZUl5Ry1b34NId+xZ7uipO56mozR7umyifPVWl46SV9JS8fKn33kRT0mIlXuR
GCwzlLrS/xNeW8cWJqkf6eHc59nxF0HY596wHwsBHaudcH3stbVdCFkW4M4/9x5qJc7icwg/4N/w
hpwoEbeIIpcat0/EPxsq+UkUlUfTZEmlm45ggaL7K9UPai8jIaRrw6YRdO1J49JeX35dqVQ3yysR
pJg/PpFTsGkCFOsFfZrYhnsi8GAzgs7T6U/3V6gJZf/JASszXccGF7BF6jlGCy8OlMExzVvFtKGp
HerrqECok0Q/6JNHXBnAIKIETvEbKmOmr7hAugTOjteSotjA1oQlDVHy5iGuo4mWPaChp7gV1zer
FEN/bZr6xoYAfWmLuFb6y3RGZDRbXxQBIC801zGOaW/9Iflu3f6lvSB9uJb2s1glTn9S1k7iNtcI
qQl02VMcH7F9j1wkfqxiloR25dBxrwDcmm19uKZypq52IYKj37638IyAULyCvng4UwuUAO5HZEgI
5R95GisheFoQTAU/grwDc0XkuBasVAQ0hPNOONaiFj4A123/nFs2JSmCAZUeObimceP6a2Vh2cHp
KrMyQxBeiDQiNojG/mN9Uq3xnRdZai3eORLCQw1kAMnuT6gyy8VN/8VOCi/U7hXCXr67rtrh6z/C
RdrGqkQ394qmsGLgre2D6jGCMYXg2lfRVet73j5RMOfj5lTW79UPbEpLO9kacyaUt2eecAwOG0mj
vSUr5LEEMjS4zQwAe4A5Wfk5/Hi/IGEYwvwq20zDbkEtJDJciqk7g7B20BE8vHAOKelSJFNO9Z2T
Ow9GrKMeHH72wIuCfF0DF1iJIL/hL6+Q8an1m4m4qX07XlSsvGBI9laScY3p2iB7/fxTm9zAPvc1
RyJ7LRFjJyrknNR87dwOnB7IO2deOqFohKCIh4FA8+4SF35m1be13koPA/RcjZCfLKjH421eYH5S
ZV2UPCmxTZkPZmTqSJpDGyEdMLtIWCKWQlmI5idGrf2q5EOwAxBIbYMu4v+RBDonWXNxIVmuIWxZ
FMahPGwPI0FZ8eguoKg5yJbOCdUyuJGi7mEcrdUGiYlpOYM8aD6TarKm1XivvGtVyvCajYlCHrYm
2OoqF7VB+GaVmCWK7Utbp22Vm40syxPwVDoZGPs4sKEpR4xqTo5JScOmKSl1IE2gErmgzUOMSN1v
MB1wj1hq13ZjGoAvhDPEfufrEtVcdl9VKK7sx+ZQRcTPP81YnGiKbSre3QfcGr7FlTbGaWEuR4dY
wC34/+CiY4Bf3vidy8EDyHcSzfElvyzl53QmpT0PPN86/ZvHN1nxYtJQZnRFZkLcBuetGa0lLqhv
zCaBK7p7hNqY7/Yr3K9EF9S0gDjTbiki1z/MsgOGuo4vIzkM8KXtNc01/EPqm2PnIo9QkqSFhMjB
laGp87oVC9Ubt/VdEIxk6XpuBXZ/SxC9SPs+RA+ILARVO9U7v7Tm94pbsaiVEErXoKV+GaeKdCEn
4qV2vyYVp9fPi8mi30eii+c0ThMxMRVZ5wunGMU4kmWTRIQ/tQikHVNwHQErVnN2IZ7BU58Z9COQ
x1TIRkwh9cMMWKEhCVryaoYrfuL/EsciH8uyTUhK5zoVBCf08CT8cIOCeFr1c0qkBnjPntAJ7/Dv
NwsVhyxWzxtApJFM2VkjBMIvV/+UqT0dkz+xxz3bDiSM37tl6I0G32/CBd8MjQ2PQBfuwS2VnYm0
3KwftJs30DOQcC66bkm/w9cHbb0ltl1Rh+BcGYan1A4o0QjYCojdKI8PMhsPEZiwCVpGVl3qE3XK
MpRsn0lAUX5E4R8Pr6DSwTQQD9CbiwTpWlI3MiBPLIRriepJl12T6s5iG/+g0bKSTGWIzcRDOgoh
I/sa92UvR4a1kuYvpVef2ZzEpZONZZa7ysz+I3iPTUsNeqFe2oaH0TEGfS7LqOmUuPYFh8XBOXYy
kib6b6PpuSCcTq4f8h4Fa68c3zsB+bX5Y2oDX3T/CUPbB0P3HpKPx9to0sXHDuO7u6t7SC/tdD9S
PP7q0713vCJax5RcYZdAgTVidQsP3yNBPa7eGqv1B+Z5RkDVd2lbpH7QQbK9v+Hw/R6XKtlQJiFW
yNTIjPEbvt6v1xzvdlS6zyLyqqq9yeI3ewHRH++KBP9EJFqVBNAaCBlyiTfXABr3yxbZwtu6xD2e
m8TQsrHpRhOA5Iof2Hc62Xe2g4A+3z6XwOW6B2SmSwoDMB2OPwGJMD6n49QnObOMv+EMjBT4PM+W
Z3CN7tomVxx19yjhPX/+ijC4epqxXn4mcyHNOBUBymcGxbMOq7mv5wfkNhGggoZ3x4pxz++AtwEZ
y4A3xMtiVT2Rzn4yMmdx80gErnbJMcG/EGF2GznAl6V8VTR5oiOKb+gEofpWxSKE4PaEYqlp4kAE
8zlZ0wS5jAATB2B75pUHjd6QgvscmQ2Nq6/eeeMlYctjVU2T/kiP62Fs64R60WfvPc6yhHCMFMzT
185NxI9wwE9p0Rilqg8+1vLWF9ZGDII51h7fkxw+33m9DwpS+QhNh109TlKgS7mF3srBPQY94cWM
L9C8q97kAAe55KLb/j5+OCn7e0Q7I9oyImCNXGX5qnEuCooSwqoUqOpguAq1loFBiJLC7kwjsg7d
yFKFybkRKzaTmxRgbdyItM5lOtH1dDFXVOO2ZC5ZWEa+X0wSr5Xuri3tqIswThe3YDb+nzvnGRtE
2yL8Mb7s/UwWhoWW3CKIYyH7byz8mA2H+Tuvw9PIS5MjgoUQq/VzqbzXF3N9rBUjX1MB3hxIMcR3
7Th53m8lwJn+JGAOoLUmAtzXru7lgcOsFhwtkeaZ+5ZDxt6dSvdRAikPwe4DP3fl7/8z47XUEUu0
NDSoyHITxHAD1fKjh4coMFmW2QOZbktQIKEpmzIjW/4tgmXKvqlJnPELHLqALSMYcrxfXhDisdfk
8E/EQx0FEJGQWSClXLnQXJqrYUsyP4fXlJlc2VPWGAtPlgYXB/exQeHjj6lQy8xMzVKRUxY8sKte
WZiPrKQZLsBNr/uH+uXs02PCVJUobdnhkH2e0LzYylhpbrcjVeoXkinhhhMxpO7ZMNwN3TJPBqNH
lTYPrU6dFYpPnorY92uzps6B2QZGCQuia4GRHzUY81dztKzaT+I8/1OJPfwbvySNjRxt2kJt+wBX
yI6sh7/Dni1OBRf9q5RTNy5/6Lx28Rra32s7pV7MrMid8UCts4OrsJcNoZtfWw26xd51Y/DtFwc0
SRC9BGowBug7rVryZ40sJieZpCrTLz5uhoJuJntcXL+MBwQZ6odew1Zr6o+Uke+pu3Zv0RcNMF8x
NmzFAVODMSqybc66q2xnvc1ozzjll7AX1YaQmKY8K2pXGQleiXnTSCn/xzcjRNUCqiiJocS4tfhd
bgVN7zX+kycLt5yognqdO0UJRYuQ/DctSWZsMK5/RGZiAVFnPTptSNxZ8uKoenusWoc8RLdEyVJ+
21pkoqTZw8867whwFkv3wkCdzk4ynOaKoxLNqIddHizFw9rMkFNRcRJIPzZixMfW520X/NbcJC/l
sZZ6ykN1r3kiZlNuTCoahXQ+BqO3ogH7fRqD6eIWzwrwU3PWn3G9h06Y+YM8ApcxYamqaMaeKEWl
cjjRMdTKsV+wwi8swoS03+qe766HT789eGybHRSKlLWZLZ0dWObn/eyuRUKjIwFjLWLUVY/+Q/Uy
TWKLm4id6gY84YEP8q8gfXIohJYL7n9MGVufQPRjczn2c9BFD7jACq489takeVh3FFqoW2/xWRBd
cBtqDcCNGXoI06w7rA0PnXfWXHDpAhR1TXFvku1poePIKqrX8UGr1sfUFcLO7OE6oospFEQFDGB0
EjH2qXxHHJJbmq85enZAmKpSXpnuO4zr5v72IwUmcwz+FReDy1TreZrvbS9TItiDrTMGqyyDnogS
XspNKwVDeoyNPHHoY6oy52CAn1fw6Y14gfVeVZb0t0BY2eI+UI/QkB0gxyz+dBJ37pMExWLgjSWN
CPuDCEmQXmrex58foorTfjxDcoPIPMWuSLtXSInFZi+tuFd/9PYpPjaDBiLrD5N8xeBExIguFunm
QQrP/hy5fh14zGh9INUJ/ARmlSuU5JEA7D7kih4EC1QiVG5HCzzrK6Q5Q1rGcetlk6GZmp3i/qxK
kIwMM2EwKGzrrxzXiMtRk1sT2b9yNxXUU2d7/ftabpsnYGqJwgurhKuRU0+b98O43Sq8KOPU50vs
8OTaOgQDxa/Wj3yB60B/OTTydSKhLwUJSfq2mtovJ3TdmeERhPmHizRUNe5aBnJyGVsm3tDhDzvY
hL0yf34xZzDTUK5bakkVwcdt1kv+fxx7dhmBe5S4Fo44M/vI+Tl4rnGhpHBC+Pxqa1jB1o2at5eB
ettKXoKkGfqzVBcci7A6rK8z8TYDwmEncibG/SqEuJvYa3/01+5YTZyybQe3vyfK+sKozA7nh+6Y
3NN/YMN/uuGnqYlEf83GwKlX2TgoEEuxCYj2RcJVb1m7fduMTch2NiIxWm8PO7l3ccs+e1qZMb4e
fdr9dspsdtK8c67nHzy0M3mZqcU+jymw1dIFRnY5dnlicRxMKNSC2Ad2kMFxZahAoElp87cFxLxB
Ks56yYnOCH0rgFuRjAklgVDoFwiH2sCmgy9q8IKjHsFJYSLG4G3x6qZvZHfklFJXawg/EPo6w3LV
6nHrn02Kwws5+Euq5XE5Lgegm73HGOe011EUuAid6kg/90lQNftxn0clfK5Vm9EyzK29d2ZKVgV7
9UsiR86fusKMVYom+xmX7vQApRQmodPgkmOsBbg4rXcVT7+6rvDPdNJdPtEMNQPLwdnVacrQ6l00
lHjSePG6BZXp5c8zMnU5bqwjhTHtKEUk/a1LBD3+g0g5YoJVeel46BG+biUrRXjTY2zp1Aq3+Cnc
wjEMJxA+aCgT8SQ/V71aPyObgiUh1Xd9he/cl6KLUOXO83RnYG5xvx2B/JiDehaIgj5qngCLQuOs
FPOCpN9TOjysZ9TdZ8cAPxSRp8q03TFlHPPr5c9uPqDERi8CAJC1W6bq+sUj/c7W0xX98zH+/q3c
EXaqqoeCNy4HL+sSZWhooeVlUtLwo7Tj7qjrQOfBf9xvr19zPC0nsoeuL3bR3pOWh1/ABvxTZRix
rQRFSZzHXna7xV1AcxztkYxE4CX8jny3cCFgLlIcPS6LXgAFkZNvENjDjvB409ksC599gnTzH/Xf
Bt2U8rJRCg2AE4weRzBUOfq2cFEN0BivvtMlXJeT9Pyu9/8+a0+l94eftI5rF3y97RwRQr+1nGCM
Yxr2yY+3EpkZaPisKbMHPQgbsuc3UYbjiPRRZ5ob1DjGYkHl2ktGpP0wlalKb5IF1lDRfv49JiVs
SFwIt8XQE9pfcBfdvpk+ksXz0/j8pek1/i8dnvK95m4/H683ACIkW4o9q3IiVaI6uTtdJI7aVTvr
P6myDT2pABfbStmmtmzgSCrcZ8jcxwM+1WeCK6WsqxWtDsZcZRHQY+MBADJEhuE/2Szu0wG1pX7s
pxyKP5Mug4Xys1/7nj7mM0rUxwwigXqUSPkTdh0jqEZGDC9UpN5vPuDEMw8fNaGqfpc7S9+7rUfm
a3JqQZUfPs1SW4A2Jxb458L1LRu0ps24QHP5rwGl25fRR+U7mzP5LOOq2QqierhGR3S2NNLbohVn
D8OdEY3/MQ2BaY4GmAIX55g2GQkCqbzseh0+dde0e5AMOK+HvH6ryVaMTrKitQnddlasXKOy4GxK
SGT0ngMuCBEFEM3ELo8s+qdEhViaYZOfzweJbPwegt+0y5EJC+bQJCwRSvakibUQideICAF/ua/B
8ECiFgYg2MW/eiCspZ5tStSI8X74nA9l1eiPzDVpoHF200qoeivk8nlmcs58Df/jQd/39hDwUKRC
W8CNb9EJAneyYC9VY7uvYnVD20V0I/5/hUJnnHwIdD2IDhP30JW5Det0qFxpNj85gvGVLVb8V9C6
7AKVw5QyPQ5WSnJQ6YfMEuudY/acF4lxaVwXYhtHaWDAmF64PINzdHRLq+YmfxKj0C8oQhzkeJ4U
8wKpqrSaiM3zhq10x2Et6JIFDLvWlO+CKSfSz4dsAXuNcoUyGEWEuIHf28WO8bVNfO4pxofxS4b9
0wAmEXGwYz30RlOh/hT3jsV9yzZzjCuE6aKBzHwqNUlrpbAFQl+t4f19+3cAo/4ARJXwdp7L+GBI
qprHkJzxcKgSL2ofhLwRYDvMiMxw3EZ4YD1vKRKPejiyzemVnRF9+qeR0976gjZTymbcwBdE0gy2
ATHRP6ChmGoBR6Sb4fRdCD46nhX9adzQl7aKscFkbVbp55Zi3iTTVVbi5iy9aNWz84vzZVmbKCBl
trXSzRF09FvrT2azjOccy5Pp7YN/GhEz+fogBK5mYBUcohslr8kWDVzRDtkTckxtiOutRuSJfSGs
ZbWa5NhPCc+Oy674e40qkMwelRU1ouI+NgM8ZZwnQQsdi12RhgPK+LaKNSSbchejJsUL6QE08pw8
5fI+T6kkdADkKWHKNoimyeVBiDkcSs+kN+izUvj90hV3nuX61CYylwc/CyDeSxz9ITvV9vQQ1Jzv
5SGrrWHjx78D83w/nR0jMTGlXtfw4eaQNZ4FhvDz7sGNlinAXUhEq6leGTo1bSO9KdaP5Pa9flda
COfkbGaDXrWEk+JyABy2m/Dl/XKrZ+VUQ5YGgcUs8uItm/0A7KJaj4mFrT79BDiVsMRu7dQRmbaX
xJH6i11VvPWsJ78mDXHwW2/vNCjMoS6hk5c/KdmbLX5xr9YkhPMN8ouYW924A+gvPdT1/KOMSrT2
7Sk5WYIEb5gmGyfieQpw3Y8dblrKQhigikO4VncQyg1RZHg4EJ82LGpEZqaaY+SLJdWlz+3AgIJw
Kiz1jKEkVodIaYGMXzMeGQ/0WvsdefI4AuY3Zu8GQE7w7rarSTVtbgZZi+GqmOmSQUW45NLiOmBJ
uXClutyWtaPZI8zL0ZgO4V+nwqFkcUtEmeFQjD5cpuo8eshMMo2jxdAPRSnGwJkFW0S4BH4oOMjV
BIrlkoe2MMFw5Fsk3LRujzZWySMRo7GasHC/J+Mynhok1bWlmzM6VG+/Qh0/1gOTe2NQzv6VR2Em
F4yvPb1dxhTGplTShSga67XRsAbalKBXyGC1lJ35XogXtxlDHgTbZ2Vs8+b6FSI4hqSVTDpaF+TY
fcgTVe8mJibHLgK+iCqobrnfjTSnlXD8ptfjYbs2ZtCif2JxXP8j4jHciyY3BCTfG3g0xK912IFE
vWapfR9mn21TvtKcahsu7ZeIATX7PGWP/CLsuVmdrJkT6NetxRcU5VujjjFJJ1KArhU2J6/I3+AY
ntd2M/Saq6qAKd2Fos74qb80lRrz3HeikZChugSs47GQflbCFy8XsZuQGue2DcD1AWv3o4G1Xciu
5ylJggsC2lwAd5hmV8fM3hBJTQMVcB98qv0S+g/oFSSx2Y2Hw9+AaJhMzvWL9T6hBPK7RNCcvxJZ
G0E57XvA69x50OgtSpKDOUmmXCusKvyjLbKmWoCTPlyZB89eLs5NuALsdeJPtqNwFuDG4n2Folt/
hyBQz4/oJ0f3rsfJRIBQ8CEW1kx6fh8LgBHFEi6XJbBOLNWjoaDMl634r4XuJHqTTHzhAY7uZcDu
xcfInC4U0iS90JrPGiGJc0gMst1HHx75fqNpQyB9hBy9ejWqB6K6JaPws9crPbwVySLZLS3D0V8n
TmBA+pZM9yIkshbOVfZSb3j3SUX2ryP+rrGpXYEnY94MsJob+IJxHLTcbfmeM5yOzYcjSYiIEAPu
/nhANEusP0EwgGdPA8Eq1QwhY9/3oRDxNFMhkTublX46ll3jeBlIzcSrD1S/pa9qkRbJ5bnQqptr
VEjdyp0Mx/DlemgTYjz6wwUR7hHeGOgZeXUguv1VG67CfGTh+ZrA/1WwdsUswehOuhyo8+psJ24w
YqSn4Coag7UO0OlC6CRy3ZeliHly0uY7HItfo/dUp3+9QMVeYS+WmvS0zLczNPp3IOJGjf/69nic
SDwPOoCOjjx7yfNc0AdHjoFiGSeaJjL8i52d2r7nv/euUU8NeqHRG/tvFWCT8960rv4JuObZuvvn
guy5Gdsj+HszUazu2W3sGKckquu+CN3tMniHAHLoRx8ryKKZz9G0AgyldlW0mY0/FUnvCYvtjdI5
qi357xEBBzE2OYAfBroqNwxU0Yre07fyBtAM4VW+7CmZTMIGlYKEeRBe9atoJwfBN/3lICGxV9kB
OCbYLwlr9aZpVcfeFO6Q8iELNkLwJQFKa8VfS7nsVlsLje6lWH/jjG7jdou3NAXcfPJvzYPJStUP
Y2QcfxdcmH3yu66VPU2oN89dNwlPIV1ktrc8YNuHqU66jNkWyTIMy8S7/8/3lAqXr/NGGTSGQ7gC
m4/IsrtoHDeuJ6/y4Eu/GeD49EVDeIxZvtYN2T2/QU4DWBl1Hvpq2Da47tpxbtle/zfO0rdXUV5s
+GBEWGg7x46heVsQbq5JpLTFRzo2L57AIbz0ZcaXDGAvr0KXvBPKtojqBcGY/pqeiA9fheqBUF0B
F8OORRhHRItA6UKuMXeyMg84V22fT/t59JYr/GWINteIZlCMiLyaY2JFRj1oECOKpuIcU6C/B/6Q
V75gAd4dchWSYP0U0oJpYlo/hhgdEdZEH0ecQn4sAblN3rgwGBZc3UGpj++b+SJC00nMeHtZ4HNP
CFTHPmY7NGAGFk+qHc3+skuSPuvr+0W45NJNu4kicI1X0DZUFAY5QPP3wZ7aGazjxICafR5OhdTz
0Wzp2fdtCBLmxIUTdeZ46YhsP+ZMTsaKo9bVLKsDomIiFoYQTaSbleL/yqqSus+/GT7YdgCpaCdr
Y9EdF7ENE7847Mw9H6hNq5SbrOMtmQSxQIE4VX13rVyvmBMCadsuYPcCN8emJ9vu3a0SxcnlVW3Y
L67vFfDvcoAQ/KC1Q5q2c3zIdPzDYWGGFgIIdXh7hQfLACVh4NvvnvQD35Q4QV0UOka0UeDmZigl
vWUhPNErPisNrZn98MBAD/PXKd3e90uYOgKwqOHT52fozHzbuAIAuco6I6OhcaaoJ4ubls33yasP
JULN5HHXdYaMVepJVZAiybTMA5i8oqoU7I5ML51giECPxczyK9Ri+3xsTZPmLQKc4m6sM9x73rvA
JSdYuvLZktQP7dpjiVuB1eq6SzrLMMsILD+MaSvaQnLEQhMx+M1sC0UmyoXystN9D9AA6L559wpB
sBo6I0xm0pSTUkS+UH3C0f5B1EjGhbzra8W0bRWJDHwzD9i48v+nv3DFKATwuG8MxG9SW+D4TxXA
XCw+JLBNZje9fY19BeTC/VkCLRV44kg8z+BWa0j5Fua5Iu11qPtRmpVXo0qOJZzNPpZOTcFZ6Dgv
jyIcfJDDHmsCPVBKvZtSnINPJ/uSQHMp+c0SM2JKjRnuqqvSgYyzSFkG+jbiv6JAWRc7zlogGeD1
9WecsCo1KUNCHmrLyYg3bO1QPuNeZsECPOY5kpfS8TR7klcfvuN+bbyc6QjpIx22po6xBMJpD+i/
AaBHpPJwTyzVv0GeGVRX2QuT0ZE0DxPuBKlAPO29BpVMdtVzZodlh2WZ171dD90vQMoAf6gZ317Y
cZWv80DnKiZoYrkprZhvBRrw+nFFhIU8/r007DFMj34HrVr0Fidqx6J6VZQjdyUqegrwkZZL0xd6
kUVA/HSOR4x6iO7PVnOSbGqfjefMoFvG0VYq4iWSbe2lU2Ha9vE+iB0ZiZ12uHBVzydpV6H+9o1q
ohq9M3CuG8BbFeiqni7t3s1KjVBH9f/WhcaFedYzSMZekUX7YufH/R0QrMTAUJiap8Pkflym/WJ3
MIsscY9xwJV5qHmLapgDCTkpSdlENGgm57s8iqcmco3N0n7ffbkPNcLg20u92bsS2ZqShwvFgrV1
BnX7OF2ezlaZLSM+/O4oocNUdfGl1+YOonVk4JBjVbNkPvMW5nACCFmzFX5Km+bXtrR12YUPUMAD
GvPxQ77ghS22D/nH/cz6ofws3lAQZ9e3TeGNRUxh4//95plmbHjzHvQa4uNkqgJmTf5E/rgFjGnn
oGf058PaUT273r+eZpYRtiohgdRRyRXcAhhdba039FaKuLLzXnAAEp6dvEExbnZShrFWbs8Rhhfj
8dKB3n5wCVSpmsTCh0leWQ1nCYG8ljgF6h/Hy0ufLJPfawjxiH23eIxRfkc4tZxdZ2QmCaj2DdSz
XK0K8R8kcMaO5XnPvWCy8km4G5UWtAzHK6kXb//np0pYMp4OY6WyqkdSKe+tSfVzu5NA54dkwfKn
OqvCJRlN1t0zorz3CVjuwVSbjYaNczJtB3DU9VgdL8DRArCTf5irDiu7mB5n0vkcEH1kMJ6FusYE
HfW+SKX3aGglJkEUg5DU97Ls0DKmbOiYmrrKQeth6J9AGppysrsFSZXFosw2zh6jtuSVnkf3BoVk
6SZYevCQ6efYBAyLc5Ds3ILcOGlm+OcUKhTyJlAqxG/lBkCjBF3cm8Po5JS8dzzgjqAvPDFRZIe0
aURSmdhrq3KQoX3UbbEwGWOxehVW+YoDu1fPSmXwKnPYwMaGSixtsGaEhBM1up1B1vnZX0kAX2Tc
ZfSpeBi99cRo3I32UcUmD5ZvGU8ob1IdAI/gHNdSR7GXPC4J22DwZ2/m+90q3lSJ8O04rtJk41YS
JbnILdjfeXLF+vDNIOZnE5uAHGjKSUMxI45UPQ15D/9ilJV0WG9b0+fFP9P6Zq8gED2giMdOvfAM
0d4XUoaRMT+/fps3LOUNnwXyDnYkIMPJZG1zTlgZqB5PQfqfy5WYESgCnAJIW13V/ZSgXxZh4k1U
7XrUXZiB4/CmLXVAnTTuDfP3s0oDcdxcCijKzJdy6gai2RmYwxH1UyWhGY5aGoksT0phFy2cNyxS
Gir4m9lC9wYp45UbDjUAcdinLtFBQKYUdZ0qXyZnI8mhj4e4L5d7E3g3npqdp4CG1iQbsOp0T2Ot
26QSv0UewrE6sFJg5nExE7AqBRsMZJkIIM5x2oBBkiTr1NumC4N8dAwMXrMioOcO9iy6R8OE1veN
TVSxr7GVEllWsykEQpCvb+nAVMClMBQC+UhrnPo9j/SXB1sCLowwKmgUKaScLBjMZotHuPFtBlKN
1aF3+QzB3LHehWCtHK9rHycPJkQHNY3yvwHB5ra3JxunGmZ+5Ozsc/3lxsFMEttVoLmFBWc9FRun
pDRhyPak1MxsXf4N5PYxcMBGDqCcbR/Ndgkx2Yab3dQaBOYaCph9c91OKDKOP6+/JqqnJIjrp56L
6h1ZTVnoxeDxxN1yTEKPU5ZSWVhNjoVh1Z99n0SUbUwYKCpc0sJdeSXjgMwU1gstkxc51/EdYELu
VUwCor1nGhf7OWqKG7LupfkLI7pvmpwekZNzCHizVGEUM7n7SJfrOwitb+/ya99GaLbY6sG75O5C
61TLTJpi5fKL7IUmz3hVEvtf0ILmMpfyovz1lnoFtIGJg+fRjs+E+bw4Jkj4BVX9gppIY6NGFN9k
JnzCYVkq2nONzVbOJev6tRJygJyPOQuImJKzFifc0PpISUfG/CZcxwwm3+mgyWDlIg/nzk/uGzJ7
4F4xF2ftC93wthYX9oaauXANWl0o/UblKl61PkX7wtBKa/WSx3AODTIWjVzRs3/jLTS+0cMCQbrz
KobOaxNbQH8glf7vkZGtZV+gIpZb5trawV4oH1aNJXL0hD+CUvk/HcpSzUykFVvby7GZBcuAXEck
/e8mGBiuvGXEy73JlW0uhhGvADjD+ET7sjaLaP965akW24tg7EbbsygMJVvQOm8EoynsgnUzYDcs
eWMjPZJK2tkscDgp/09tX2pPGDH2hlsb7IoFPZAYT6TyUhdCK/cUXvO8sYyECqOlNTgmFmudDZg1
ZdcwAt22aqG2NScHX0/pAlGJjL1uUvTfcnFW1BZwl9ymQJroGlTIEvh/dNidzyI+hGo79X+1t52O
wj2QgnCCEmAzDIjR0OJSLajEWIve/pEqatBWogRW4ms2zXr6FDzAg+2VxrJqslPCS/0dh6ishPhK
JynIQVqGS5UugGWXGPV+hFNT0eoJgZdKfqRsrYQPXJMnNkaeZ7WFXMGltWvWy2iX0ukRrdOVVN2D
CpekX6xIkXJ9U0xaudmPphWAFr3yUmrwDUUkARZF4hE2VbV6wp8WGoVjJV9Zenc5IWmkNm9/cTw7
HO+sAyu7uX6qx63ytVNmB+W8snHdgjC/K51E2PoqtWMrli+YwirWIIuJYHElFD5NiDAe+2DfTbN3
l4RunNM5xmPOArnvoOZpb+ufkhU1zMRQIgbgX7ilr2NQAsVw84kJdi/aReZRyUVBZgFH6gA5qhpt
qHqxThkFH1A+iEDmNlyRrj37JBMejcs8PQ6MCGBRdNGs2jYtpFenU0pzmmOI5TwqR7x4f6SMEmsD
n3fLGPaHgNnQ9icjGVHpKnCQw01KHJsTZx3ZYzF9waD3i9AZuWLgMduxDiGXkXqOIytlapBjnBNB
o0SvJTw+5/4Nog/jp5C1iS8GYjrLKSXLUiCCt9iPWWT9L7YrpnmkmqJACICUosqYlROO2ZWKoDsX
T/AW8OyU+IuhPNTYUVLUCB+LPMuNqu8i3e53c40x4pzoKTp9w6/7+Lypn5LhCR8SUtanrM0AaPXA
mTNaWL12Dgb4r9OilDLzEyapL+4IMAOMNO+wi8yjymdWZ8E/CxGPiao/rmBdgFCCwtT4zQpjkxyi
m/2T05u2maW5+tO2N5EmjM9T681md4H27MzXZ8ICr4CH6FO31X0JbneoN0Hu///s9rWEVQLgWGbd
tZ8st4EdNT5g2a33BkkLTJ2rCzLVka4mXQRA57CLXiX4G4ZZ3+WaAaz5HUXLMQI7KHNbH5tWf04A
uabS14kX44hLPMrGlrb5vbyxSQ2AR+Jf85iBnCDxNR6Noodh2FSzD+H2EslCoIVfVQKwHPbD6ysR
FhPyEF9AvxMEXyv0y1okx8VAA/Ok09q3kjQmdtTzGRnMu41UwhVfXXMjKRiuOBI8oPBgavt/Ycd9
6N/9p/miqMChsYqQC07gvJvokxTj6NyhJlZQb9yK+OxfL9FsY6Qg/uuwF28XlI5y2uwDvirK6aQ7
U74qH9mCnKHaOboWP6YS9faXzDmLaeemccR6Gx57xOY4JQ6Wp/TqxbNxMiuyL833u2fmQGwosS/n
bBn0flABSaFj1agNj3JP+3aXqv3BLWRCF/ZeUXCCqYjG/yULUJ3YKg7yRferAr96LK5P1L8mPgfh
xDSNrX1qUiysdG/Yh/Gc+675bucnv4gWlJDgSFD5iAz1yt3zPdxD5ieWecHQIOEns2DjQLncbdoo
fBvYM2MFa9hwzkibwsgQP46C8XHAJ2XWYhqHpqmpUa1OnW001TBBCJXCe2WF27u8VueH9pPF+qLX
ieRZB7qVVdqCxlgVJUhWyscwnenDu0gl1rFuW4p8LyluwXgRoX6Yp3We2RsVCss93D4KiSyK446N
rMtlEOvQQklpBhgSao5+v90aS9LFpnMIBrs0crPIEGzOgZwVsixoX/ImDLqyawyu2CKBjw90mADF
jnuUrDIRYd+KGBLzpULAkaW1VxjZO/A6sl2UyigxC+hjZjjjYM97QEVhnvDoFGmWBzedrMj03d0q
BxUPu3mDgnmJ2zlsdCllHAYk3yte1fhB5fde6Km7JYSBqSF0nLYdeiObg41hQdSa4VFuvGSfWlAM
f5ybG0WzvBm/hMWpKkfcR5alpCH6epGSK1ZyUwGZCq5dhs/Su8vstWtbeMHInBomp3naJy/JJaA0
aqPdjG7MIFaC7cDXUAGIyp5TydT/NtjoIbz+XJUGruO/3tsPrblo6nzezGjTPX7TYSKs0hW3OjGY
OHg7smxQAB0rg2UTt7Gx/2v+kn8wZEOMYMFemt0hGPZjYybkMLYWr0aEzH/cK53EUKHS2R5Vfehn
iDgC7flL1wHfWVI88m5mjjoksTIof7bDn5/0u8UHlUOTLepJ0WLNqK7XfcrhTRrk3hPp92jbtePo
T8htNhHmVW1+OIXLx/Yr+kfmIC4Y6gBsr95Mj3ubOFGmt93UBZq9APeRmAFZzCGCMO21qhKVgAFP
BdU1WKpOZz/Vo8Err3PEFXJ8RJ4ch2RON5r4g9zBGXTgtPljd/Mdvvwqo4iV5t0895INNHWtBa4T
K3YIMWiuirIVF6t1TKXIgUIQ6EouAzgekMkk9eT9kt46n/KzRvCYTFJgrHvJV+oWXJw5mnis6zW0
b7wQvorVunFw5biqzzdCYQ8c1nji6SBzwRp49EdTUm4Cwf5h8JBOoh1v+FooxKsUxl0LTuefZSDD
HCque8TFkHZPQSa8Nqg+/2ta0+qD7dC27C3OK2HmxhNE+Um7f9w0UEfQYd/LS8oAWSZb4Cqfs+Ti
ZoW5jR0ZSHoT7IpfG5ZtDn9Ve28qSu3eAOPNmbKhbSpq4ws0uyqEdsHTgYZPZClnL+EBek99Fap6
7A3HkJ2J4fYfFtce9K+XW7OWsn0PE3bLOr9gZHlyYsqbhXgbkGauGEvpLp6LGL3UVHldGOR38RAX
omUJ8+7jUl1lXXPuGsEsVIGS2EfDsafxg7RRSJ2x2ZfniYWXOwjw+CjqRMcbr+vJlx8+6m3TIw2J
FKS0t9xyb8X/csWhmQ764C9epFNhNAEX5NgouhvbzM65lk5T+I2ZB1F2uA8SF9VWLw5qKwF/wOsG
GJcEZ7TJitf2AxUC0xos62uJt1d2KfVKQlbmvu4COxytZR9EE3V5gi2OMj+N8g3ylYALUR4EVRYr
jgQtuNgYP+JzNpLago6gbAdfBi2J4ogdgQRj5AxLxLtc3XN8j5y03cAZE7hOrWfUujDaOkh6IeAb
Gp8NcUg2gZY16Cr26zMSjb8/OsW1cdYuvCyVOeh58u6SAlkoyR4/BKlRwTQJ+mszk/GPwCgqunbk
2APBEGUvPlJyzrtLm9pHezkku8MGrANGHlt93UAvQJkWmD3Z5FTJfiwhoCvf2jE2nXPrqPGVCblx
smglkbrr2HLHqVMyYxf3QBElvUBRIrmXaB3+GzFXjqPrN8iUZmZ/EVNErIE7H5vnyFEGZo2nS0zP
rOjnHZTZbUL+VVFoaWT3X7/aI4HekAeGFb19CuRswYx0rsRlhyGAAQkjtvUQWkiGQwYaia4LBMTt
xZ/Q2ZEnFILXT21Qsig732g/td1hhhNUk19yWpAP/oL8Z8c5Im1PtPtJvBXZcE6rw5CAxP9Tgizf
hjwDTtF5NbWQCWm+dKkgM3Li5iY0BCOWP+fTdgPq2rZxYSLFZ6y5hS0LlZ4f33DBC+MTvSaW9ncL
6II4C/RdwW6oBWt71sVJpYz//b6Zkp4+UibRhCqAOd/uIb9K/ks/oclPopwgb99vLpFbNUVnTbj7
81XZ0HBXyxl4QvC7IyM1chHgH1f4+C1agmhrsGFtmpLDQkgJoJRsQXieesKSfsFnTNg+cJFFH1WV
AOOgCD4gcvCSCVLmgURID5xI5h+p+kUXYqH6Gj4li/iFtZy3OzVJxGv+GDnbvb8zylMhyhIvVc04
fduWS6Po/d/Fv6vKeLGnVjvhQHax8fNYKLsQvt3vhz3bFsl5d1fekTxiN+cg03oR13J9vgC9L72d
7c41Yklb9JU/+dW6hu7fb9pNmmM2j78ImONzOVLZude0rLXEh4HYruW9ZRd+YApYdY9oK97uXlLM
Miqb+GgjvhtYEMsuGYYDr37txTgiKlYYQ+zdQZ0feOqiigzL2sL7IW4eY+hAJJhH7hyG6zNbinnZ
hnWDy9smir/R/xHLh1NafFe8WWbdolY4RIlzHXbAoJCFPJ8RhJRup6p+B824I7SlOsaJExMaPrk5
ZAJfaFPSd2Vo9/59nRa42ZGZsWwjKNKjXwoR2edr7ADeg32aSB2h3kaNn8ftE2yXwJ//SIm+FeZu
/Ru09rwmTs+qpD7PtNift3D0Y0zW8WO2OEGGVo1II1fRVRNT2mGzhZeUwpjSUVTyovcVm3GKuQd4
0POpz4HWikk9RgCFvvb0sip6CTohVjec0/cr83fGqeLHh2MwTBmyph7GWn/avwvM9Rlbpg+OdTuY
d6I+1042quJ5v6FcooQFUz+0omMWGTYU6cE7BwXAr4TgiakRULV7u8lJ2p9zWOqDtrAwMfpxUxof
QCbIfY87ciehYHXFC02oMl+2hGpHQa9binJqmf3+skwqxU6UmjheEn4l9Vv1WNrp3FkQ/UheOtqX
krvkGLZ71vYa6A2U0Nz+qTlYZphtSI7q2wN5URCeoMdam0r/iaYA/FfxCr1NkbscfXYacVFkiVWN
N9MoEr8pAyLkX8RFuVk9heiNL3cDJb/lVBf174goeFPyA2T1Qdf0BLn+GADxUcEjJFmIICU77oy0
NoXxXq6rPFi30ndQ2VRGVL5B8UlbNhrMawQmbqNqNwhuOH5xX1Gix8r0A4n64HWmUUPLwcqmEEhf
ZwY0t7VM/emAqznchBK7vo4mqqAv2H+4f9D2J1FG1G4hqrV9eltuJCzYQNLgeVTrWIm361E7pk2s
qNwp0Zo+3jPdqw5JSGZ9ETQszBpBuUYLHBbrfcloPxmx5eiARIMVexLYAtqsDzj4kZNpv49gFujI
S4EZH+zuOgWTO59j76ESJ/t6wiRs6UB6eAaxqtuWRDXFVyshhNnSNCG6OnCoOfGQLiY3xmVG698D
A81KYPfpH88uq+YDphXN8b8/krI5N6wB7X8KOwhhTaqpvBW4RPolkblBjk4VBVPgHowtC57keZKY
5+cPrC3wfuhn/j/kZi6mAtJAqyYNq/sctNV4MTyB/YOqoysHhIXyo+n4D1kV9G5z1ZuOUIfq9Gz2
pNv++OmpZz4hCLwxR5ad3Oi38sGX6rwUTxeGUdDHmr5GmFZQ/F27Qcnm2s9+EeoEAzELL2zdg+7z
zsLmL3d3D/tE0WmAWRwRLlXpq3OKH1M00jNcSnHa51xiB6kYokMe/hKOxTSu3M9AQK6D+Ximx3gu
eiZ80rd0aPRURC1b9bCn9/NiaMvM0qNdZ3NQo/hKUYwTBpe/vIWCout8sx+h2niSUUX5LWzHuQQ/
P6MbwR+cIfpbNnSSRbV9gNnN9b5yIVwdraag1meCAIaK9H8rEGB1GkJRlrrgOo8ecvD74NUOrdoM
X0bfzwQxMoxcMy4+qhN9+XF7T6OD56siCDjdyCsSwlkeisgmuEZxG/V6Wi2tKJSY/9gsyowCg8FJ
r0aJ7JQUwF69ClhWmP3NtE0blGmQJkl6g7Jiok8Ehxf/iaJEiREEnycEWwxEtoqW48nPvvZKSes0
hPzd3l6syPALb50hnTtNPj8/qUzSIfugD9d8o3rXMWnKIt0ge6AYY087rPPRCZsl9balfR3yPcm0
R5V/2nwHsEA4eRx+InNkGyIL49tRi3aLenvUsfA6F5Pi+2Cjk2oemw8zf2EE8X6gkAz1NcCHNMef
uzCFQLFqUQx54Ig1jSNgBkOul38P+uLGcVENLmAD4OGZRukik0HPax9gg72lt7h9kOZvbHhLQWih
lL4ML9I/aseZLTP1QXryCrEiWC7NhROHOsN3v4RXo/kPO7ngIcEGeSuFaKxejR1/5D1oMvhPj2y4
WixnhsBy+Ogg+/OSxR4pIx+GNs3atWRRtArV3PrFN7fYyXY6zbQ4ImHW0EGWmzBtrCbHxarBzG6e
+hbJwRG65Hv5DNOHYmvXQ11QZurEoD87DXQ7U5XUMz8QKP/pBjuMbcFEq9uETHuooC1bKfvnTlYV
X1nqQ1VXLkIYpUCpQgR1CMcKAH+O2yVqYt+7WiHWXdqdMoO0hGrqWlDfwHn9eWaXTJQRA0tEPd9z
do0xoEeG1XN1EQYJ5Gf04nKzESdITBdy+AJ11EK3+haMyAkQD4Y/sTc4/95gDD35nVPkNOCdbIxm
b+K9st7FhHQPkU7AscYushR63C12Xr2Zkx+ETXbE1yIRIF/u+REGMIMxELobl028AwOtRY5W+cal
SDw0UDWB573FtgBySLKa5QYh6ipkuabKzFpsnBPiX2bgOXI+K0ymUfJtSZLzgSWfb+iAVdqkyNpP
pJ0mGVyt1zcF8Bg3nOpWpy/BnoqAox7J2DB1Kc1BDXj3fGGpKoqeyWou27m22Hd/2/aRc5y/xknf
XC2cBChkv6yffM44hYrrinyFfabx96DdlabD3Pq5+a2IdbniPMXqt1yn+MG8DRIl+MpfewzEBaiT
4p6/NhM/bFSu0MufFN+VNG0Y1Li2cOiwnuHF4caDQFBpbDUyrFZhKCpUpGOQX9TabDzeQSOU4jj6
gkYflW4aS5Hwe3pqywnEk5PZlqAYcA/Sep9kYxCGlDYgIDnNJSeaM1YPz2NMV0HkwdCQMWNZzpIn
8ifRnkXEXJJ1CJD+mJmy/qiP9I/sAqtSsQvlAgBOWL7/CXiAXVYJYDQ7q5ZNLI9OWjwDINX71kCN
iFGNVsjqALXqEJaYTnNIfPIVNXInkCuSzdib7HQZvWiJ7tkC4HvyGyjSyJGguEu87Os2W5sII0tj
M2SVNIbs1LXuhCcoXRPF9eX0K+G/eotN6HStxkiBuLRZrLYCq1LD15v871I48NdlexJTWO0mW8T7
Zqn1GRO5WX8HJpZeGsD+JSpCqlreGL6rp19OqzR3nHgIgUs37WidRFMgMuUX4GwLcbxudtWekOke
XAALOPXSweTxRHrSouJh6XV18c7BgSrvizEHVyv/xezAevc6Z705ItNb4HWji8OC+wJ55lPt3rSo
1mUxwlWRG5LTYoQGcoDeI4G179j2JvCk8oFFrLO/KZWCKaZeedqIr6X5XS5gp2E7KGsgWc6OmgLT
ZIcmkloPUMV39Er7wsoztf/Jm9CGEnllomqGPmwNSueuhjqF1i4mbl8Umeu7xXZaTH/w1uaAFFtb
VqHgoom9E3fauYZxesaDBnsJSrBmJ5k/dpuXqCFc52CBa/WQdbHj/64JwDZBG9tGga02K7fwiZxh
9/gcf5s/jOHUOmMMYup8QpQfR9DkTlN3b9VugpzhJRa7wC437OEj/bc5b9GVrA5PjA/TbCKme+pg
IMP2k7tVfCZ6tOka619RUNMdXP1NvEm6btwOZvblu0GQG9d1tTdZyjD7Yk9iHNQ5frYqVZubnO+h
TidO89SDptr59itxzLIjWqN5qOUKbTZ1WQKuQ4QxTt2aYdoqEAUuA3LnuM3iXbH3cvHifOiIVAUL
kJGlJxaXyEKQ2aD5lo1GEVrPrOQgH2VVf4bFuyWzRUGCvpp+Qfxagmo5LmSxL/Q8Dz4/QkwEbeTU
2CIPybFzuqr/ljVYeuzEpUDDCEXYYnO0M+IB830WOYyzOvI48vbD9y1jMc9vz9E5wQeoFMNlayYJ
n+s5fF6Zta/xf1g1KzLQ0c5bPPadvSPPR8632wpkl6kkYCWLz/zUCJvunu49XIRriBlfDsZto/iH
/nYWdjvjmYKq9CUbVwXBxVSioNWLiP74inEn16Rd1+kS13XG8N/JEK1CPkM8cR7/yzSrdp7a4/r2
wpP2V2l0Tpl0OufZYPn4wpji8EqWT4nJdNRXT2meU/nHqg23y/oo+8h8lqd0VcwEtqL9sIiluvMN
ymYWs+T85nOoLyeoaWNtScLtEVg4TYd7iKqaV1jZaKV9g6dMQ7/XhHkGvK9v5a/MG4iqUp0E+EPT
CxJdC2+6gxiAoZ+7A58e4NfY9q809R8jy3vRZSQNddE0S4S/navcJhlwd6ouCj7GZ/ayScwQs3v5
kNgsbkGUI0nyX+cOTLU+qhANf6lMOhUnLQAUiYQ7DPitbHURQHjYJAeHFh0zIjPgmnb6mUkhdJHh
yjIWiP1GwhL1FIpvP5SwfQs7UyVfnNrF9kC/z96FFDOx7+o2x9XC3uCLpjs23ROS4Gm/na4C3Vop
p4ruNEnyiaVcFDCAcEgkMfcKD3OBZS0ZIWWNaQTiy4sbsw42+V/1G043OWUmADUJ6xP1n+qJ7ZJ2
359N6dlttNRi39e39/Kcw8kGgPim0kX1S8tjjZbAJDfORSyl7J9QN4ALDWgDbbDcw0ETjrFwVXkh
MdSaZlT8QKqS52XL5mLtwDoffDcOoxVSZN29hKxmD/Z3Gyrt5JCoeY4yERRs2AxJ0Vc42fQzGRmF
PSCb6cq6EllUVMnZbiOVhY5usTSCY6OoAc+rr1t/kfzwkS2KUIXqZDOGizJ/9PKw9f1hPWoKkcXq
x9+cdu37ALcZA85g/Y1OHPJY7D+22d760OMdMgS3y8t3flc8Fnc7iAXhQu508jHC3GvYRQu0kEK3
0zraT9FuCSAmKgFeHTN6ZR7w6oYmCcix1K0j+RCs7kZ+Iwmt0u2m0K7wfbW0Su3bvoZR7wSCL6Eg
gYOqVAgiSsvi4bple2tIKfJPyQEG1+szY+Ap6w6rmDx8ZKVOJA+A68L3zGxYn+PtUx/+Tchljl/R
1gT0kRQdKWAYHkM6FEvL+7Hzschg4rwXtTU6LCOoJcDv7BV3dWaMeEWY59jbNy7/DyW07UWwhQHb
edNB57cwLRXDQiAt4a6IuXiYfRwxqXaMdud2oSH75HmqTDpI4Zhv7dheWD8QB31aYmzdUfMqmzam
wQVagtoIPDOcPyDK0DNwkeDd4pa0FLJ16hjiB82A7jTP8B4ufNXqn6l2UMb1EmcltNe/zEggDMJb
cijVYbKYcXbyKGZyciovAYI2/cAKRD3G8R49NxinNqp0H0w3JGvQPQ8G5mwS8OpJSy65NpUQ5y5r
fBS1MnQS3Ml8HTGsDkMTeFvzjhAlIZrYZ/HFRtAAyfqLjoMGZbD8tYlJhzP1Ytc+rWDefqYrcZME
2a7aGHlp5FzezMNWYbsei6fOdvH1aisZLOjgkcck043NFkn/D2jKlOhMlCuNPT1/PliwYBeM3syg
HgUNEBTBCnOhTAnujR93Nya625nsUGLaNU3BniYUHYx+UlQRtLybbAFvo+V2RnNquEtorI4JzbkY
KeYghHiJixBDPpCLIu7ZxDwCKFZ1hndSC9WyItLTyZcnm6jrRcrs4jhmA+tJ1xY/u2AP6V/rA3KY
+tBVnvcO6YlD5PND4JRNCqgUY3PqBTZ12r6of4asJWHnrvUTJ/XWvxWIzdBCPQYEkmvbAMqiGz9l
QVndoHn/iMtsqoCa9/2oE7IWaFeiECYhcyynS4LkgEKAZIQFp/Y9jss7iZmHGcaawJJyFibJwZPX
XVVWOab8KOKF3MiBqUt/hEeXNgmrAJkuXH4V52+N/VROqIAs2xv2+6KNVsQlYmawx/n3VNixRcAj
7NxDo/H2r39zVsDr6NJKj+F0KULOTwqbFtCQY6SaNGPsQYwAHXDIdsXgc/Vs7JrzekkYEwwcWa77
SNSAoT7bJT56fEttJXg6DUtVGtVo7MlTTDzn7lQULoY0ShuAUbAcpkeYTAfdKbAs5q1++yBDIitt
4FgY25/Dk4Rwc8GuwfIVF4pGxZ0LfRgZ1o0+DIbn3khxM0CPmmxEAr/T6XMhtHvx3VdeSLDjAbY1
7zg/NZdV0Pr8FSX+G/gaNy5UyGTCZJ8P9Y/5eP0xji5T6/7PQS41A2ROFvsTz9FM32k6eYq6EN2K
IPvDB5qdAOEXxyoARrmMMu9RYbbTt1FSuaqGFpzZa8vdUd4x0a3AzgWLFxTjtetGB3cxN5UUat5y
Q9kj7W6ZY6V4xfVShjynkqkmeCCGCLv/LUNOyCks36iV3+R8J/rvA5sJdWbb7XBdocDmi+Ycr6LF
gMjWXdnMfJkRxrWFrhbtL0t4oIPRBZDv/vaUpj0FBekwzLniAor7xsjv6Z7pH3B+Cdkkl/AV/DIY
mlNBGbw65/4Pe/YPGtlRgyg4LzX7wgpNQNz/R9nNAjzHNz5ptrQUCWedcH8Nj3cmYa1PF3OMmkgW
mY18KwkFEk52Jtw6DT7Gsejb4WsoV9U3IY+oryF+1Z8ZKgGR0okHEZweE0BbKGjIVc4VNtR3ljTq
6j/+gH5FZViLXHp4SNYEzHfupEgXiJNlk+1fmewb7/3eJZEAkOWlNUXXQRaDKcwagm/XQjqO9KVX
CPo88+Qlul5pv4bDxWvof+2j9qL14A0KzlA5U6c6ny8f2iCgPujopgemXtjgSEW0V8YW66+qpUTQ
YNv+sI/BMGGJxUutkknaiA5vh1GD+2sReuckX4qgfTDVL7ucfF3UccQIqNLXs2FASAyDRwxRKNxE
ByZ3SqGUVG0BZeG+CmR4S5v9XLXDx4i90JZhhsVkfXQlpfCXPBMM1rfWJoqFotVrjXCmMcXTl0zP
FO3u/039tAiAI48S2I5R62veqkDznWEMmNFVI/kNqxQ+kdSmY9TwVy+rt/7kfMWC84TxIxzPgQxb
Q9oyQXa0RQTMId9r1OsMa3XbVwNpgyCRFHoAqUw0mgA8BWTVIAMal6azfJQR4PRBaojtAdVqQ9Gf
X2hu+AWIdoxxFLkhu4w31Kr/h3jcV2UGhkLiPRxZ0bHTcne0one3SMBgTTd4krceMgViXgdEbDXQ
K8WpIkSv4q/rdR76lU+1Yw/SFijqvvwV42oTAYzW468alZ/QdDJn8LOgEl44vtMh2deXQNYiAnZL
fsmKntG3IAMDPksyQGkeEyLqWziHVC0q5i6wcEDpbIVWL5mZrYLOueD0x5KQ7LOK5qdsVfg2jB6d
TGFi+3L+/4MP8SBQDKi1oJ4GCzbRiF5qEYC6eC1GCz15mHYtPCDf6orB2a7HOrEOeVahO5hV4FiG
7D13fmUmtrYQoXU8KpwbN0CPSfUWN53xrU70x2HzrJpQxOtKpKKUNzgzr5FFssScKcDd4LYiQYK3
bWrKCCa7yvq9JKX0CMKidCMxC14xxVb56ZVuoVMYSyKeZGOerv6cHoOE90pPDpRRHu/eJJTYschS
SANNaaP+5uNCwcK/JXlpLTOt7xRYac62bH6AnYWMeTRnNGxK5uujpuZftKBdT8+MT/Q83iSs+wUF
ecIM/8dLAcBsGpzaxebv2bGkQk3W2rzhGw/YvmrUwg//0YZneKOxBkjc2MLL3QRTwx9Oty2JahOh
TfDfY81UTYLUdGfY0qJg8iwB20ffW1il3o5zKpsvFd+0ANtE8TprNnJlVoLXCIRinhbHjgIJajY7
xa636fGaq9TI6lfZjM7e2tvKOD56w2HJK2fQT2fDmGSH+TpaJRYXFGKz6ZG00E0obZ808BjGd2+b
cltUnkoARmVYcSkKJEoMOl2kFSUIOwEKWPSHCOKyY/0C6I4fN56IR3+MktYfqSkWtyFt7pVVCiLE
nQuJsSjVckDRdnZAHUYqQcZi8JbjQPo4YuCnc8lCnSQk+z1wKVhIexZzQM0C2Gc4R/xYXTyCbBOY
+mqoXhjQv0Bfv9Rw2vMSClOBLFNyGFFvRbNdwbioCFT0o6KCoX81FKseyYuJ/3wUqpSTofVnkZ6H
Lwo1jR4WXtLcV8l4XfPu3unME+VBEQX70vwWALKhPRV3ppch1VQ0uX0MOEgCed5e8gNBk1cirm3B
6tLhNgne9RnfqhVOsyjQSYNSI7rBxsH2vNONlQeiKymwfc1OxcoKoQ6cpsWoljUC0cJMUbIuKmgM
HrDE0eTpe7Jd4eVbM0OFZQ43BeD2TPNZ/trTzQsjF+qadgb/5fRdEy8B3c4tAP/YkpHkrZfbMIIK
va98QdPB310YA2oEBLD7aL4O28dn6chyBuOapnGTWJLZ8OM14hcNEgJRuyXcComGORKxaQRhlKqA
hDwKsbVyW4dnMaZFX5uZ7igdykenfIeXRohMEL/wrlfZovWDrKODkxvn18tv56lHMF97+3EqSu8u
tuDiCYu0+hbGEDbJHGeHpOl1PqV0v6VAzN7bZkGSyQ911S6pejV9nY8QqPXzFszXfo4I+l5LjReE
NxKrasLyAkyloi1JoKbaFmB7tEDw0U27PpPEM2896OK4QnHnT7eY87F5y90gU1a8a/RpuxsEeiVm
lmcflygYHVp2Tm/jp4F/6YXVZ6DBwaDhwdqkcYKKR7N4qaAWSBUcuPwPWMuBgFQgYqksZFhioGLC
5Jz7dFPj+Sy19ziRmr01ZSck3FeomGDPtCYNP15wj6TZd7gbZ3BiFXlY4015AVLOVuENDESReyy2
3d1R+HuPx2AdLyBpmmdfnvE4KHtQMDvz60Wrx0SJU3HFUOy5NREUEmU8/ngGLte9cwmx/F1FvoFJ
Hw4bBXKyu8rbDK3TtlJcTymwZTqOS+yrcL79Rsn5Bg3ZQZlKCEE3mJ71HFstU2IaTtV6woXAVYkC
Az8qvMvqmrIjR0QF80Wc7n8kdOcjGZdVGqRi2bq1GO0beLG+62y3EBuOmPTViQpKW6UmaEOoP3h5
PvAxMdqwvCggewztyioNOOTtuv4UJrKGwJWJYmsEudUSa/2Q1w+rjVB7oxYBJdb8eWJ/9VwPV6OA
l7LxZxlfxxF4XhfrlR7tPkrVJeR4HqjWl7BE0bu2iNV8Dy9jz4DIhTuKbKZLda+CWIfUnwAAZiio
2W0KT+FqjaXB0LuPNO+v0Wo95bp0HmfUOO36fKoXPPkBY6O371ld+4eB4nYGvldXrJcR5TCZn6l6
H5EAd7LDuCVMLc6dHiOJfL48miHT4zmmx1YVGUydiFCbsYz4mcBZc175ua+5UZS8yYTEA63WryBy
eZb0jhJgUG9v6Me01AZsfF9s2nalletF6QzPvgRi975cVzfbApHodrVgSfKTlNEka36KhV5mGYfA
3rzRVqR208DddRzPdqZ5HxaqcgVME0mD7HE2qYjyJQ3jsryW6V9EWAufsan3p1aBRKwmQwbhg+2b
iQBbwZo8I4R3wsMEKw4oOkSVVWDtopRLSEXG2QXbGcRLM7qMmopI0rv147kqNzkwmbWm+Dj6GHn0
DksIHsrxOIH255tsWDtTYlRSe0iz6fwzvrsTDl20cjzdoMMUwXzropu9z5Iop5KtMPbYdXGPcqgQ
ynav11ab1yrdscJIo39/pKhdG7OV4X/wNunlRd41a+FPIjZB3F6zGwadl+tvpuo/hfcwQBTI3HkF
2STnVI9QXMnkWCfX4HecJx9SiWVyd+vnHUHS6V+qvzVRLPVImUwa1wWl7XMGXfA9VSbOYs4eui6v
N88m7BTlRPd/XcFfs+Zhngp8DUa9FoB9fYZfWqW+ZLSW8syHI1ht2+AB9Y06PTib/7I4ubTzHEbE
whQuzZHDIAQI/b01i1fshwbdhrTaDZfNPDgOBghBWo3a5pwxdeo2lK8JiiilbBH7Yp77D9x+X791
Hb0TYakwPdMBzJXsHDsprZ/bc1HbrwjmC8qgJ1VO6ZMhYxyvv1m0LT+G5BdQDiHFhBRfiE6yDEV9
aS+wDnrduMPqWxw/8piAnVGXkzxA8HW+cOSnwTh6XzslNWx3qjBsRECiRaI+fm3YVES+NlsozZ4k
8K4OHpunzioVYCGhaPL3wnK+MIs1etTSqNoviNJyanEQ71O1ETQgXYUzNvmKsmlMOvviXCo4Kgd9
M5z9EgecFIfggU73rXeyJjtZMz0jKNpevLtoyuqO9//K9rF25NyzOB5ZtcPsXpKaC2Yb99TJTucR
wIuor3EIocNGRzkxbvrvccC4AfU7swjJ1KvDSiP1vIGlEkGl2fSb7hROc6ntC/vbZkQw+IlSM0It
dX8wnyHRmimb1rCw+H1ssyzU2F0nJTztLZ94AeLIytv7LR36WkASpEJisZUpUrXZ9YFIfMHu6EW6
pZoFFg/EAIQmXc7rgJvo8S3zaNteNZ96rUhl1j5z7oMKiiroB1uV04kFAANbSCRwxeVSvyIE+Iht
VnJ30SDqdy1Qq48aHQeQUluwYf0ghOT9mQbinFj7gG1EtSeeYPdyTBcofvK17LOWi1u9hF9hF8bK
BumePyRz9X4OCJYntGA21wYm3nNc9Ztf9QPgSieGBvivYt38lQQgMemgDwgIlqz3M+NFBDN6FYcD
M1CeUNOOivjtCKHL8kV1f/feJ74ekBi8JBrrIwJvLrM4fgLEArFzRDHQu0OF2KYYxoXIcfFFFMHy
6aVLyiFZlOhcOugQOYYF+hxsdOSmbgRGirxHVfkhcW2hOTaPN8JXqYTSRmoELYiM8HPaLHzhIe8T
qNXJPNbGr3wfrOK0bgB6Ux4At6fi/KNK6yVlxlAd8BZLueiYOXDXUdPAL+jjQ/3C8j+dihZNXZfN
IWwKaziKaRHdzjG/EIl+OhsawGq3RfixJmlnYa8RJ8H8TSuDjEGj56mjbI2QgmqfOu+7VtLSgfF6
iNa5LLxsOi2V3hcpW7K4IqmUk1+HPxc70tys9DmLGqgA1sG00NTPF/NWoPY9APnlgA5WAl9M0eBS
ckX59zyO07Rz/sB27VJRT6+IE1FMH87p44fn53WHcX/dGwEZ1x69//6B1RDV2UvInFd+9FanLWj2
YNZdJE/5osEKiwpo2fe+Xwz1845TPiLUdCyy4ZexyTYOOKi/P8Je9ynnrC0oUDUWnRKZcsoxMQTU
BgfeYgRbF3r3CZrNDMbTsdGQHH1SN+ESCks3DW6QkMWD/HzlN9BbnWGjzfqddvMkSvQNYAulNfmV
8DPF35mK0l73voweCh+YJHmA9oz0Yc37qOju3i0ivXj0xCkii4+MJP56aQow/KIB6je55WMqKbuc
eJI7+i9HHghPfonJnPfz3t+KnfQVBR73r2n/Ub1uZg8ylNn8ubkurt4/WA4DyMWUQ/0f+df62H65
UrfxZKsKdsRlt1DF+eLAlTMtwooG7G/MMiQo0b3eHXYSlWi/lY4diTHGDA1rB+tWXZdf7HDY/ESh
XCMolA0icJ5f0WcBBgaKC26M9YrVsO9yKrtMd7he2FvdEtRgo1BSrxdKMVNwHg/UnDVNqvJgrq5Y
Jxc1oDehrYIV9CtjAkxXGlY7SHsZyzrIVWQFb3i01vZoftIUJnhCEEt54FtRINq60IzYSiQF9n5q
kpB5I0KaWoWNLTF0DaZBl3KYV6i6Xzz7PcGRb2dB/XdgNCytvDyKpWHHi2VYF5WyWCxnOTHS7tQo
33UvDI+X/qmXAX+vc8ZxbOgGLOtHHUvQQQwJLG0ECqWCuAFl2qHh/XkCmClJulvUjBL/ZwwXa1uL
rbQRHwInS1MeYPvOrf0B9huJzj3D68t/ip0gjFJehvJwzOgFh2Xuio39bti4r4EmV+mEz/Yf/v3i
jy4aXpsnwTSVKB72sY1b25lAA0rmhalVojaabjhDLN2MbPBZhqER1HCvYOtnOUZ+retTNYVvZ6ju
5OToF0jEMNB2RbCVfhGfw26wuJdPGX2qhiBIRzSn5vAcQuoveq5zEKX11P78ZJzzwrPxqLZ4dGKj
CcLmQpcfXXcVLjLXGCGE3/stA95+H+Y4aJXNv50LALoO+IAsHDamgCra6Wn7BIoaSjuHi7v2vOLe
eADndgDsYXgKGE9FdkW4Uj+mk2ERtDVWUDLvokyB6jn1owvpTDpsmDViFNbVqd0zu7dK5/12Ofz3
Atav9qDH3VrT9JGEzzf+5Ww2iGJMo/kKD/IdAk/o4/4AQcMJQq1/JjfRqv5F6rzoxNQ6+QSOeBcd
okpMEQQ/fDJS8egGttXndpc5Kdaz4aLuqhodypXDcFlp8L9HhLSOnunerHNRM9Wf8lIVf/rB5q/r
o7mXAAvQ/wn1j1P2iwz3mZB6ACVgzW+qzGa3tA54QpB4uM63ZmpsYQEqgDk4W8k37R6Qkn0FIc/F
jmDjmFNIbq7pJmhJs+v5Fuf0kWUrPON6eT783DYP7vvvB5X9kG9ZMG3fvIy8Iw2uz6/ouj6wZApq
BKXRBgrkXHQCiy2g6ggTa5hHtlxfCTfmpKJBDe2Z5Xo+8vAzP7vhnXc+h5qdVE3AGpYKh94FNICH
P7ajyO8gPIdsh//NM+1EFTQnjgfcW/vQOs/A8DnWWlok/n7gU60r1f2neEAUFxEG4+1J6pAkJ1dm
pHem2mMnbRyxjPjC6b2SJmIOQmoz3onBY4Qpgf55ySiW6PKd7KzxwqUlpx/b1oIeQKh2O+Pd6w9c
F2tu9l3N7h9acskQzAfEaQNIRjPe7am52Qq7Rekki3kq2EolSfe2vCF4MIuhbX9EOHOLl+yXv3X7
CaQU3ggfrebVEkcmeCtX5I1G8t7SUp2Rz8FhvuWPUlbz59EYfKdVbbtX6TLkCeC/emMSJfn9jspj
NZUOTcB97fIRXa2H+yMb7ZCfwxbkzwgS0btebCERwIfip2EuU/uZoaTSqdsOF+kwqXQiv0chI05r
6R7Di6v9L2Q8VuRpx09LIr5iqwWhw9RbuQUPKcwiQ5Xl11V+aTbwd4dacOv7HJ57/5I9xHhwqql5
UVR+C/+QxvXp8AhmtT7TN+N3UPpbMz2kmX9xH998urShyX6ofl3MsQNxQI4N8711DHw7nd5T+UlE
AbI1W843Taot5rTov/sj+Eq46KxKRXM2l8m7NCbOQI4xmtjs31HSggpxASXUnX4rR8pRVPtn93QO
IrNIPscvNELdIOtwKPOGLy4ovHy4A6GuPzXMXq8Jq4zGKYox1TtXyNvdMizR26r2rHApCfXfeVAt
F7ck4M4BHDr7F/vdDCeTqUOs9n+z6caj/9qdUBsPbiDKYYxowBHpGJ9CdB3VscyYZViPA1o1mi9b
nhWl6KuMnGk1mSHX+mLzhL9JYcQ4DNpUSU03SZs/CK0LvGaAsgew/Rz3Mjq2FQhJfoE3AUP3VzLO
uI/Ts5a99o/uFps19lfL/rjAaf9j2VaK1tSKKimQPtl50ml6maDr/IcWdKkyasUXOL9Y+DhLKC/q
yPkhAW8lD+NIbOSrb8YdSPAxRHUJODKO17LdgyF85lI3DhhH1vVHp6a9Hd5TYxevt5U8rPWJ0LSN
XHrAwntXgoeUF/J8X9ZKQk1ah+lZtYEnlDNQEK4unZ+2q8MJJQUC7TLuJL29/sdQLluR0cOUcCE+
dApYW9TVwOWwKaa7feabrfJVpYhYPM5XZzSBvqpz18Orq7wCuD9kvjqxPZG411rXfczE8TykH//A
vmZl3DkWTM/zt2kYQwlYDzBSk06KLhZIXjqPqzTvKnY5VDqI2dycQ5U7eTWoiqm/74T/MnO43ge6
ltURpgDIJSx24529uQMMIXNeWzdWcd9HELDZjTSC0mnsiPx9/918uvtzdCecVtTMP87PyUM6Z3J2
9ZPBH5OP05HzI6OrpqS8qPMGdmwr5rRmLO7HBThvW91XsqGolVPqvxW4NhoB1LGsea8YfDteZz4s
ycSYPZzc9mSP1GKVjPRiB1D5ZAu1yEEPu5sSGJLntL80KD7rv6x2V69/Ll8wfcQ0c+PFZIG2t/l5
4Bfp0HyTLCAQpmfjNOEeS7nCDOPeBFzpN8L3tL0QQqnNoo7RgdQsJIIogXPaRmUQtHxjB0dPriGH
9bqJeFoeq9ZsN9q37OdwfublhFKPXYb0dpzSeP9/QVzGWOF0UsxCsYKidNoLQud4YkdT7dG72ups
76KiZTSQRvjNiepyXf/djeffSJImzFDI4LYXUCcDxB7Rv3lOzs6laTlHUrgkcdM1QGL4CFj2U/dh
HO8BQsHo0VCPD00QdJbYUs35JktPauoVg0LSjzcLhlmBxQVhgh3MFFDvxooMQOF4H/5a7NTOpXaK
7DNUpNMHGHn/xofRIQrYaFvaWhQAfikB1UKtva+gUQBlpJxJCPMr8D7EEbRzFeypOnOQ9odZh4Gl
o6F5Pt+aOI4Kpm7dgNkJhg1MPNf7TAHfFgTbdVk3bCrwWIsBQovi7/m2PUbWLkihBeHOvA7LtoNz
VL/7uHSKanFB8//gbeWFddunqjJqx5Y4VhP8D1ht8RYoKUd4ezCAo1WrU2v256c7OU7DYfIkfkCp
1x1QbEbQNzd2j92xZswhltLEOVlJCnn5su8gggTXeOdBgOsae9C18I2RZztW8HUj6ggRokQcDx0J
UJMJbiQMw4ysDHmS1R2G5lcW41m4LLdZKRTFGPiWsHURgcihoR+Z9lA2OTzDlVsMjXu6F+4ZrqQP
Mzcw43AxCrpxOsyQz7GfnVlrycfDYNWqyhsUmgTb4TaS5F0PJ/gvTYdmb+dPXY0XegPKTG5h7Yb1
S0vtjHHsmJ+KyeY8ha8fxRTV6zO8UIFtwEmxRjk/gFyWnqwg/y10mGc9CM+AYS/lJPgSvloT7jek
jVETIKiJA/VPhm3ptkML6i/CGE0sV0aHOwm/+k6Xvvo//CV0l5v51TP+n//J2V3ccTxFtIj2QQTS
RctiyFj+M1GHj9yrZKe3Chac+jkhkTV/kVifAd16IlsFylxb/roTB2/omYmFN58cOpmvdmg3e5VT
TW/0DeA1SPVovrzXhBuXIBDvDqk47zzlXZPvw4B5jLRug11qHkghIFeyQ3UNc4u3sd2AvWypR1vj
w+jQe1Lo5Fwog0GE3c4NBkhUnBvGLTZuCPwoftjRDptlM+LKtmeare5SWTPeFv+GaQiuw+ObTn4R
eiMX1FuQjGIuTBb8a8IjVHyK4t2GuQTF1Hyu7gm6P5Eu21vhs9AEcOWbnRbWV4oYm3tJ55qmAGqD
3wwm+Cjq4L9mEpGzPMG8i2BhoD0ivJI1KgLG86KME6Fr+orXLNilWyhFjlwU9UVlb//EuDnFXIgZ
9YrJ4HNtB6jhKh+YgPUXi3XPyyGyS3uSBMiAgowebimo7hJIYrSncUOkoMttLLGSrkh9ton0Jjpb
Do5LhPNHi2LP159q9QNbeTkF1p4VM6K7wBhr+j00kcXKWkF19/dFgpVmcFfo+xyjmZt2HJwPT+Rj
8TyD2FK1U8k8oja8QPynVuVVG0hExrAZ7cVIG1s12nAi65PV5SbJr2foYd29mro7tgEdLiruyEzM
HdaLZRLMcgz6T32EMrTeSPlHZDpxIIvOR0YZ8/HIUtCu7lddZle0lnYtck1hVzoowbcGf3I0G7xK
mH1ElwraWE0JQByrZfUBMpVqxbZB9cM49ECfCBhklHNe3Nn0l9t9bY7WZfqqKTAJbSodLPGOjEMG
cDS/SrCZtdJOWAvFsSS1gjbCes7XgKeqgWT5L6/bOpYKJ/OaTjXXv+giXVox56omI2AZy7tCLqy/
44qQB0acg7gt3CRJMrvc0o4pVCK4xGRA0LEK9zmxBEkxp4ePgT6HZIdpXIohSWPWHigAtpdGWLUo
Sfd6gY5COPgM8rVzs/89nwP2PrrshLO8I8Z2fcQAmLH8w0LdVTFulDiD/GTUvdXDuC5M4XQpdfDy
b+3tQMqOOzJIb6HhurTwsVB4qRAKGfJ/hKFuq9x1oIE4uQIjlFmD4ozMBTzJ5u49AJu1EXQQiX8t
UAwq6yBUKlG+xOw5C4gTUPhxGwQchvk6eU/pQN+2MlNp7UvU0L7X48Li4sN7Y07NBXD8IbHy3zVS
zyZL6tO9GHisSLV4bUOL52p+HVqMFgeY9DGUgwQne2TJAnYUuupPBqW0d1sJJvaaCSdVFih6I98a
3msLfXSMbwX+vQpFuVNdsXRacRxOoOs6jA/z2FmSu9bNIzjxwXejocJ4RphTizEbU5IcvTPfFUDl
b6DlxQ2tSvcIZp6vaGI7GZ7Uuq7TJBiWiB/ShKSJff8Oxqe5PtP3D+bSIa469/OtM4NPlthT8S4K
QNaJMTDwapBxRYo87P/iosEkA32liFHg/OsVLhHT2GKo5s+QO+5Q1wdiVcdl/3pUPjxG6jhkun/o
wuSdbJsPDhJZ2BZqOGmKQYd1Gm1G5irvg7e/bhJz7IM/QVul/aW6uf2hXce3MBOaS7WsM1xdz07Q
RbxOuAZHFJMCekrjVO1HMIW0+nkMJ4IvD3nV/WiY3WNJV2mWkNQbQ1mqjSj9aELzQaZpcxdvlPcQ
T2FGywLiDrhptAejXb7nXtobFOIaZrxdUiyhvtJPKpEKoQmHzuvLa83Ipn+MhWtajZLN5NTuYIEW
1SLk6r5zeDfbFBMxK+fp1V/qPR5zUOZKq8Io9IU/l5GRloqyQdwDaHPDinp670wWnYTLeMXf0Q9+
Bu2X0J7SsdAz6OFwTgcmgmffm0qB4B1Q7CGCAiXVE3oPUW1Dv6XhXe4uoj01d1t71lhmh34lMMqq
NTWrPf5Of8HjRaxlHmT73loOP41AXYy5Ajqodn8+e2bT94FRqY8I9A8SlEtfBJ0O79h6sDTI7/Pq
fWnyFSSSfSI+/uA2i7FVAI2IEtjWBCi5J99zD/SWeYFDmAYwpFWd2M8ITchfQ1vLLbQqseqXtfw0
+gU/lm1qF1CAnk2/YY+PdnMCz/gvUwa5MKFknpZUGGf3K0BNsfHF19xs3ckObBPcRx1TAQc66pWZ
cxQ4Nl4OCTJpel2c6FJByVpcXoUpwPLZAL41gg2ICP7Fs60zintgPVmTVsMAx1+D50OM63HLEq9G
K0s5vLgQO3313a66N2kCjLvq9luKLBRR1EKmPUSHkoeg2YSQeoOcD8uG3CUio/c24A/vlJo5Qb5b
SDtgUs1uiu46laJXmMzxrZ8zEy/ZXYIDy/ECuTWALOVE/nzC7MxbZDrapyqNznRNHLF0yRIrJxZ0
5Pe/79LO5idPH67qu6y4ui9gS6Vt6PPqFpp+6G4X7jfhkJDL9xdwc+I/HEI2twJTGAzhTfsKakBK
WZcl6niWQyk0JKi8oZiUhNWrvfnky3722vb624//Zf/rZZ1A25henujTA6Hz69ISQGL7m8YSitew
6OXGL6/PLHwayGWeWkeTP4Nfq2cl3MZqFsatpBILmxtybpvabBNAY8L1tW2rvhAS2chaYvypbNeu
03smYWog1EvMudVUXRohnugBZm515XNfpBdLJI3GuN8t/oDsRCxwaEcD1naZKeOi0pH1vScIOv+O
XMyqo+Ciea0rwfEJarssD0RPYehhzqSKFqXNUWlzlUlsKhfrqgQbL9PU29JMrSmcLx15kHh7L47d
oY89dfUd2mQlq4pi3pZNAkmCBTxizKz5EPbXOK2Q5unT0DguHgl2MiJ9YEihJtvfP/w7mKejG2aE
xi0jWd+qHUWeYqY5etIBihl/uqJZDDQKSP/SbsaEtT+Hs5jTVp1IupHNVmQHw5c3ifZyiPjC1Fge
/Llm5N6FyhRdCl4QEB+K30N92pt8YzH1W5AYPEZ8mbIDQ6hNGBv4E96P+IJgohrfQgk1BdKhBUM4
96S/f3EaRLGb51dUdGV1ix6GGl6ZCjMsr2ysZqaf0tf7kB66KZ67JmGG2ek0jI2BUH4mrjUrraNk
hCaqa2t0RyLBny/e5LrtNKiqBq3Ng7jIBGOjPZ7mj7OGhH7TnYGkGXWmr6x4LIVsIeMpeuoqcybH
gpCRImknq84g4YH0YgJRdYMxT8r8W5dDVyFbCj5LZMGYxUmMoHXeIydw/9J+v1aCosxvPszRZV8a
mv5Ai3sCr3LnhjGrBiR4ZDloVh6NSVNIoTgGB7IZjJfa7k8fiaoRWPNDcC1qxBYkLkpX1ySvfex8
S0AFphdtgIW36n4I6dANXlbymIwJslHYVCRZ3tdi5rpKyveDamHuBJviiCaCuTdmqWOOb2bCkdy9
S+sj+b5AZmnaQITYDYyYOyvYGleRckopAcKeS/lk4ENTkTiBW5HAfQUnNIqy239ef5W8f3OuT6al
RAUMuKpq3pKFk94kfLDE4SGe90F5g3VxJJ+sAyUhFRTe07H8bJwh/k+2W3A9uxdUNwZdGjfmZsVG
knmsS57Uz9Ycmj+G28Z1BsSDfyxKv2Ghjaw2jBqO+W+I9moCzcAFaSxUXrBOS95+6AuuCvTFm4b6
gP4+ynl4JFD1JShOaWf0uBYs1FhomLoam54y7GDV/u5BAdwCSO0ncqkkfuWm6Otx1wHk1CJFbO0N
/W8emYsj0axGxpAHZqSE0l0u2yV7MLSXemOR6PuuOilZgFvbv39/2LMa8yKTTB9XDYYI3g1g7Hye
2fGO2O0AOqhLYD2iN0rDt/rUzQmAqCsYxGOhfI3I0fm93IY+nLGDrXpC04KO4RsjS38FjZa039wF
ky7GxouN1h++uBgR4X+JTSgsGKRKVsdQJCgcaT166t89kBw/DlkigrRSAAw1ZTZXjYa6BUufA7EP
Zh3uaf34T0hbkFn0xY1MglM/V/UdY1grZiwEXjqFTPEVDYdDZqn0CXlAm09gEeAH92LemQOuIRbR
760pLF+BnU3T8p+bcZfqiSn67tredBOFjJILp8GlER4n6qBKMvQZlTCPkHKgHWYxlJqBN1ce79bp
vo/tYqaFTHKmvoHLFRsdRwO9rJ5MOJ1FeYfvTFmbPRYVu3ZmwZmK1yU0odRRTRxS4wuD814Ob6Te
qzCobepYZogtpI8HxXrFaW+Thwg9lYJwFdR3+ngcxQ917/ubtgMXUHrmw/zgeBpGkjlV4uc72txb
lL42bb5dVjcQz28dwLCLdjB/hi3ZtuXHHpizhMf1517kEeZGI1Jd75E1TlGh8TEE9WHqxkA847gV
xbYyUr7mMj5jZvCZeA8OzB5Kt+gJJSpyGSvb+5Tt+zKeKemEfGoY4fb6hGdcknr0z6dxH+C138VI
JXS3Qfr9nryrWAi4h+eXazumgPS0ebVmscWfoGp96uuRUNOhUVMAIDMSHBrezKdpePIK2X+kbwsq
Cx7B7AUFxWM8x/QDkn+1Kk01g9ytpBEAn+/zqZXV0WF70yBpoi/HIbBcwV42sqFxUEUHBS0JxM94
snT3Bxn9q89KuuZtUvUHLESm0uANyYlRYSdGomZ9v6wggRuMBmZj6jr/xTGfSOxjtb7/Q1clMxkr
2hn7YbBjLibXqOp2h/9omr23mnr8NOvLOczPgSBp2Xf7CMxQ+aiqfm3kupx+1G4kiGmM4meoYiCP
FnOBEmm1cTDmmLF/NxHVKK1a4/jYcws7ES/ei0EjxEZhVEwCmWIVXXZGo3S+yncsuDy7RQlNfQRB
8L5anLbMXQzvSWKwUOJfdirS50olXYn7P9wpYR8Yu2dno0V02cs182o/NNaSfdY1PquvNXDFG8kT
mT7x/soBJugaNCP1NPB96WFaCiJYtgWLDxFDVkvgSGAj2w4DLdUC0FRMqebrQ0mMww+HWrhM87sc
PVXAOTxCwXshDqVrUplLzMba9uQ2rKRX6+QDHuUe9gV2iVa9ralu04GVtki12Yizn+y0T/bHYf6h
5Jw/Nnr3WqtTy77bh5M29MCgS5C3rS34iz1+fSVWyMSVxfyIg4VduyrK+R4oV3Uq4sz84ClXvA8B
uIhCWjh3+t7MQlGEtFUvxLn2HvPE0sj4ey8TXKEfgjHokImK+Jtv0E84XtcYmQy/Vga+XlqbNEEw
dooyOd65nM9ci+dnlbUeg3x1t7vtcUgyN2ROMXARbSqp9/om7MN9VupcPWp3/vTOqrF1OgrDmqht
rMe/B+OcoW1cIMfBUWumOMb1uqwZeLHo7Rzf+RHO8lwi1o+WmNH1SwvHKSqTRsGaRVgW1cf2V1W6
TI8tdI7uOr7GMcV2CXr8tpVFs91XhFYPb1u+btMAFlrfaxWINtV1bGaXO1a8FVTPJ5A2UXboh1mv
i3vPPSiIf9MIA5nJdIUlYPc4cDwxdxWBFqgUfzIjfvqJj0qJQ5EM1fAFX4FjVgD2pNUzWi5Y/h5D
eh8ggv+1MeLSGHjmqVff4uXejD+tY4MA46qIgKfqalCmLBU+CahUfW7INBk6pnEgwtqQVRPu1bd0
n8b/bbzuKAf4GK3LuUpf/y18l+rGB3P6ABRBiUJ43VU1Z8GnIavujgQIn9Lj9lsjwJG1n1vXidev
FHa9e/NmdgHz+k4kkePrInDeg3HIIdAKkH1Ri6DQF7imuFdp2Qr3TcQCa42FYCOd/zrsWduTxrOT
SUDQvTk2koYAAlTbzWipegAgIREu7ChcIG5nlrf/gfPsPLdD2ilIu7ZjtCkYyYFDpBQFFfcbzCpV
eZSrjYls8qoQPkAS1ATLAQzauxpxrJReU3xZpNYIC8miLKkkT1sqqRp08phoK60y/bMqFFdCFlaz
UndTGNuNWkEmMU3E4Rj1Nw7DyBwE/Q0sikXpwhKZpUiG9Di7DH5/mJudtMOZGyqQ6oQB+S5SKgLU
8tv4Bd47HsFLSktxZS2jO9aa6sP6ZXMZSlYxwp8vAMpngMXKeGnlUWfIXSkkPLXcTGoSF7ACuRay
XI2FiEhgVQg66Ds+L0CSlWLoImHKUKBNlUhcalJvlAv5tET+sIgzkdeDOBfl+F7XZ1uu1LbIRTRB
JkSiBIvmTt3d7sdwhUJUseAJUbROzRJuXnsTh85LXEYzLPZC/ffNWuIjef2FfePEQy12cU9WcPvL
woYel2ttUGtpXEY9xA4nkoSEbucuYuc1VFP55asNE+j9zIhnta4Qj6ymiA/LhmvJkcJx8SjwQlqb
ZsdvGEsXY5V7wTNojHRGD0+BnmoSN8rnp30IuqzM0XL1S1DDKlLrreecJOb6Rgxh/Lm+yFWi+Qu4
S9GfmdUuVZ2pJTXyKNdNq7PKSHLwA5QMeYquqDCOqb2PcHrTuvxO4kaXRC/EkSL8pOvgMzBFvJYJ
tTr4kZ9RUQxpm9kZ8pAmaduqQ4yI+x6N+5mbIIQ+ypYTTaIYD2CMSWe2ALX8mw1wGUXdwbdjEtfr
7sdfNU3Q8NCXPDJokYPDjvVRtYgWPQxUJ/J7Vmv5hKdwkldriAuPvDqKuNaeMRV0Ls9s8jzWGN+z
NHI8g0yoPmaHfJjsx5auVZf6jo6vdGRPCv+iW6fpXyQmwRbPjYWlmH/GBtBEcLNzWnliOSxTu2gF
srzD9LAhk7jD1rhUNPjZ+EYcP6qoaZwnpxNCXRH0mPnSb9RIijJvl/dTpiyRqLNX/rgCfPJsHqCu
Vk33w8/vvoKlcS2/zX3SJTnQnwYaOPWQLgOp6Z4fu03SS7RO5GzgUwH3bgLHf9G2OvLQ9wUEz1Td
M+8HUmVj/wL+AM8PM8TVR5QUxp+byx5Vsx3X7O7r7ifEXuZKjO3NR4WxWn2sNtFoLYNc3uyOCs5X
wM0K3nvaOJMV2QmovFQJMdoL1e7XQ1vkgjfA6z/4qotdEJ9LOWFYd0NAU7DEnlzSRWvxvQQFbsEq
cqdvjbKDjmLIuKzd+ffDQcdoOrKETs6zY9Z8e3AbmIggV6ZfuFVLZnF0QYCJD78c7lcMp0MwOEBC
kVWm5M0JyOnbov0GUbBbdlDGZz2uVHny6NmCV4WBu0/1i21KyN+jqidgowO86ws7vT4h4Q9QFrE3
pUHvDiRjNp54nhcBGflSTwnB37fOLZE+4lYErseENM9KI1IgbDkDEeUBzDSBZ4r1jKENbeBu/6lG
5HPX14oCEdvhRBbABIS58RPgiCOh3OxlGl0BEZlet2qzDAGJqDKKEU4jP9Fd5vcyh+eqsqE6zak9
coVbNGCYvcGkwtIiTACJU2YFBJ8OCI58GDT/qkv41mXdkNlLMTShNYYGXvYsN48gDPmmj6ed3QpV
fZdCzxhQUmss3yl3Fx5HTvcTbbs+ZedZth/JBK/2VopgqRRImPpJxoMZjZkyloIzSNql6rv+pI8e
z7bqoF978b48ov0y3N6yxu0sb31sElpE6bqWt8G3jcJFEepRnn8AYON4L2/oKNyoRYrck4wbse4r
fwhWT93iZl4Y9vjNwZU7DHt9Fh9JQ0+ApB6roedSCxzcI8QQddi5RqJwn5UDpOQkjEIZUwI4+Nn8
QbxfaWI9+Ixatj6cW4rK5eyBVr85VVOMnZodELHoH7ewAmJWMxsGpEo1FNJIS8ZaQbMenGmg16/X
dFCVt6xTT/AcLgXb64sAw2W/u/7AoM+t8vYwCd2JE1phOfZD5MPIgWM1XnI7SHxYx3pdq6OtyFpF
5bvKGjwbUAz+hjUyNuP/bYb9iyMvPPicAhaZjR+rtMonrpulZ6uTEhZ5FUzWyHEUdBB8mYUM0EOh
Yv0uUV8YhKo0GpXLztfgL7EpnB4vVDGb/HbiVPuVWbNd/eBx3CQCEQYf3XXnVFlt+Fa0wtvDHsEq
R9RDWy/C94eM2MKIBGQlvrGD4icN6s5QEiMzrmcSBJvYlJVsiV/stIIOo3C1fs1JWUghSHwxsyIT
EkbPeKlZa0zVDHo5VOu6Bjm1jbvHXMU2zRUyNIVpPw92VM4BX6wMTtl8YLbwHeu5LA4gALNOyaeE
EXXQRHlKFb9noubVVKaYRAcb91uDw+IN11m4SdJcAOapCqgrjLSoq8+2ag3x5Q027xIcdrum+wKb
saiLtyyCHjALiNkH1IbmaoHFiGveGsZUdubxDAcMNbXb+DDw8+tl8Z3V7v057sByvbYPDDwYp1L3
7wb0twohxWOFIoFyxNr8gKQJmm0fsb11vYpcL1AyQelq6T/2vBQswD1qnW0zcQk7pkuZBAtjhgth
ljN4T4Z9Xzg5m+R2RDziJ2GfhJk8KOZTF4EnMBIQftsG02IFVls8iR2YhFukW59iys6yx/FnIxQf
Do3p9HmvqYkI7SDF4bhNYSzMt9l49ggv3mZqt2xqXrx/uJr+NguqiG0GADwROX6rkxpwXX7qj/0r
a9UKAXj5LJZGhexdv0afdYYf7pnck/q5CyF2MpiXZzUeyOqfW25QATcvT1EDkldhNMZAye99A09U
sYJ1ltmfw0LS8MunAQut216bovfkbPrpKBg0ZbKEoX18N/uIF7Y1+1FwTzRl5rWZKmRkd8URXG6N
F0wSe1rRhqM6Zi35eJFp+apmAXXsquvsmoZAPR62I/wd9wkMgN0RBJrsb5roPPmGCGll6CouQyBY
b4QeQ84AGL1PfpvkkN5/xwebQ2IYJXZ2h7QfY/fzwn8X7Y7veRCpHW5v79yw08JtJl/Q6JX50fi9
sTDt5wII1Ab0W4k+gCTWetzDa2JdPO54AMw6TEynIV3Y69p1+W5bmL7nZg1ro8Ka0TAGTJ2Xdfa4
1hUv6zicWUvp06gIGRMAElAtsXNfMV/MX+QgGT1p1PWiphLx6pv13EczNg0KjfvkCErSciAK8ga7
vx+yU3NWJEsq3Xcd+rgcBeoyYIBJ1Xc+bHv8QZrJeNkbSocRpXYO51q4+mAzoej+BnxBGgJaUKp5
uB8TrEQQQRb/Jg5E5RZXPlZVndXTViEffTjdK3ldkau5vW1K7+vezYweeRn32Qen6BkflssNTv7f
sSP0I9/YvhZ/6JKXx1AjWMIMDdbMpPMho1rvGSRtaPLWwWJxov+SeKLxralY5eyHFldqq78/ClR/
sg/ZBB+YGD8Pc4qfx8dOGRebI5kMnhzjHkXPQY2hFjLqdpOYFWZmi+en8j0WAJq982/GW28LbT0h
TBmgb7fJXTixwQ9ZH9nAAUA77kNPmpYlanMouhFffu5CH8pEzxNVTPP5r/wPw+PVjLZ3yJWoXK1Y
Tlnjempd+rQ4bFrsXGxr1DlTgUay8EFJd/YX7vez97FHDaMWnX9CrpTlj2ICIFE/5xgDSeTMroa2
Wzy3rTilrsKBpJixigPNhNeXIORIl7xYrQ7qEB4ir9pA1UtMa8ezG6Bl5XMInNLRnWpvXuSQTixz
jgLygXNmGJPqgTYKiJ3cJJKCC2tU3a0VL3TuHzhKH4iSAoLGINKvXwO/dzpYhZi3myoOxEbYUkqe
7NlkAB0jzCzRB8bE7m73ixdLFHdg3BzsjONsGQjeiYF+6N4/cIfiCoAAac41y46kyxM2XwLLeUCV
lZdNkiKjqie4G83iNPUtpheyk1oMnoZ1oU5UVFQG2Vn5V9cr2IbImoq8K78xdP7e+Fko5c/ZM2OJ
KRj872Yky8jvv2SrA0kUuQTJX8WD/N+ogWnDHd8CRocDAyAJqgHXnLEcF/sclRovnwIuBJnJSdYA
Xj8Spy+z3gYL+rVzpso7r5LpBe/DOeEFUM0lG4qLfFxs1Hv41V9fpk3indkM9K+4TSQxOKKFeqKG
nD3YP0iT4D+ZkNghY0Hp/5mzqhRFzwdhpd4GhJJUm7EFxNDmM9oKWqqGRDxAfVnw00Sor0PBT8US
CVBclj3rhWUnbSXFU+9Y0TpUinACsh6JBkWmZEgMvMot2rwD/27DyevS5yqYQzwaiHwLDbZmhwBA
wzYjGE7mrHprvdTh5nQ/8S0G+bDrWUD81yVaWP01hN6501KbyK3bh8ibcmeF3iTPYGKJgaOsB9vU
xYt9b3tm4U9F0HYRgkIv8hCpijPCbrq71ad+98/mwuovMKyvfuLM5U2ThplspbMA/A50dgLyT3Gr
m2TUEuaGyOSR/ES9jIXmR0UbArl4kuge6RGUT8CDaQB5GDgcb4p6BifQVSE9lEAwz4R91rvwBCpj
PgXICRxti4lv70KdWRb4ZnNfeohlE5y9vCy2qXhkNI4iVVKo8DYs1nps2SvU6g7tdRlxcr7j4TAK
z39cECvBR0DPpiq5WM9rYOD1bixPjIXtoXvXcP4m5e9NCQQiD3VAoctmp3jV4bXZdy6d9cGF9EmO
ClzTXMXSVvtUWWpvEYlRf9eUqIFhqZ55FNMo+y6dye7Bx2oHlxZSSF97bHny8qHLO1YmFBC4AO39
+oOYzzFLrw11zz0g13HFMoxJhxZNXdIPzNz5P4z5JtOy2Td72mEwDAvyoL8LTAm6UVSzJVIbVgjN
yth8kKdw7wPF2evta9W6RIdsDYDqHxYbsBJ6eiwP58rUhycgqz+k0o1p73YXdMdS/PHkBQoctDBx
GO978YyS+PoQBPw9fFHRskmnV3A16zg/scQu6PyjU7hibwOCvrK7UBAcIFZXMkZRiiaTXxyw9ffF
ilbOQBtmKmXEAhob01Xm13ngEmbZ5yi+PCbsG/rcOPc3oRStJj3fGEv13MkB351YWJFZjncaJ+7a
epuxUE4xrMf1MtzoGQjOUJC8M4mEOvgj+mazYgMPBSowt5wsJ4sPqvFx81ywU1tvlFmRebEAUn3T
aTz508MCWSLaOCUpaCsB9vTGSO3TC0haML7/QH3UjazBfcFtAmMPYHd+OWSAh9YfoH98DwXd5fbp
dl2X9BI3gEWG+M6uvo4V8IZbuQe9eDdl5YRb2YU0/zN+HPXDHpyMeQ91wpdMBF3aEcfpTdaF7b8f
ohmfdnlhSRHNhIgz0EbcEzhs8D/i1BtyJci4JlPbDYW4S7W7OZu7xDAVMNljlewoS/WXZMv/b4He
MwM9jtVnf0ZoDut5bJKcK4jKdqiGEIeKY3/p4MBpZEN4offseQVrb488PcwuQji691Xu8d4dbCPb
BF3yGA0Nl8e8QiWvexLr3i79wKhYHkpKFKRLTUYIn9Jtpmt+36LZjmCTHGnIolbwMxLpO8Lvao6H
GM7HV+6oF44LEoE3fCYRnUuBu8xjn3ffbRHU/Q11l4xqIcGixZOfKZh3AteHQzfYw6k6HkCgR2zI
EJnj/OddwqEHF2XLpUWnlsvemAjK9jwflUjPinJOmZ2PZvdPI4BJtBITOituU427/XuBdavJN/g2
Cr8xRSsZDeDP6TOLTzh4kLjnl7agRebAJjU9q3VfZXq9DzOsOkczQIft5cv6gwF6sbJw/Pa2XMm5
8s3ppHRm52cMTtJXSsClkheoaWs1zTHwLme2vAHdGlKhGNfY4Agk5GBHignkfwM5dVgYykP/bUEr
hKYXlai5T0GidCizZksF3jGZdi7SabBoulq1D4PnWr59lkoKfoYFht2MEvcMzLS4M3oUjWG2Szsw
prgrzcj6zSlqH0UAXAbQqIPm5qjAKh3KMWxhDh//v96dsft0Og6nTI91fnB6qV2Gy53ETvvkL9Xp
ol8xhVN4X2K2JrlJN+lTteXO1UUPujNrL2pnWBHfuDHv3LZmU/JMCHfk9p/8ad/SMM2TI+dmIumF
owV3fAJURv2HFbiG6iQLKkR9sDgWppc0eQMgKXSHArln+K7Hz2D1vhKEj6l3cIeRNlXX4L+a08Uh
+waMFY6HLvE/FdqCMuCFUcdDgbWDNRR5qbnnmYXgExNv5r3rcsA6yuBYoFqVeW312nL60ExpA8l1
m2r08RzB7sRySStgGSoOUWPuPm1GRU9eeRpZYeD2uZvunHg9oZQ1Z2oUpz0tugoDr5XtAGDdc8m6
DAdVbf96zPm17ao0XPKsJVVV1OlzsVL5hlbH2EdXBG6YjbAmfn8DmqZVgxezBZS6B+ZSsz3WzadM
mlk9YNl1/sCWn8F43ZQkEck4E0FBXSkcWB2Amm6nSzVeqjpkjBOo5MN5rKnZX2bxAviomWv0+Txf
503r0dEm0a5Da9ulprzb4BweEZzo9w1dBAVa1QRuVlinanqWlV6EB4CV6155/QKS9qdM95AoBo/s
j0vPgBnoYk1cPMn3j0hPQgy3ePOOES9TGfYpTPHhB5uAPB7OHT1atzmulHnf7H8jrLCcFgfPyMPS
TuQNql7ZviE1GS/WyOJfGRjzgm9GL16H7LbLYsKofCyETi3DKoZ9ndA1J2GC+652af0Fh35Jh1+o
eOrmpLR4gbsIfH9lbd391/LlM223NIhsf7jOGOWu6G7iBeTUtZvmmE20iNOt82VuoC48Tut44aMn
aST50v32QmYDmzRHmGsVuBfM/kH4qlTFqH5jPdropiDwWw38EZ4nV/wy6ImzTvGHQxPKSPZMS1/3
qM2UuUvq2yJ7iWwHbM4ZUNL6IjletPwUJSkMZRFrRx1O4FSymYtuq2I1pKEalVLzM2a243BRGlgA
a2/QIV+bOGOI5V7Npp2yxXY+uT39FCXfs87nPcBK3PW/eX3RrbcaUov82YtJsBZBzE4nEuA9NUrg
3GzYqyRCn3Q5rsHXl6PbgrmtRke5blj9SAIMID6GdxOkEikoa1w8Kh0vEqPTub9aLQsHSW5k2rvN
SyCEQlD3ciDg4K+Igb803C/sV3FmRwolOxdPHsFqYeTpedJvXS9RnDLkEGXwVqBESEJ/VWSgV81M
7G1XbymZjVEKYcMIR2yMh0AVf5yYYbCTXChVPPm9+V4PYglpEhXZinWb+NJSHt7P6aQeQuXB7w8w
IdqOP3NHiclV5Rl2e17VOzQ2gPkO/6SIBgV8QGIdz+m5Vvw65ZIaJDca7EOCSGG2LCU3toK/TIBi
3/wVaqTPH2oyUlNGJinNKKmBSkZSovMHepkpZdjbC/QgARGMnd4SrdbQEPbYVIK0rzJ/tS6zfI9a
VNq8Uo0CgKaP2BYUhNg4XEICugQBfmITHlR1V7eSyodyuqcxDhL80Lpt+lONGBSNouO/y3VEVPxb
nR7Cs1miZGWKoLVaLBXoBhNBfMv1ZxZygv6T2RcTW9MZLTvNGLcCubEgQP5K6zF/kthz9GjxWIFs
PSOoiIjTDoj7edYUhmYJQtHNlVsuhQL0VXguNIuSZBrP/zJPaTztVPGX8D1sXL2nvr7zlbdRulg8
idfRRGrUHDxlXkHJDdQ+usd7Wtav7rUTo5voUfJ8wz9ARFC2gIcnhuR0BWRgL8FAaCQhB4lz71jZ
7slcVOI8qEIs1YO2X8e+bvprof6rW64+kVpFDdmoRfVBdQnpeBRPrnZaOpeHS3HebUsASbsqO+Ge
JpVMpUb72q8MhIk1VSKTA2Wz9SZF8d0sSCmIJoK9UzUnV80i1erPT9B26ueAISk4b8M5Dm5PEs/v
D7e7RBOMRaddpcbhndci6sCWiR+a/Oz6aZ1iM4WVzPbTkytYaWztaXqtWEoxMWFcrinq77yn9org
vNaWyliJ6juGKywSxGNaXnCNGAwmx9P3Ab+Y2oESfTYDZ7m2iONoop9hxsmQDw9Mtv9GW74X5urL
Z0tufC8O3Kj1787lN64V7kmvRKyqFoI+KzHnJpRES1cEpY0hXQ2EZ+aXe+vEPwkXKNIEfMkerVnu
1Z7hrYeveHgX7fkAeAYIWMjqbE5m6mBIuX+am9LK7FLlP/ovHmGvaE3Hdv+NF60ANHNZtsCfSxsy
T2n1Ip+x+jBm5JMxbrA/g9YScGy8I//eHkgNMOiTloqxhKdfwU1DB8fjKlAXa0ORLmipcltT+yMt
kti7t62RzR3tU/Yt44BNy5Q5cuN3i4zDuFJlsNW4ssHev8EQg6wEcipu8D3YPX6P6DcCYjf13uAs
KnvZr4zvMJDeRfbDWPmugx8QmKdCdTjsXS018t+UnkTlya3vyzIVuPrmWWaUYUmo8nWrJzt4qYlD
DqwOFrdWnVTj6PintmuzYB7DJIrjDXpDPoO/abYqqpnjyOriuwvrLQPjAVhXmqNWoUXlz4jJuvmM
fIhVU/Y3vWBY3Ext8JzEvu9lli/k+hFK7G0VE3qwO/zQq9YyuYvMSt57sXs6aE7nWPo4LFM0gUcl
Tnykw7sVQ2zQ3mdBJl0w4jAX/4/6BJ36nTZrfWdvMGvPRTXXQ4EY3mGouclq9d7AiZjpP5uDzFjE
c/5MDyPavCrqNLxdB2xEGIuhpvd3R4bII/xTQYsxQrCNQ9TG5M2B6z/ypZf4CV9h6nj9cTl8uDb7
prRukUjJ5jewGiOGh8udt6HS11JuQocK0hLKXNq4Hc8ZJl1xXRISWFP6FUgHW4cU/UNjajsJwj6n
Sot4sfARU0OpNzqSQKAjPpVr+/0AWlLxmYAOV+B9DjWndhFCMBXJAkwJNmxrd9z84HXrOX9NbMha
YVbvRWeO5PkLu8ayaxbhJ1KRLL1+/Z2Kgmj2OfPAR6oYdMqRRuJluQ6qLCq6/r2BHS/n1eeHtj+D
urVsqFDZJ550Dw4wpFlJDVTWCKisBOqKnBVSrilsSUN8dEif1XN6Qt8UuQsX6p3Of9GuuOe2Qu78
3NyRNMiGTMr1guaVAJL0zC8Der3aUNzaz6JVjI3Eqszku/WrxPV56yCttCfKeiXEvkR3scwcCAqj
K1bvOkLo343fx74zQGFkahaaUy1oKT90SroZJyq2QZEwPm/MQb2kirtve2+pjPIIIgF97dzomQIj
3GibgbdYctzjjMS22LAgluXeLl3+OstMjLX/qfs8mDmC652HrvplDDzZqtBzYUauuIXWbdvSfEZb
wz+hjE57zLPZ8Br043uwsnlOWen3J6EiL54+Kz0cU2FfrZXOLDNvPiTm33cy6nyib7UpDxVzJrAK
6tQbYGKQUT5GQt81fSk6XggafR1LsMlQVPYNgZGmw1FKNG0oPan6zUxd1c9stQyvpErMH2wf2T1B
wt7uK9Pdzx9iFyoFR0K+RIFsVTWD219OI1zKKTOAOqDclD+DoLhmcKMU0nlZjy++CsstdgQfOxTb
gisSoYvB//SlpY6oFbqmKh4qG1SykCzSjHFCUKkuiEREGCiJDux2qHtTP5tv9eP+li6Ln90UT5Jz
B1ET4/joek6P90FQ7cbFlWXoMLIg0EPxe6OOVe5vWIgvZKsjvwm6Qww76fAMoMnPvf40jyAE9nIV
v0+7+Hep75aMNP6/0+a/H55fmiioiq7VRRwCPCxpZjElAlR7BBaxOoOFZm80JvVZYXhhBj1fYlA+
x7nelgMnfz86xNStpwmHCaj5OIcfcv9RM1+74oUxtWZpiy2+hS2c+B3pqxFesoO/ECAe9/gQw1Pa
exwqkDNallfCWnUX5mqqWDDkZ+hsPIFNndf/EgJAzjOHEMNLdJMGch8Qqxy4XQ8FXsfaXOiUe7Sf
u3TQQs1WBNW6uUFyt6884pQM40fYeCdBJKPPZgLKHIUvomtZ1FJCaeLpq/NGhMbXoCmlgDZI4JoL
AKxGx7x4YRqsqzfbz9q5s3qsglNpvtmioLyl0d5GeMdwP4NMu2ihi/qvy4SWqbN/LF2TB8A8gzMV
sQRhPAp/SVwZk/y/f4csxHTbcuCOrnTsHiU9e34uNsOa3KRkDAKfa+pyruKeqA+2OkC45bWprGav
XX6PcmgIpWFgQr36PfGhtIJLDS3ATpBJ8qYSpeC/X4+OjG1nL34VP2rxC0sKU6k5mcbeor9H/cQu
kT8cajg6KKfOFJFq9MBrCDXkeE3JlDe7qtvehNQIvKrwDbPMqEJVisDCUsjz+QmV9+mEexAQ0Nm1
aK8mkagXwL7chRDrCRkdrW1fj7ewMHNY0OmR3SfDi8Yi0UFt5J6fOwNExU4N6W5J6SU6VTCZ71hk
DsweCe1qqMQ6btu4j6tuNno/ZVbLAqNmlb6J2MRV+tWhZvTnsFNSM9wZ2Jild6PuNAIU3lQRhzS7
Y1gpvLtYUsmz2HBtD/OEcMXy3PIV1UeUIAWvSCG20sCJ7FzDMXfros4QE2XS7eaTRyzSbw/PaVDW
FBb+0oP0ijNz2uGYJFQrWKTTfLrwr4RuEClhtX3nDZnXb96BiVPB6VTxnnOpEAIeHld46dUkuXJ8
VgSiBNkhLSAeY460dWqVPdhie0QTdvsmj9rCEoalPkn2OTTBxwrC6UI+GcV6YGKJsKl1tHDNleDL
O/4wg1iwrBjpY4B/Qxt6yfMi9QRfV/89J0NpawGNVshrrFdA4l+svjId1pLldEoFZDjnGHkGfjDd
jQcIv7oevyCp2LbY9fZFdX0WvWJgEmyptfQYLc0CGZOlNYXGFb4NiHkP9rm3AdqfE6bNzY6u5qY3
43NsB0Ok32Zb4sLCmFHymCyvqgEeBtfrQR1z/L1Q2Mpa9nMXrypcoO8BYoy+CB4Rg+OEKi0crMWV
Szb9BSt1cE3Qo9tLflpicIRAlQMfZ1yMpHN8JvLTTXJxvHuM7O2zuj3c7XEM4iMpPOw2IgF23mma
+Q0HSqLE63M+/TbKwiRWQcv4tn7WaD8pZTsDLyh8Dug3SbZD3YBxqDz8xe5ksFcA+cMnaYB8UYbu
zUOSJeE2NhdQofzjeuX3VkwKPPNO5QNNWG6ZQLYqiGSg/ieXnQxTl2MJga3I8oMUoTLT6MLhVRtU
W6FSc3m3GIdv9YXs7O5Xi3NEPCLH6JsgZXBuvv4jGu4iywHTPGVMf9571HFUfxD2SOeg3EYBeRzU
9T/mupJUpXRntccVozLLAsLuZ8OubEuJsWki5iGTrnW+QHlVyFXnt+8TFnneXAjpZuQltyUMw98y
YSD7/lcMqYmcxwAD79unSpY0DiAYFSgGBonzX7X7IJN8IGTKJtGN9LMSCf29foF7Ew+hXDto/389
oSMFjlXCjrWhYzewoxB8dHL1ZfHzvvVuXuIjgZD+X0qf4VAXfRfElJ4qCjJFVMcYfXl2w6f33crk
/NPBQdNvJVNhlPIB+Qz1c47qlxjzL32z/MchIgRWn5ZAEbApcpxMulLQveNns/flyRhJgzlNhpOA
5p9yrPKGxfCnVouKAB4BheylhoqNGSODUATvMRiyjAIJAeaEK3FfJ8AMsFOnm5pBOrM01im/HIwi
2WeSNip3SsDEXqDgzWw12rG930IFvw36onyH6Jv4AAXzNeUuyNgijOP0mp/75IUDzyx1j4HpCf+7
cq/00cGfOO3ZutOAV0qkCcAk4f/u6QW7mOymBzPmOKoZpdhtYEXlNYGcwKHuQbophvRHGgegKbyJ
Gv7Pl7VdANCbOq3CuEXsLwp6XjhW4/g611/Tkqi01qb2g8x6+9QcShDTJ/GVbftqMCpvgZlvdg/h
2eUzGdjSQ+hETRQGaBDHJmiLwzi7qGnQmDsSLG3dthSRvNTPI9DPecvTrvpo/Cd3aIPcvtKd0TSc
mvqxJsMPbOsgi/tuXsfiS+nTvpGXML7wRaodCNFkvVWVDllTT0vivrXxJt0pScGKjStZ2VFP4RLV
yYlvPRPfokkZMMYqSz9imeAP0iDEZonhP7qej13oR17PAiq8OW51GxgydQnRjzCy5q2BLLMPHUVL
8fhO7+cSbstHoM1A/6rle+rxKAuyDzLdD9oPIJdv2YJOUMg11BoI2Laryo3xF6+ILxuTwDBDpwkR
lfD6Cc2u2TjbMaHhJizGNgHjZORTuXcXhzToIuGtJICQqL+y5D7FUdDsN/af1gz9dgt7t3cjhpYX
POMF/3ahvt2c3bCmgntECXWPvG89F4jfS4b257EDCJv0EZjf5kBr/+B6mAeOrvQL2rn6gVYb4Aal
5bKAWvSpS+MHVMHr+XeRrMgAcBC78m00tOSlrOnNQkh2PNNOEHTvz0VfikYyA/tcz24NFk9LtCIS
mWAkKVnG4sRxbaqETBPNo5zXK7AWML76FukPaGyXbiYuFzvk0fOjeWESzPco9xEme2D19PLp2GZ6
uTF4VBSEFfpVP4MosGqt4L4rw1wkR4eRXhPZ/k19IwBSUJ/dXJRvJMOEichMyMMLPvfS8SOEbCo/
vaonw6ftYKmMzZa+BvLBTr4/V6ButzePckzojcrTwTbdzg0ThyRFhaOHs293cAFrm+6k3QSQosFE
IZDqEGkvgeWSFiI7DK7k7AKeLrapVjdNswcsrAD3KUHUkplj6pCgdPq6LDAblIkozuumr48L2dmE
dU8mGtJT4T7eWfbg+ehNvOHtzSjSGCgwewj0FiokTcyYgxB9lgoOPRe0VdHPzTxz+mH27kdGxg54
WR3q46oVPW/6neJN8M8MFAprGTo8TPTTf0AO/uOk+qa148rtQ6wbEy3N8or/UGnIlvp1SbKZ38oi
exX1SacAMHD4NQ6h77s5HprAB3O9dcXNWVAK8Bto1U+Q15bXYQqAXuYMsE7KPmgfzsy1LhwiWY50
YLPZd8QToBsPrdi6w8xnW8XmslSe331hN4sugdcN1K49Bvlulg8QfxdMOKMLex9E83wD/TOCnPVx
SmqW3LCcC226egLVb0sqaHcwhuU4eNrul5lAi9EYMoOJUY3dT1YrSVtjOKLX+sL+H3n/shwRaLo2
WF222Rgs+TytOtrFXYpzqq/E5VkhaiRgHIhadgbGPbrDFL4o90xg/m9QW0K1oQ0X6niNWcNR5m9E
yjSlw1ntaepoD+OGA1EfmfqXL2T346py2QzMV+PJIeS4VKWlW7orfoo9mdwUN0WnnTVV7ZpFGVFh
O5zjErL1Xs26NSULhtdRmZAcxW39CBNlYro1HAb3zuazxSDdQLl8pl/wYkncrV0UXKSnSK8LHUn8
zbid7tIvcmvRfXa+BXiXemwADooXS1ycx1e8sBv+yu1GpsAWpWkBFD+oA1x/bWa+Y9SLGt1Wn9v9
ebSi4qW1PkR0aKLPL+YrSgS3z9lf7WvkKersxlavFA6TZn05VG9BL5SRqv2YDVusaAPZ6AxORw0q
kUP3o72TceBaSV8+m0jy1EdOVSo6dNlpK3oDWAjsi/OWDZGtMQ+mHTfsbq0zUXCYaImmPXyM4Mvw
ZIctYpevHTeTxspNbeCqyu+eHoPYRgHZHx0Kg0CYGXdqUjhwG5pmK56SS9K+dPC3Nkjq9VWCCJkr
b80gz2+mFNKwwW7Zi+P6cv7EY0UGPPVIXaMfKiwwV/J6PiMh6BL1U7EYRytXBIvchiYUude5mwli
YibHUHL7wHo9wjw+roOpMWPGlSV7z9qJOD4HMedAiCSkGdH0HV6HnHI0HSfNd6TUPRu3Lk6/XnJx
iuNDHAaS/T6ckWLvv6fzCsIkEnTjcWUtmwRsZiMQJA8ZON828XwYmH23YR5dP1FrN3zZUL4Bik8F
i+iY40D5/WouWndqpNNnAppYA+B2RkebDuL3khzAwMhphpLgLvaqA/liI67kZsDx61W07L7LuBMq
gdaoii5RDU+EEe4tqWlygAyENFLBJhFByNLIR2sfE6CLk2h3eQhWk3XUOBt1rySFC9aK6gwT6H8n
3J4t3OdhDCkjCK1QwOeLjYGwslemyELBAoNvjryeUFYfJP3lp3Pk5FPTnc3QgDUKoegD3Q67bZIe
olWhdsUAgumf/TCoBDNnspAkrz1bD7ev04CSdj++2mKxfTJH+hRX3UTUjyPaYcDH29VR1+2pBAeh
YDwBoBbnJABUQZtIGlhq1Nbfi0riasT7xhhNZA3ON3jQhl3OmoNSNNc5NidQhnSqdm5DOJG1E44b
4AHNkuTmA70rMwUQsyME2v4qBVoiSFa7B2zk2unSQZZd5A9KFxnIS1yF+oomLW4v859ogFvlc640
/YtgHiJ22OduMljOsdYhY8KKaZsc5kOQsCoFGm5QAHP7aqubInE69NVa8xXGc/3SfJmhmyNpUSIW
roUe1DoQeP6VJ++fFtaOcXDRj1V4ftkcpKm327zTcw+1S6zSCd0ogO8ADer6yFLYTSgTmOqZtfte
WG79RtlRb0o9kmsiurS9jwiwtBEP/Q7+5arz3Vqdpec88YrA0NIKXvFx2U19ciKeas5dVr72yYnH
5sC3BUS3sVV8TSrTGQ0mkJp8/dF3O9n4AnlQH5gfOy96MpUUPoqv3ML9go6NJlGcEAUq00vQ8ugt
yKlIdc9rmSbWDipi4Get3xIT7WXN324batkR/ywsKDtNSEsUD6Vib+3I8sNPzPXhSgaFjBsW9etF
UZ7PoU02nqvE7Xyf6vWCIVxkMBejQe+cvuRN2oSsR39fFQKRiN2C/xtSqpjIU8Pa+LsFs3FQ4pGN
4RpoXGjg79UND8qsOLaxajol3FIMeMpyjGlh5tKy1vgxIG4VD9jRbfHlwFjon22myZNvG5Cf+brJ
+UUXZcHUcwW2namQyww/MgzbFiSFyDMixl+/l0jtwHDA2RboRJ143Jwix3217c1LlRnn1VCdZ80Y
IHulGT4lKno7VbuAFfSDSvcVt61BZVWkAb4wS1ONYPzgCJ2anDlAlsEcT01ZVpQVNoH/Ktq1P0kN
/2G2QNSjwYcs61Jqyk/CZfTwToilAGWWNBPrYvs/ZIRW7SROiMrs4XGEqutKJ+UYOPT8FRgTtUpF
agvJQDFlQbnl/mRf1xx3RBQs4Wt/VFN/wnd4vrFohcszdLI1TE8gEnUNj6rFR6ZHotr/veq7qJue
eBLfe0UKaW9NtwejQ4+Q7x7jEonekvyjkUHSdw/yVC9CIz752ymP793gAWtBcYQScMA9H6bUYSRj
T9sb6rnnr3K8sjMAnMdOca5Yy7KOWWelcIRtWUAneg4T4U09ooOHxACtAAExHDOfkh7qI+EQht3B
rRCJOi8MyCnohk9YCqTdMM0oJd2mkeflNcvq1Fmmv+Tyh+bPvtX7UdLow8TxG5tEv85Id1beQucY
UHortaX4iWdADOdadZEtzO+dsQyh+MEhgoYWoF6MQfw4hV+Eo+dFKFVwE5v02v+CVRIZole2sXVQ
6zLn9Yqw9J+dpGXG+1yhuQ5co0egEEthyQ/8I2q9nn35CnlN9P7FVfintvYJ3ewC3EqD51l6QDQH
tTGdp/ruFetoU1p+JiJwCaiYUMigSuDKYTgnC36/gdgd0hN+ZvhhAmcsMbs9PUb9OQ4ETi4C666O
nLVULocGccR8VO5Z3bufAmD3vTW47kkMZDn/KxoWeAdoUGrSKGoOkM7C32+PE5cROjGND0ADzJ77
Hee9phrJVkb7JWgdm/57VJjES9gAhuWWoHzbgVDFhc1PaZ0fVOsiDMmx+JsJ3wnb359VkhgXWosG
2PZ9ehx9K+mXiO20X2fpo3Bh1ylwhlW00N9xKgPFfnMWry4p5DhkFBGRXtv7QfCI8Yw0SS2TNpc4
A/ifqaHASilvoznpeS3e2SL3tXFxSxjkGcDOdSLxRyv+oRsnycyfIxVOZQnowEqQJvoeFGd4TMfs
MnmXFkwBBeCYv3UNcbasWPSnVbgo5r1r2HLZDzPWaIjvDAlHvQe969x3T50DD1YwcKVmz3/LuICv
vdyJv2ZZUY+E10bOg8PIWg8pYZYAHiMKmelaQQ0UVPtjwjODu1YRGpzmmor3dbUqgp6Yv9Um/LTi
RrK4nYSRthcSIvQpT4j5dR6w9hTYCgHLZPOiZjJbjKyXfoZxRmBJTsnRqYTnWtbu+aPFVSaetZS8
4v21LILWfAQBG0fdrPocKPQcrpWUX8UD7CkdhK/p8NGxvtDh3hsAWVTNgiTV/Q/N8Z20qjL3fCja
FpF/Q+iSc5WjraIZtOrjflDH7H4ms+efFiG91Oeftrw8FrhrePa8A3lp5ofugMxH4cVlDRwfXdbB
KQJx1wvrKsAHLkqZ0nPX9Q+7Jk7Ta63PKo9lSQNfhMSopUhvR4HmhfvAO9rOUVNdaTQpZRmtxy7A
yiQL1SIPtTEfnz5+pQb/5eSdTTAcVuFWV3W9pZBRaCsfHXZS5AiWCDoCldwiP35lbAOz1bhFHp9K
/SkGVZ8n3yNkW0VZYRn8jFexwDmof8w9sZCSRgNshUBGNi8uI5YNBWzv1lxL7V4cS1A6Y/xW2f5X
+U0bVVIY96QvGmAXxzdfdwVsmjo8fcApEc6hInvQqRrk+ouloOeC3qI3I4OPoMLfEQact6GAS2w9
ni4llMgfikrXu6OGhviuIj/CKMBcg7kfbadQwgiBZ8+9uznPEDOKj4r9EJkGP1vD6y8hcNEKkV1b
xXshEsRGJLeUvNH+njnMu/nYSM5V2ac50mrAcTpVohBxkZhVXz9LuN3y5locumJKyEw6tjOdx8g5
9ifJ330K2mxFdYPYQoXi9zKbY2msF0Rv4TolI/QgCVqdCJj46DruTw4VeUr58d2bTBZqEfz/GY+4
cYGuIlXXBfBRldau6D35YbOgROGYz9LU/9RkoYAhXTLFVYXjsmb6a0PaNjnEUCDfuj3JdTtmKnBI
8rSGJZlgLOxdJ8JkTuuJUODjFE2C95so2KVIMLXrVoACs5tn8nMxEkgwF4LE7VKSajo7DqT6PjS2
sU09mAhWzdYiX3MV79B00v7Ju5CXAyIjL+MYL3YmZqpbq7FRbHW4j/VZgaLmK/vw9lVsuRx2VduE
0V9xIzXpDBX2bkWzEUDciIP1xSDfh02Aw2mMBHK0uGVg/US2VWrx2y8CkA4CYCvZhayjCtp0n8Dq
qibWr0O2iHljIDX0e2EAQf/+HnhJvDAo2F/oBHTVMf+GNvkhniwSch2asAwiwX/cd3i6cXJLsuEX
NZRKCBAGgdh5wkqJwKRZf8GI5c6fHNCxWOSZVI4kDEGScCjRZy7cQUTy1gREpou7jg8BLFTAAKBM
E1MTNRJhsnoj7DUMrKYc38n7iviEEqGZxabPcwV6lyU5LdUS1K0iRRCXDoGKnEVtibrOdrHG+age
EkwK3YuB8awJbIFI8rrf0OHp/3X9RIlfNVzyR5eAx1HVJmcFhZ0IaXuSC2fDuiX1qstL1CglI0zm
aaHss0ZRkTqEFFBoHo7p4jeAd6yWor1M3FZ9ySd+aCNsVO/kGBPomk3u1nKX2ZYkm+cKFBhpKKOq
nP6ugN43s6hy3mdOCHquWpBQNDlbrVim/UynmcWB+UOsdbgmnyJlTbgm8hUu4N7Kn8+KebJEjZkC
e93rmccrSoV7Gc26XPgK74l6jmFfCPZUfTYwYo+8Mry/7hFD23TyZubKbt0PM+0s3P168h8wauve
mjmxQ2dA2as4lrfSbdsNj8iIs/lP6i/fStaBuSm6vupK8OAelknd3bnRzal9+wwOv6Dv/kAcGCKF
mWvq1oWkiRLdulpkwCYIPvK5a0ZFWwFQcdmROBPq93dk4tZOnTOyjb6BemeWBt5jxQrCI8gjtQ/6
04qm0FgJ/OFuZxuJQudEj6enKKYN9GwT6kaLwCaIg8aQT9ImMoUgK9XV8PardPP7b2OPqmsJ6GIz
i+Q2vaA9e7Pk/shhujmi9F+mIH4uq2tcV9ebHVPpdm+zGph1ZaVYIxmCR7Q5SIbGGV6N3rbBBb3d
oGSu0S1YxxFah+kUgJEfT966juWu4oScJrcDiabMNUiRfxusaVKlPdGfXQjVPV2VIKerKTfqIcVC
Om2y+1ZzJoEzbXTvLzmoAUNg9UpoM6gNPpYMd5bYKZWyEBV0NuIoU0O2E7rTg2E7X8aIlnBtK5zH
wMHYB7TvVV3jL/kd34ipdQz0a+QRQwHvDM+EQpEmcK7S2OIj+8wrHd4/POfL5N2LPkuj5Lhpaz9w
ykK696P681FbUeZ5m+lTRIa2ew24Ncz6J4PMcvFWkQxRk3g0qrV1xXL9R1TTo3guFqrgAzkBnrzh
XMpVlsqNrv1g8Je6AP0KQfBbCZYaD3o+fqXw42p31iKG+Ef1UwWrpuQ+i7weOFJCzH4XJra1zp7z
aIMHaLuDNpHuX2Ri5CrVOqo3T1UEaU3/KRhlaoAppn7gmFbke4B0tKr0O3/dEB2fYqHdDjY3+Xh4
UVgsXqqhKexFWXSi557xmOVVAavCYiTRcQR2U46X83r0y0uVSp/cHDSmOaDDIB2Ats7L6kZ1JIT5
kS3Fv4GnVomOGvswb7M8ufVqL/BNVtLiaT4eywz9xlMqlf05yghVIAtjo0OVW+cLPtezgap2LxKj
FtTmPrA0XG0pL8fO9XOu7XDsQIcSslr8ytwJWRJDfWvRalbGdzmFucX+nWZAMKl8Eaxt3n6i328T
jcxEkJs8P6VK2/snH9FHDsqkesMs668zko1ybeuhr3sTualDKWOnxsNoWiGzccH3t599ui6/8vR3
qQKg7mGGN1cBU81i9EulY8bpWHBUDYnrCwXIwoYk5mggTEEQ86HJbr/g2gRkX2glYbeu90wCci+B
tnFMAxm/LaeaAIKRoq1aNWUIjCfNRaNBPxZuWpNbPHbqJL2bzZ47j7UaTcu8L8RpS1dbQxrNyugC
YVJDSIj4d8+OI+nlUXCeT0zcG9r6D4ff/gtmf7Zq0Nx6l5YfwAFBA88gUvyezISCPC6CSGUAZEOE
8Lu7n3rJ5RrV4YP6B8uWlOTZgs72QyNDP8+FRwydjQroem5h89kgYCvt/rem0PN66vcLYjYWq2C3
OH3AxJDGyVXESk7NHuFKFHOAY+/SRUdHThe+hhIS8+5GbKvYMrbJ50KG+6ACvwjY7JXvFP1Yl/8n
5/OqqEHa2i133NnrjcJk//FU/Rle0uqoad6Pna8IuOzBSTTRRYwamenekt+gqaPhEVr1hYJHQowI
7AxF61KBCENz/j4c8x8MUUH70i4gyOHClN0LUSpu3SfySsqTBBciEYe7rXjKHqUPWo2BWdEm6Hth
qBRMIw+l0b49zBuUBbkYOMIYg45iw8CcgBZx7zPGr++HwuXDlUMXUEjNTcT6sERfkqsn8fxptti3
VUzJNfsVP4kbsY/g7TnkFAZsM3pn0KSXPTFlSrFMzFMsGjYfpTjeJ113L4aEofFzgy8/dsw8JlGQ
+aBOkKRmR6G8RQ+jpK+OtYynw3OSq9JIN1Gwu1ZxhFjl9WSmq/p+OpV6G+lbsGM3IgSeQtYR01X+
PNQhBZlvDbcsutafu8RPbsC8ijo+8uraqQZlappQp5GjG27MPDUUJ5O2caNDrZjQDyMMib2JeFVt
jE5+CpwyNLL2aDm4KoH98i+fHVCHmcsX1DNXORB2cDUCuOEVsm5wXr6pdQwOAWxQVYAzRW0hKMdl
0345kp6D8B8+vUUlflv2wxIgSYqanDNZZqnfExYIyo2lc6j7qrZnDI6LyyJxQ2ciTIodCiloEmJc
YJHe6fs24PWo2QQLRkQBlrCKXtjyocj/Ju92l6eq+zgiIINsxYajBBgFPeEavvFgl8u3xzgTsM5x
aQgitG2cQqcmEPdBU1XamPt7MjaJn9DZlrdy/HOf7ShWSpNcZnnd0MZ0sGA6vHHZjXlcAXCKZ2r3
kCLHYBYhBC9LzwGq8Ae3SMup/O/+Lau9SNSUwrVXdQ1edzNXF+sA9dGuU0fmLNfBvbY4Rg/RV0x4
dA48unik8iZm1tNFfrJ2WWVJyL8LH9x1MtCt+5E3AF8rpyYhh5xiHryXIeI+4CDSmYK1zzCmXrOf
0ROb3tSPCC4z5DKKL003zS09qzyfu8lAOrUVw4qhIOVW5lwcO3hoAJhknPrZy3W31uidrc4b3E45
+QjqNU2jvfIMWEXbeUPvelmkUzV5EoksBXSJhpQofWgQ/JBC51BcAS7ObMDp8Zzqc8MGrM8HNCnK
Xe1vvYI/1o9Mn6SW6q3Q7wWFwa3d+fF+ISdEkNd4iDYr9vugK2NCA92voFtzp8NZBk/kkawfXgVh
DYIdmaCqRqu7EhAIYxWSQgNLeOlgXlvA2p1b/6fd1hVS6V975bwRcoW3Cb7hQSjT/X7YRm7A6SCP
2nyMwjFI9cTT1HTRhOe21+ykEZySh4KGKP9JD7NQJUA3JP0f+2T/yiNeUYDsCD5nJXL/cwVgQ9TP
tPgx8k+b1iLygnWj/6Z0aQ+ELJvq9wb2dYJBYX43QZnMPDk/7LggsUTUb3QAl7GFSGzwNzh5IDbb
Zknd3DCwnhevtv9RzPOXz6RwVQ8pWZBNs9LIczo5s75JguM/AEsa+LWGAqGDfEM9jk37ZIFeq/x6
ZlOZIJ775WccIbK16aVK5lSSg54gCmCzmuv5MC2Q+l1u7p+VCB03Y24Dk2WWJhGI82vNghZN3bkk
7ctOBfHpV+xgdGiZBpH+94dPaRa4xh7zyVI+OPaIPB1pScvR1Br0XtHWO0IbQ1xPJZZAvFw2BnXu
hiOjc4SimAX30p7EKoH7gfb+vZ7yeGHyUyUXhI6A3wLHke6ToD0grrXMdcvzJP4MHENRoi+JnPnn
Wy2frNi/44pQaAG1uTx0Yk2chXDzpDU0sWPk4RJ1SL9ZfOWImSLHPAg6mLna/idkJ6H/1g8lJtVD
mOQ76Db/2CXTnyr7rmmDM2x6f2E2ai+HHRr3EioQ1Z6p5+bFx43QcrKmZpRlo6w3+QVJ8RQiDD1q
z6B/JzRhWPZK+4a1M7GGNk01Hv5s3Hpy/mX8cMO/K/6BuEw43KgxiBKbTmwJAf6exCRFp2HAyOzh
CgJ8bv3wF/pOwo9ACTEnusyF0ZN+JIoDdrckwDYm0yf6LEGQvvpjfRX6OtU6sgxi+6yRHNDQrcBm
bqjlxpMIM61LECKOgwBJMz8n/tf7qXhjEhA04egL9G9OXztb6t9rl0G7ktSNRbK3lUQi5BW+zewE
4eDvmg+zWEVZfksOcwKrdF3TJkqI4YXOLHm2jK9jdX66p4tcYqz4C6fP/V8U1YwT5qsAAkIg6ee+
isefaET1NBdBBLl+Q3o0sR2SLsa+W6ZFukQjTHmaf0cZFbdejKTXlwdqf0LSCUrUjLyeTJRMA92r
q2IsUYzOarw+eaf6iV9DDKWvrsBcgYIblxnEdUx5liKG6xtVHlfV9voHsqi2CpHEtDlI3sDijSqk
gvsyLxZi70kgTLKkfWWqSzZYS2SSqi5eEFiXJ5wVbPN4t3qVXKB39CGfVfvl7KF0yd2XtyOTezb5
AH54KDlXwQGw6YwheqR5N9AMiViCA/EQHvn3g4D89R1oT+gIWnzfSUp4IVFsBOULDr9XCaoVKxbe
e8Cq5avAOAdGu9478ZWVnSVt70xqBXegWEOrdMe2/lPLJ7TLTYMy2e2qQ7T1akr4B9wJVuZvF5oB
AH1q57Hourj7iSHdOrCliDyPkoDqes0PfRAskW41bM6t5oLH5ZKKkFh6rq756a0M/PNCnIqLpiM/
uKYml6Oj+NeGc/8fFlMhNPUqqspTYk70m5M92jlgPjxulAUna7wQ6KKopTkkoysT8KR27N7l3JIR
AW8mKnrZzvF++nQXNijSTG5y3JaRkZvbL+PnQpSK2URW8LmVHCS7cL5gVsSjZbPVRtig3rFNW4vx
72P4FPiY38lzaj59PvEQq3lx1ZTA5DAGReA1zxqii/98RWjvUi68w4781yaY6nwjRGVWbDyIMawJ
pkIn8xNzMgRY4gD1miujdXXoeCcZt4TRddkuf1AAxdGpYuSy7WU0Yx7I4cqisXnu37ny4F/Eux1M
TIvkXcUsYa6B//xxpmP7DuPJqwz12fBEN4gWahmxkYWc30/bmA4GGWytKfRfQdKBsyx11teC1J/h
QuPJjtDHgfmJmRyTAvVZJDS97qQly5yiapmP+bgxDDQqms9bm2mTDL3M6SVHDFfw8AbfVDTpZCn4
IC5RRjjb7saFvwvt+9NCV5cjq1YtCTMMlemaRkgq20m4BSK7oVxbngfn1L6WuqjdDkSas5hoCO+5
u0Qhp8kVgNKFkPCGez1sfuM5lJVfF6qDOv3S+222RNoAL8cdlqwdlBlDRaca3D8qoqGpIVZ4dQiG
Thg8tWPYEVk/HbXd7/gapP+71p8qgYY4zaBZ2q8AJ7EuyM1gFT14xPcoo4D29a8L9X2hWljM2MlF
okSdsfdNWZ/XvT2cr1cLB990KX6Fo7IWZyxFzHTXMhc4tMFwE6BRdzJaMpjmGHuZTAODWril5nrq
fi8LLYhQw270lQ2Gv+dkxAaLaeOEwcB7t6S8tMvnbWHxh/EXP4prLbypnpSxygem9SDoWV6hjWjJ
rH7sQFsSabmgZMXFPLyPrAYh8dBJ0DCwnx4V4POfLvEyIpwJwV2oivCOFGk0KVPoUz5/otKrdjEK
L45/9obbkX2VoH5tfaFxPG+figGLAgEg/ZZIpuBW3PYtNa29/TttQDedgyL9QFYQBy1UKKdJceTV
9bz6dz2DLSZ2VGVXLLyLuWpNyUg6U6/7VBB76/CO6Iv3H+XcF4JyMXFitWDw4M8cBDon3iUHWiIb
+qVVuKmRR9SSW0XrBIXYUZ2Ca+BKB7x53+1gnVoYrW/KuMkRsC9Aj6/2uhGHGdDi3KIU7GrUEEyl
cwA/Um04sl96zGEyT9bWWMy36LNrjs1lQwjrB1tQCZ6bz7+ayKWxeStzIuZCkdjmVSVKR4+wNJQ4
VoCbC20QI2egkGAYV5Og8V/llS+UnESdmHve8zjdBXGN4y0B4/WYHl5iPBoKWIDIu6wR5AsB0ej+
PTpt/93783CTx+wAZiNTgPM3hqL4PzwHtGyFhrroMOsnuR2Bqx7om7Z/YBJqzGAFJhDMIo6X/b9q
ut/Yi8FHtm/7iOGNXTlFQxlyKsooLFBWNz0i33V38H5VrYI/qr004TLJ4eOvB8f8CDic0zDrSWNq
S8xQpYcL/RudEX8a+CY3wgPToGKBBH30ojGaZCt+3SZsK9MUiSJS2MOn7Ub+mX2MK8zyX7Rer/M0
AX7cHBL4iFVtID3SXlvAXsHj3yBqTDCuBLYxlP76oqhZKxxQ+hdyvGPyDA2MpqcvY6KQdyhvm1Hz
c2jVuEQRQi1kz5ZoC/E0T7K9cqYe1+mEWSXeNpCEpeo2aZSzMdMvwEKJqDL8U0nVOindltplMxmb
IEuDH5oT1+IlgC6W5TlCwLjK33hMfrXNamIgOdYMJeJcfQVIJpuw0sPUumSRI0LWUv+Ti7V7k3X1
VcBFgZEZBQCoCNvDMJs68AHfbQhyuZgwC2jv/icgtEwevZmBPm8IO8uGb3KeWC3pLndbMxmmpYty
YuU6rHoU11JztyfzGJwLjIz/25MDzfwG/B6Epgz1elM9hqLvNJqqHSRGtO9KFe/rmNxCZbslL1g5
xpcZLZFIIPaoyMsF0LBQB4G9mtvoJQc1c9Hoqi8g+E/RqzZmUwpR2r/hzoeq+Wol98QMuOpwFxZG
nEG318YsviRd3fEp4JFJ9UQ/MJ0d6jy8U2loeekQ+qG3DnEMMDlJr3bZXrgc9bhKjqkaQWL+SXwx
2dZ74qaj/eCLMijuMGhMLBWwVHAgGIcF0lcVPAw3m9E2QzQDy842p0CmaUX7KJ2z4IwdJWlVJ9lj
PteYXPr8vBrQoqt/dLPdMqaaIBP+MxFc+ya0f09jjLbsYTyt525uG7mL7qsEwmtq1wNeBnsf4Uif
zTUc7DVEz70UTpfzpfpmbjgGGzVK8HetnhHRgIUL8WRVy7vOFYlPaNR5VFnGxzgSleI1feaOdC8X
Wvw1glqxPVMA4bbSbENvS3wwvygzJRi714O515AOAsoLNW2h5YSLg2Jz5feJ4BEooFm/E0vLoytp
vid/w+aC32TKvcZnoWACEeD0Pf9iW5e2tcXHbeAGM9SvRZDlFFQcAptEpJPHWt/l8dXecaLfqp3+
kdl2/4MUhy6DFiBWMp2YEoR1vI8H7Dk2nwD7TXQCYSlM7oHpVmRla1M99HtgSwX833NPgJI8J3/K
Xp61z+rtizge5HFEt2lXkvV9TmIdHn8SsyXAIVBoLqT1dfg1E/Q8DA4/a+p56XILoSb51BkDUY4M
487EnwYj/UDpNZ3Y7SyML11iwDUyEH4ZyfT19yP7laHImsl73BpknnqZGADA+wG6qlTehnbicPOn
8PFsS/ezusFLjiHWOAOw4JJg7tpb2LuRChZ7AG+rZWc8QRy3FPnXItvrRKEX9HKwlFI6onOF8clu
FU4f4mnNNtatTusmKm9pDq5XrEiu02qXwi1MNe7tH9rbXFvdfJ1uSgqxyYHcxqTE0xpKhbmuLMY8
PWdDZIO/kuacSzWUUujzqN0rfsvuG/z5oRaOTx/auuhei/R4yM2uGXHPNRvyc0m735X9h1mrJ0rD
IZxGuU+yLZEGNai0hoV0ybOTei7zA6tgqqS+u/hXLvdimnmC9eHSpxtMxJ1YGhAv5ECcjoOIV7m/
2OvCHfZW63LrYwIEXfkuEC8Q6VCEdbrIoSueetcX2UD8XAyotS8EIpNfKUi9xSJ3MoClXDp2uRDa
pqsv7I1dntqIEHrEIsB/tdVLwH18jhmTwF3aqIIa+vvl2TsbD4PwDp8S/Svd2iBbUjJ9b3RISlEH
TanSJH9jbA6lWJ54QP2cDXIXtVr4y9HIBSE4xsseBLJyDW9OuD7M48TfM4jQUfH7YDCMYnxfner0
G+Q66bX0IEqbjk5ERZ7UfYY5xa80Ak7ExReBfEUK7GteoulSOVdGtWOAITcd8ledj24lpYiaoRUR
h/TMCJc4PV878WYoLYJ8e/7kx0ua31j5YUam+E1sXc0UIxlc9DewaXOeGTI60A6IDAeS22RaOoSf
o1Sme/e/+t8ETK/G+XomWSlepzBodgtbhHhgP56A9rfh7rj5HI8sCi99i3/CPCoa0NWy3Hogr9Rb
YxMhArzqJJ039vQHUYBQ8pKej9TCk82Y+JExUGVsZG7FtwVJM9OOPyxM7s8Wcacd70rZBkzgzoMz
Q3Owv+nLJfzM3+nnYsFURxaf6KxGsANCGnk8tdx62ZrknzIjz485YoOgDMSOxJ4N2aB+UN/gpNAB
4OA/wGAZMl5OXW6sPZnEJtuUNB1/rAulE+J5606T36nCDacur6JKzT1vvO3xTt1/2u+h2O8bwgJ+
8TI28oiGrSWfKovb48FQAdUqDwxFxHqTNPbytn8G1Xv88/0Wg1ORoN4GP/ztAwTJGkQ7BgexIAQz
CGJzOMQzyylUkX+H/2CxxppBsuueolJ9oiUtUz3IebWtE2Cc3qy7BoZruSJ2PlCfvjbAfVK1w45F
k2uOKfDtVNTqazjYANhlxPVxiac+FEqFnKzMy/Qkf2eD6lyZ+jqsseCuAZtdMJbKFu9icm1Semou
Zs5V4kqsGqbq39ZO4tfiiW3gEUGoK69T5J/fwWCe2MsT3wCHceGEzzb1e/dMsVxDntabG8Erqon3
3+RyjZdgdIbX+JSc9NJ3rKttzxDkPofFlkqqP5BNpsWQv028GNEPRrsvbW08+Klj+Hu6KM114UyQ
izu6MQMozq+AfDuds2IkoReFV+MAmqQw8HNZoGI31XB79omLxhKrB7T5uVZoGiirsY04pGI1xPpI
PO1Yws9XHmP3MD+2IhpmB5AzXUMNEHLckTY3NaTjS4++ZoaZhAf/H/R2m81XKg/ydcjTmL4U6s5b
BPCTctLtPVYTDPU93MStjfThY1iW43t7HNJqzERycoJGT739M/7pNuxEb05Ama4Cix5hMVKg8sPx
uvnfapCHjnz1H5HFIjCI4L13cSe2r8Jj8FBqDgNCJEQG7et2/1mE+m5/C06Yd7i+5MVltbza8vyX
PZs+CbUS9zAYxZ7xyrgpwpP/DSi0E6067nnVaGl7noA2oApq0ZC4bf/XFw7iOEpHArW9q+9hXehj
Tbpsl0W9mki+aWIz8nL1GSUIzWhmgDWLmAmPElp7Gpgv0QERLJ3dDbnxc/FtQIPqXUDNQ3l9mEFS
ZwcS0ZK0z8ZyeC4XZPcM9S+pFINP0JkjaYE0rKP/hkxoKks10WTv8EdlEXQe0fqSd4xZ5f7gAv3O
p/85c0GDI0H6FEmzQs/9VBWoPK6kHnc+cTgiUh43A8mifjFW1f5BETGEmQQnMwEHkFNE16p9xuFR
KThMjHcTOZMLJOIDgEYW8ZIrsXe3d4i0WZ7fq0kwnFyibPHjDFWcGEM/NNKGcY8qExazeoWMOZ9H
asbv6MJxkenAilL7ZDAiACiAabMAgv/FroiwI3dkdLokWKunC4xAK66UY3PCOxnQTC2izQivtHK/
nFkE6+NNSzKyyJGjqWZP4JwvbS06Y70lDUwRPOZpfXY16qBDBWL1XrTMvAWXpxFHOl1YeHng8X2r
YjDCoKsCHNdMR8RbrWOPADkD93fxj8FRqJOcIEL5Nbq6RoB23REufMbCuAtNEwhnp0ePfwK5o4nn
UEzRrJAYlUq4p3JzI/7JnC87lkbB01A3N/kQIBQxNftM9rQYsWCjFh+rIrRr4pe/DziPUBtVL00+
rMJCxAl/s2Oqml0+HTA0AJwGwq2rWo2GF6U9GvcyJOawuOtQewOKRdDfpuDRxyDtdca2PdpDAXo6
z+epiIGGZNVEjjNho7NOBTY/bS+aJ72u7hvYgzPI5/BO4GWG3ZFye00opxIeT/bFxjzBy2js1hX6
j1hnyTHITtdkC2ru8+Iv5lHPggK/qy8yzAXm0FEmVI6d0JV6Jw5wa85cVEHbeBBG02NOBPR+Rq7k
4hvBi44jqOXnf14lLJgFEsVL/HgMNyWNqQxQW8tme/igEn2o6EoxQvmNsnV4aR3Y2RTavLNkV7rF
/TdqPKpyh32at1htKgTxynnLU/aFwdJ8sX5GH79rsX+p8jiJHunVxv4coLtGaKUleszfTLLHVqVb
F/nHbqxRkEJ1B42lwiUswQtV1m29KvHf3BmgA3HV1g3oobhzYZfJZLQ5UZKm2cO42Gj2L7LTzXtm
t8xm88QP1RerDaH97TeuWfWkC5bWj8sQudOKvtMWCuCAg3Npaufn1sdOz/NodpI1RIP1PlURCRko
Rz3xTFtuAj+hArZnchHP2v+kOS5nQia47gTJDAwftfEG+C/ubpeq5AupJF365G5yyVH4wl2wYNpC
GzeC+i5T3ByTSytHUt2mPWgIGIeA4sioHZJyyqLOCpU5xbfOMmUqegQgQda243GbXP49RKf+K4Hm
1RYCKf67+4M7J3TkOLNiyr12+hO9O/aRqoHDISUFUB6N0nLMqh8yYtnL/K7tTpxytoqf5tEh1mGO
IISEAM6CJDeGEcLPsW/BTbuubkFw61rUf0i5Rej3PpzzC+3H+98lojMjLG8agbemyPZAPRw6zSqe
RP5fk5emaCtCiib1KdMkgrYvd1XurMHj0eOHABpxHNUwPo5WjTyktqipqIJ6Hd2ISHt7evVwqCqA
+GVg2OCIVast3JhqYHycuipbQcdRx9KqWQcp76qp8wZOH/DpG1Vv9jND+MyZiC8+z+Rxcnx6ydzs
N4qdrASwgoLPUaMD6pPg0lzYL87vwTJ2cVLjRPo2ugNWwecuTWNFuTJ5sSxjSI5owqJE4XQHrfo4
NRv9jyuKlSXJlwWPVLBL0baaQh5zD/brW+EFyzIndYCLCNlqbwVFdu/jwxPhXQXSu8jxDucm/S4U
AFz4VjKeGfEAPK5e+rs9ILS1tfVHVNy/EIG20/kA+WrxCBy6OgWUj5ibA5XeMCT8vjYt8X6DfELv
3k27YS2ss5Q6eANt6GsD3yLeEGKYy9XkADP5poA0xWeWvAyiEQ0H63DoXaeD3G+5SJdUGinSmfcZ
hNBTlgl8kzx3M0BbG3quYUOKdQ84s2eCi5exyQWbpmBoo41wrT9uqI5b3IdGTy6h3GOOw+06nPh2
b+606EdJKzLyfKLEVLdCIANx+7mXZQO3bmGKUg+59rtA2zCQox/XA26kYVg/+nKlLUZpETiu8GOC
OIXMk7T8+OQY6ZNWi/Es+fIqWrIf5hVVGE7m5Vd/0kWPT6a5y9EoHiJNlSKX35cif1ux8ZU65/+1
UZTfjPRUrdY6Jc2DbQffo7XLeBawAnzemrjehn0IYY7uTqciO0I7PDJcG8VL0fJJUAz2nPPBmXCU
tp11t6Y+pNVJJLJ5Lf7tck1wqThvn2XFOqpReQ9COi7csTUKjfGE0u3PIjjzd1LE8uqDbqpMa9Qd
PJfVihT2MM9BegLvcqWMV8kHCixJlPrhb/e83BAScvT7K6/q2eV2XOKwWyubb0mSWipprKOH7VVd
4J6S4j0K5EgNSbx1AXQH7EpyDowTW34iKMU6D4XAL6CQeBarcLwGljow/rORrZB4meQRx8TQyoFv
8INU9Jmg1II6MldnS+iltgdc2Vg0q0qia8gN5KkmTcnp+T3XLxyqVPQQo5vYM9l9E242Yw+Tj1Cc
7HY0QM12wtu3yS1x13pEw5FkKKmWjhRYq0jDQGd88SAi6i9P+u0FLtvZQ9Yk+BjPj5jCbxxAKN7v
UySphCqAv71SpDDNYFn1fT1/2lAs2dI/yuT59aqzYlfHtRxTMLynHqSTiIwa+h0LgIoiXG5ng0aI
u+m7PsQgBDc1OoAgE0zJkCVWkznss1TwMUdL7yg9N7sWLmK4wY6CB2BnwVk7UWobdidtfJW1X023
o8MdF1XSFLapYOt6N9qiQDeLbK+jcPyuDakXj8GGhE115BuFeny85wO2xVD+AoP8Stf0OwNA0C5u
weoh9T86oAYSG/vWDB5TK1mQB1Rl9qKRelXn0c2UDsUfMbi9nzk+1Z+EMeW7NVIbo7cqUmUhyL5m
1VyOcALEvssvElPK3NatBVDNW8KJNWxs1KLtEEmOpuzv49DIQg9/AbhNdm94WL/pdwXPuzaanHP9
9NaiGQ0nhHwMdTvj2l4FpfXsRZFxzWlLW3Oj4OybVycddSWPSyFTarIRCfHrPe3ikxEEseoqnp0i
OogFwwbKq3sq0hXw+OltK2/MSpDz3V5k9oUZI7fJbK7P8EurZJ1fHpigQFnCyJyb6BTY+kiZuaR/
5CC+LJRY0pIy7ieBjNkj/Y8Z+2e+LJedYPtDNoOEL4Lu4LBuJYCYi94nvpANPMgx2+0Cl3mdo0Tr
2T6WNseo2cA6R7yZ/CYKfH7CJFjJtND4pMd3jkxPZQzjLSFAubglbHwU7YhsRDRD56oVrUuL/anc
mntKIBtcy/DG0Rybg55JNUzEDqR69FdOL7uAozz1efXQRW8TUDo8VIIgjtpnz8Sdh2ADmGheat7W
GXaUky2ARvLQMrWJP/fGbEgFvR9Qr6NgZ5odp1CG1vxCuqVAzvHCekt7GvBapCc/IkrZGrzaw+ws
K/Q0QEv8ZoF+E3rf7dhvMH7fsTTyS/s0w6h9GC7ravhYhwHdofUMd2gjUa1sANKthK3a1ndrW3tT
gtnvKivJWS/WG3eryga4bREZ8DV01BkRoJp5uQqYCy5e+rROSpTBTpiXCGctp4PYvBvJnvpPG0Xm
0i9NFaJiueBji8MbTwZS/uDmkFMVx5VgYlOXTz9ZAYs7gupQZEt8dqYgIRlkKIGv7/tk4qybIM27
YwT+yVq7DWj/YfEIpFyPNUq6Kpuu/9SkyuAFiuaZBM7InoeKa26NVEt0+axkY/ytSBnwzHQeVvex
2UK4BEwpGuvQGLtdnJrsj+HJjnriRULC2DLiDhYRAJkiduMPsZoY6rhP1tZwaUSZf4Z8ghwThyEA
XE1jGGL5uzYJLIbiWC9sC484e8P5g10aqVKabA/EMM2yPuk13vSpPTaoUAbYRCuxy6xaHihK7IDD
rSJFQT6IaLvPCZtIm8m3uHV+/Kw7CqrCcapP6UbrHn5O1Kvy4dg3WFNfH9IQYL5mAAZUsw2CPNIq
xwel6DccFFyo0IJR4rK4fA/8HCIyeA4ln+l9nGhyICqt/GpEvSOhLocAmtkpBVu13R7iPOy5+5Ph
KHH6QU/ngRiZmjYWXIipRr+lrR4ScOrClCMyPVaDmsiYcOsCajmrzw1SGf2ocxWz2FPfZk6PeiO7
wLKKLu3AXmRPkwsJH0a9pbVDg/yDdUCms4p9AjsORL+mT2MFLuhgo9Hn/muEvKOtrXV/imN7tXJT
0ndJKctQAI67OhzqWmCdbcoTikLYqlbXCKbSU+e9kBrG/+f1c716URwGPJmpZr8xRiObDCDxjEbc
wxHQG/ar1HLQujD4U/WNQt5OS94EEDYLjbYNM9qPuinyAReu6RI8rDQ1ymBL4rmjOVI09L+nUGX5
3tKCo4PzmswYyqvI/65QyadC3I1pipojos+6LCOHfKHENEh4eXIYzmrR8YO+gpg05KQMhgszrsEl
8vdErxO8FZZFTNiJKML2eflg075wzVX3ndQ/dH0888VhEQ+LONjtumXAFMwe804//S5sC8WbEefR
83MojaWaNbjacQV+a3b3qBvtClQTWad32k4ph9OVEOKh6XNLOHLaGQ/T/w0IMc4NyGuonQShFnFu
atGAoncJEVMRVbZe2OF67S6o2bXPki/koD/B7SvrjDANT9oezVjaIWLlc9JR3ubcNGQKMRZvNLeR
ADot0xBYw2sq+OZrZS4LC/7wwZvuc4LzS8uzhlALLP+sax1TqrYt/PaezRW3Ze7+1XQSFZkVDIzF
HDHmR9SQYw0mUyNGGh5Hqd9gnezNRDj8myKmbhwewLZjC8VTAKgREsjuFH8jt5Wf/JCO2Gvxt2uU
QbBHPvMzHmaJSUpDoNty7kEEm30KmYpEBIeeDIUxPAdY3UhZfcMhAZfcqCW2l6tsGxHz3JtSxN9z
jNx+2PM4ujMbvyWim8pBsb3EJegxjXY+Lh7Ufud1B/AQZ+h3adu2lup69SMwcncnHPVIo9YWBhg+
jt4E/NnrjBKCbL70V2qW0Of8ro8rLtLGWcPstehMBxTl/VnQo9FCcEJYWu7O1ahD9x39H63l5CcK
dqGS+Rkpz1I4eUYdfj/9c6ujJIguVxGqwI9d2R0KZbvfkBM1KWqt+besfB413tG9KLaScBKG37/Y
h11GcanzonT9jN1E9MnArmb1dpJf3QOQIn2Yu09zI+qW7mubMjeV4t8yE//fKsdIqw1hnB8u9Jzi
c/pPLXIFdq+pWo1rnYfAcLwsJiLgmnIHC3qVELKKdr8ZF6+8oYx6b/fFh8elNnA8ToTVqSeg1PDx
4TAdybsYmD6oSfuXTsncHS8pgmsDSRpPUWdxpXeU8tamSPkwGLI2NdABvDQvrGR7enOAMduPmmhl
NXbHsIaJjyus6/Jp62V5xn0TN34PNLzwMxSFKZdleE6x5UpuGmHMK2Z0bif8bvcvPdY5zRkjU4/J
ayOdFQplNWWtaGtj08PxQM7jMYk+I+VzRj8obJh6p3yEZroAMbyOTkFNeet6GmAHeFu5mzceO1Lq
bX65XdTBET7/SSOazoOtV+QUzCw0xrfg0iqCQz8rGo2ygfsfVVBHvPwgtMxg1SSHEiRThMnN5N4k
IvieaFCqX6oMjRqRPMMwQIJ8ojaX6w1LTA31F9tYOSJvSjnXnbg+AQjbjypiExY50Oy2h+jT9zIc
DoiydCbPXExaS5NfmYcF3Kn2v5zS8OHJb1ja5Ijuwc/cUH/MDm2Iil2cWfpKX9a33O3TiSgULl74
lwLdgLmqmN6mEXZhnLksAEKGkqHNOQMwLsVX9IEZirsoRHyFZIxn/km0arc/n8122Kbt1hzRcvGa
92SC/vlrxWpdrTDIYd68Cth9vH8vFXbrVIvF59rSYENsTsaqWrGGzpV33AcTSsrorMCvcK7Vmeb6
xsbBl7QZU4DuJZFdxlXaX49sRdLN0KCjnb5PaYpoqxowjiIjJjuanOGjF4K3FJInaqFjf6yBQ9pY
rA0y+FaRrGry/M+7gK8p8XpeeO3C7cG4oBlR/MrAaez0s13Gs8B4/T8Dk/qW+rDS255uZGQyypti
FtbmbQUizzXGeUfutnW1Xyp3L7LHeW/SG7fNliXvO18I9k57HixExJo1eIG7fkngyqXqgoLugOb8
pbj6vHqXmjZ9KkXnBQhHHpOdDh80m5ap3WZ6PfuqS+dtOEICFEk3vSFZo8v6iTuMT8R/nfOXwSDt
78x9zuIVWW2fPEGi5fm5nK9Z8uwFTC1HjPvxfT/cE9K69OPqGQVZf1UpILir5EtIfIa8kRhcs2/b
as8wHqpQ3Bvw+wWSFix6IbIrm6SjbT3DyhUEZTCYU6f4rOxW2pxy3sVjRE+SBoxYZhzhcTVVHt5h
CmXtQLFYfLh5tqxIDVQTcVJsf/uHDKIn+D3lpwe84VcdzvAY3o52UFi2V2zHd4VrOW6fRkyZR3Bz
aPXi3XKAg49cuJShGORxv2ALDaxnsXtgY0aLT24Kov7XWDSp3SdZ/AoH7wNGCNYdPIuZvzIAwyws
abzOzh3kUnl2TO+1vT0nJFrRfasQwnH7RdhrkSufk2MJMXUdsFA7fBsyinp+iTh2GP947vuKxrdc
XGgM2PwT9Td9a54HRGRrAcIiz4O4sVc5IPsUgMR1lDv/Cb9/3N8W786jk1tLurTMEUbheXus0yYt
79hM8zP9+i6fQmWv3GWMCNiFG44T9rZK9XWrSdQRL1aq5ebJv2bhllnvK3iIqOrtznrJJFB10exs
p9K2fMW7TSv0p3trRTypoRGyFA5kRTTnvnso1KZOKkbirqCNVYXZeSDMtD1azOP/TNfbu05vG65e
12XA4oLI5inY1piNc0O2SvfjuefEs/IZHfkVPmrobuHnLjnVPv7loUFbegHj98i15fiLnikflBmY
mr+wPmQ9cusbxL8lh+FLmxZqaZ4fCAPQS+s07wIuQv1t/kQiYdYvy6mwETHs/QZhP9OwRXMXM3Wl
p+j1BnJtgycimQwwkV0UfKzYeqWCuq9Ja2nBeQZkkbP+xWE6A6wPAi+mfHQ/LxzHSngmG94dKHDm
WJ1MOy/JRF3R6jtiZgL9C4n4WDoQuRMy0XSFKuaIzMkole7IrnaMhTvbcP5ZDdIrtrlvo1nH3b1C
RVNgLZJHP2Rt9ApZL1rf4quCKAhtmJP8mmleYAdJ7GPILBpf2gWCRkIlko+p9kcPJIG47AsYmWdm
ZuiuDACslhhZxow452ubIAA/GD1s6ltDi8IwfcWoiJYXqD2n+4q9Dt3YHL7MDkth+8AHe6rcIk1k
7AGO0zG0e8Xb00bPXqoZE21nREF6Ck0voCIJDaihPw+P8hcf/a6x6Eo6qgFGoydQ07U+eXGm3EjS
/28uZLDRg1XUmtESJGxIVFKTv0aIRpeJlsQBjfmVdl3Uk1Kr9OW5bO1tdEE3OP6+mdYlmpemOGoo
GIoBBoDzo8tlp+EOzjFMi9K5HG9OvWMzxCH16akIr8DhFcTnMJ5aNI1vx+dl/ZfVq8i+SEseJPED
6ogW39lqoStr77UWam1brhDGUtSiRZDFz6BuQplbaQr88Q6Ezbv2eostidD1WTBJ/p7mDWu1sU30
87aE0w/lgCuy55Mh/eEf8FToDjlWwtVIysGLeqaSfzmYbIqUpQi9lmi2tU6kbk+cRZKFcVFNlo3j
s/wCMD9y2/D8GDfStBmFyQ/+JrEC1kV3ktYbAShvaj/Htj/EyTvnwY0hB+OtSx6CyaMy1Mgdur/r
kCck6W6MdLvZx6MFmxWQhvBYxrm168CvBRnyR0lSu848eZ5j+dNTKX8JT1glgbZsRACcdzCXG4aE
hfc+SSEzzeYmgNsq0eq+60K3KTlXVBoPKW+HOs9r4hb5y9JUeLm+GSCpmTpJh89kPdFv8Zi7Ah1P
+s08DGEZN9Dn3CE6EZGl0RlIe9NsbtQkTg6BqUCo9T+QRuDryskOkeziUkCpwJ/axjygYI32U93E
sinITxgI1d0i2QcXshTFhsMjW/TRGfqvYEo/9wgbnRNv9O5RelWOOpsEg/apLz/v2RqZBEL+eTK8
cfY7fxZDfa7h2c0zAUd/wPkjuzVuxyHxgVJFjZmC8HOyz0Vl7z4pEZgqgnYvh9gfrllArgTTKf0p
r3ouAV5mI7apWgwTdZIzdJWFxEg1aGoSin/xJ+6BwyFg21t2hXqJ+0fAs1Ra0uSX4XdPG2x7rVDx
gKVdWG7k1HsP/RFHbIpaW/yDdnV2+rdbCtHBd72oI5rfpG1PJbYaGti9y2qdkjbaSkmKbH2SysP3
Kf9iHfjh3IlnRcABFrrzlIQEZHbpyr8rKwMtwconosZf/muPh41DrO4ZIelOTviGaGXP1rIHIjwk
+f0RNUpaS+hLwUR1lQsW5vmk/pGzfhqfobPUVJ9RQ3n/nzL7RAq5uWL8rouwAxcRvNMwcE7L0QvB
iWejOt4sRTGAEgbOZ2SJI+GpINJt/7wMm8xCdAceTa1nYC0XoMJ2nBajwfr6AD3He3UBsbBU5h/B
2f470ZOu7+GiSFE2YXZbUqNecEFgmKL8cKb5up6ok1a3eDKlLNBxAv7umYS2Mxt6NMxnroOmeXsU
pY0Qq+bb47p4kr05Z9BE/T2w/ZHIt0B5dZBkR7OHljIEAYjUy4CqGxqJqXS8CP3eMXN0w2kcLiMY
csPHq48rDMBAXglxo7iXYLmTvIVEz2HOjrUuMbEtXzCDdKV/cuQfOddrHHcZXfWfn24xIqbVouYp
kZYGAr2Kgozc2tPtYhcuHNcVKi0ts33FK0slyzQhpGlGTjapBaKzYikFdMGiEOwd81Nd6mYWCXs1
6u9FBDam5PATIlZAjjLhkoN+2SuLMLXQ6l+IH0heyeQM1k88Oz3GgAdrrmnQh4jfCYoAVvOdKTbK
F1QeZeRwobGq51nZy1twK1LmGFI6u6F/0MwI9X1J/9gaG6z5FD4VzcZ0qO8MZxXl5UP/yD6Cxu/s
CBDZLtrchMNS/NrCyYumYsVhfOR5YW8xzeVZ3jtKbMG2fBBqszcphVYjZsg3V7Uq2zxTO6tB/74d
RVsg/u274AKX32CEMUr7Ke4YmWcqBd5FGxoIjOe65dwYho9kEQACDXdrpJvtVgapiWGQSHCBzi+X
iN2qqt+FQb1vtn63KsO3gIrZi02vMiIOeoi1DV8JEnuYnGqvYStZFR3NpjhBnq745xeHFiVmhCCz
urTxH/dAjp0TWGuidBMWcqxFKGBtBwXQWgWDAL0CKsCBVxwk1cysTzB6/zXZwz6MY+z8GNRMf836
vybL2SvcngVtY5pKrgIXjBPQZaS+aCknWk8X1yN4yzt9l5Kb7Ht/u4cJnZk1Ay5sgz8ajRy4hfEV
y2oRpiqhptUK8UUmjE8V/Xi6LvFYvnAqOChb9kfVXB9bA9P/PnfW/fTASIjh3BlzLGHK5ZGUQZuC
HqMY2XZ+crKQQ6cEq1ODPy8i03g/nOEQlJabBn0EYIq76ThoqSyBFNBQLjKRRl9J91RkZgfT2ZcX
zmzkriRZBNT2MtN6FtaLxDlREge/isRBk60hoQsWBCik7z3KyemnH4P4fGWrPL6gXGI4qg87igx4
CDf74PwD0VNlohFEH+iTaIah2AQR+uCKojj/TvQl4fdAgkoiZXxibXBwIZIhC54Qn6beezT88kYd
pVzGbaRPePJUqVjA7R4nTcQXeoJjVL2/uPXEolh6f4oDGgmmSn9IfYvcpFBm8N/3sMgmAKQgASGU
sv6erYTClWVpg+cux1aI/hB81m2qZV6XvTTaBohAhGh/XGFDmk6fDWZjvgdXn9n79pmY5lstEfgS
XK8San/QIJFfL7fRCn0SuLpRzSETOYYIgaJ6rsVzZpp8eKysfwn9fRyNLqrXQp7SZTSK1KklvxjA
W7v2ZxSJLhROYoWvN3xiXkx7KnFv7/gfoKqR0OXYgejC4mz0fsecwhzdn45RBf306jTWuSfCqCFS
MCa1I+eO163bnZ3FNF+g/jwa0WUvYAGDAl/WGfvJXlAPFqDVRNumI3EMkmO/CFR2xR7LHxDpgjZr
NJ63stTfhnIzeUeh0ThLf+tg8Q2b7bKliF/gfQI+vEXdIjZhyv1p+QI/fSJjCBwQDI9itftwbYa4
TlN3KRrOCkha5mmpAlqD89Tfr62FQXLnhMaXFu5+LDblANa5eb1OlwvZF0xazHoC4Sh3tKa1pfZH
E4mgaKnE/VlCZU8OdSVDw0saoI2TKjGNLDBn4E1og1S1Ch2SY3A0DlBflqjxeuHB9z7zxpox8iPe
uvkwGuJUdVFVvJ6iSH5Gu/2Zsn+QhnwGZwTIn+HpygNoGdgtM39tJBPZvU9cNJfSwb6LR/IChl+x
g7/CKZwEROvaGQav+5sJHtL1SOox3o3EgoYHmNj3PLVtCnqNpNyLlT3xhZg45M+jjsrE+0BV/vQR
v9+XG5CjdfnFLnQWZcNbiS9eOM6orEHp6tVEhbdF7/Q+COh1s4uPYl5JMttC9/9MwxFyQB0J301v
WMeZOK7djBUe0rbVEvJjVDj+xq+tfSAS+8gMqFsuwmTS4gSADhYDVAtxoUImrSKcpH6mYojZ0XOv
zQh5VTBwxajfAm7rJmIofwC4vwYibpUNx4LQm47oiAKTpc4fsPKwlfYeG2skdf/l1lxEirOciMwS
G6VRpZ0saPHLiVoXxJ59IeJb+E7L+SlFP9/AAUHETEOEAmMlwyaVzFDKwTjjoLtTVCnnxOh6zeJx
pL5ht2Na1z/Enn2HjmkZQuE5BuL7fLBIxxYvX93Y6vp8g3wQriUCuJ6tK3BqvZwByDng6d+ZjBz7
3OqKxu+P7j1BUkVCNufqcGFnv2oaYoOvVQbeuMk5WgFgMJeeJ5jBqgeK4bMtzWZ5Q9aa/HBVS/ge
2KhS3Y5WtTkXbV1xNigociAbBw/uGtNIWYvy1r5t3/INQ3V9UHPu2rbLHZp5jq0qNO5yGrMjVrQT
u4eamzS9mnNwqWgduCCvyXlKEkq0putGUyBYEeYg464urrX+xrY/CqYWe7F7quFUmr84oXFjjlc/
5CcE9c5Ci17aRk0pQtahgiIlhVt+x3qvy8I387f1MVfTRBjQzTqxhlKB2CZFii7T1QA8lewi+DP3
ZguIsICxc2Dh1ftkttr25Bh7GZTie3nZbG2mnwGZXQYA8W/pky2UkBYlXssi9yboJnuHH1oTWrzg
UV07UkSxLefoeGELhO037ct51kHTyxeRkBzpEVC+mZc9Gb1G9VcP8GYiE6pkx/Q2/wMkbzlpQv8q
oPLM2u4QIQ1tsD4aErODRGqIa1hY6EJS21yppUwa6+f8JBgpNF4/bAd1zsI8vYZGnR1Bk2+1PFdI
zfQqRMYr09+bcPmCF4LFBDC6mOvfB2Z3BKQu52mCtp1rqRLXdzy1VBwXkLsRd25xKvuEDPLlJzr6
/v6IAYPquePzUOEIDeGtEjuqo3APhFUj+kbimdm95SHDgOMZAAcIzG6sptEIwPTnmwjosU3DHkHM
C2PCjAg7KobP0MufDaGpgGTaXr5amV8cVhhq83XkNdC4ZDWIe6xHkdQwZyDY/bg61PICo/04NN6z
vxHJNMnTpFbMuFWZqHtcXbm7gaFBiUnNEr11EAHOikBm+4BFuV7v0FxosvQILYhM2f9gm3Q0U/w6
sXO6JCc301PdQjTjQp+8R3Ac0H0+bJZiCPkNS8YoJGDschA1wPrMixdXx3g3vkyGQjoPe1PYp+lR
RY4QlVzV6X/F0ZEeel6JFeUnvX9YW+8uNl2HlVEils0mhaiLkauWmCCAHu9HZPuQ8yT3sqTQisxP
j7reV8sxm1m9OHOSVo3LWhdHcCysupLeYLPVTkOzwt6VFVSVogVh8ei//cQM6cifS5J+ZkJ7kmOc
2uyf+Oylafev2LAnUXrH7c0eED8w01Yhqo7gMV3pFagGVaLeW0ifttEH1xkyigrih85wMCsQ+BRJ
6wIDyZIAgnjHLm8RuM//bhlcg78lP81ipZRSBufKVY59gUcbo3Ii+dkK3SIZLPw5LR7wly+D+ZQx
K33VmWsTdYzR2fT6YfMI7CQ/8vrVsDuZB5kzLeoNzynF3eOLMqoKZcMvpiv/kygFvfhVuEsmye58
0OvSaIxaWo9eATIiDaoNRu17B8OT2cUTctIQib6S1KJXlH6xR60ic19UEmsCPf08kdNMgUlEohV5
U3iTx7WrM4J4Hc9xZts1WZuUOhrcVW47cHYPy4y/8JPE2BiaFcN1k3qzduKwWc5ZpmGHyVUo+tWT
AkfH1U+gw4ElER+6sZ//VIAHqa1BIc4IDnsxTevb6oJqFVRdkB9x688oQGiIRR/kcCUamiUB3WSD
6iObeOvfOzSwm+1RIcrI63cNouSnnqKLVxdPLlp48kQZo0lh3OJQfpe1JEPncmF2xO8g7cxdX6EB
xjk5nrVhpiGG5mPkJaM0vB5OM/VieHvj7tueBUWOtPV1YjuZTSz6zbjGFZYEz2EqXucEA8JQS+Qn
Cw2zcc4amZVe5KZ/cjhK+AKfrW291EUEWZ2nhqdWZV5iC1wb6kvL9wS6IiP0LgVPvkQc3IOxece6
qfCUcITiZEhwBZND++wlZpDFATuDwZ8QJl/TJO85Q50XaoNjUHAJRjt9galR0GRZLashQNRwfAgF
zbYGmdQ8w7vI+EjbLxc4WElDwgNGGNSnWybBtkCYL4kb+AOqhVcdeibhlkBU40v3xvEaVCMkmUhh
7tP5xOBrfUzM8iEPM3LJE8gi7o8xYCLoEGit3lxrB8t/NjourfULgBbh2/C7kLWjZ8aFSDsibwUo
oI04TGDvi4bY7Gmzv0N8Mk95WB3Q9mHTFue87rVbSEP7UgJqvjU5HfQBTRjWFM+0NxerwUEERodK
bQYQmaFji8bIDECt2QTInqyO3AuAkDD7+OPnzp9Zkcn/UxBpcwo9pIQS95Jggid7xx337bpbJII7
hyTJNJvZ5hY9tPqAFXywLrWXKxTncgvP6R/EPXQiU5+Suv+UD9qYsR/8CgiOSQ3LGjLZd02+Ndf0
/rcsFmPiX39CRj5x1oVufMUSE7poTpU0inAWb8Jlzj15fXdvKa8NV/yYLirsS7KoZ2Ys3MfZQbBx
TtNapuUCoxrITzH7j3olQEnxGxeTqAfq3ORyQlyCDPvmJLWrYG4sNiuO2W275g/dBGp3LKvXJJTy
4P+Th0AP5HRoKEu6cWzvxbekOEAJlgM4QAxa1nVLhTTA3RCJTzrE0VXNM77sD63mSsYd57JcXTig
ucJjjO1f9dxl2H8vLjgZdJydP3A7gOGQ+TUrsy9cqFW71dmPRzwJ84YYJkchj+PjFDNm8R/z4a+z
l2wmYv/nyukY6CtmS100wMdIsRhQJSr85WGBjebgMQEO+Y9BDBlGeX/Lo0kAv4l9v3X/V26jtkOq
bs8pH8+TLvadQz3uDOq4OJ8VQ7MRzXGw21tQrUe8QdEubKZzMXj1bxUp7g2SBQt6VlS7W+EYe/cR
6w6auHBxctdlcaOZq5BPLrejI/05Dj8rEmjBWvV9T+2NHV8brSkuoOL/nVVLrMJYNecdl4o0VwFL
MSPH4lf7EysgoYzyM+tsmsl68VpyVftI2MrFDop2rJO7R5fMhKcFeNMAhZuI33FkRo6TgKtEnEkx
UkdCS832ZBYbaIrxFXEpLM5Wexp8RQtIdgP3KVBSnr/bk1dmpnU2DCV2zycyMQU4daaXKJks9Czr
p2VuUxckH8Xct9GFFK/JDD4449Qo67oAFcszK0KWu/rVr4fCLqfwBRt/KmVnqBxC8+6Wd5O2LINC
Fz9bz+Rhx6reYN1Pv8emjgt6ml+lYAJ/4DSOO7loB9bXN4sDLAjE8AlQBeP+cxt9KPZW09eNYxgv
AKnIZt7Be9L6NXcOiUgDsJv0cCP2KI3IB7j+wZdVPemRrdYVW/xkwlEtlNZH2egv4Yt6iOPoghiJ
lpphkGS2Y5Qy3HXuT4bcXOn/DK2wFFARrBJgx26P8pva26xKFlAJ2PTKbOjuX8cgPSVmdLLT9Hro
lcKww7i0S0Sy1snAsMqj8cH/qgtygRPLhOR1HV5W188Dvef7VmVmGqYQ1Ly2ciXrkj8F3AAURNf9
xhu+6HT1N51c78xI+WP0wiGlti1/VD5Q8wY1CcOrl3p1UaZUE+DDPRPJz2lZGvm04fkxIiinhccF
k9AHBsY3w5cWgnmb7cUifpqaAZAsZf+yek5cwkysKIWdGsMeAiX5uskE6McFyTQPJLHF+Imi0owb
LIunItu7kKc5SWTsFwd1FdsClLCHTUFdxgdkVFDlZwi7dmgCKg7Ht2PbT7A/1U4SxOx6shKlu0tc
Y2a6cX6WDO3jf6eDA9lghwr99DlDfINS1Dgr6CY6V7sWdOnmfB4qRvSilX6WHo5sIw3EkyS7Lmgj
vc0XersR2mxGQIRavtFHakTMrenPIqGJakLv/mlhJ6ux/b9pMmMpBRjD0eu+kTkyXBtMP3osmAZ2
zavYgTtuHZfnUeRrhEdMKSgFC0/k4fJ7uFTzQyjJgqtCsQQJ7zYnfy8WrQ/GpR2gnWhPd3ZzzDQK
8Mczc60tX+oZyFec8zTNQY0msJbMqlS8kF+QaTxTWRDe9B3dfLUKSO5yw68lVinx4nGSiVJm7a3S
IdAoK3NnHlaJsrYXApWVCBPnNdvu+2OGeAbKN4di6zM4X/4UZ8lu7rU8KrJooF5hKzflWwDbc0PB
Kfb/RK1M8cVTZkEXE7LP+na3EY5CPp3670tw1/Os+rIosdqXsXApdPe+HUfo8km5KsWS+ccW3e7y
9TR8evecSj0UGQA4450Uv1+YU9GmSsI7QT3ghjOQIdvgjukihg4BNPeVI8rJjaspWbnMnrc+bUNn
mYXPCYEw1LeZfOKn4YdZIPBGKneAp+VWQjg3gtGfYR0cRQmNsFFGou6OwUpB1RzU0pAZUwi+mvOS
6Y4mZMkDnCLwyCmaIzMGSV9pEifkh7xg0CEd9flfNxv2XLmTqGLzOBNLr/6LvDtELfaBtiPanU8M
ZwVmTomgFA1ZreCJh4wnTyI2iFyHbpzG5Xlkyn8A190Hb/2MzNeeC9FniDlG45k/ySZ7JepqFrJp
O6WXl++l5yWHpbAJDqXafRXCFOVWC1Om90+mAP7XNQBJP8kaPOOaUZhaL/2HDi+ljDAS9bUTAOrK
50chEwNDpNzd7sOBeoKDw6J5rRBAqeKalFMQXdoFBWSq1R5gyqcsMIHSlDuew8ic7AlYSsa9dZbX
VLDsHZvLqBu4dBtjxdBM/dTxv140DdL42bgpno00cCvPgfn3Fqz+GD4GukUMEriEmvkzWsUh0R7R
d8H5SqUYz/CBZMpoI2RzgIogaNMdhdwaj7o0+BuBDaatGE7yfWmcXxBkXip0TnqZ/hVlOSeUYfZF
Jzm7AIsYM1MHp3lwQDc/zKmOrYEMjG+wi8YtBjODqv/TiK6e/s246R+hfq25wrWzfIaug13BDyzy
P0w2zoDokqg/dqUy02v0cCC5fS2CcYlnHLUX8uHKSV+0LvR3eXxwxdCn2uP3fC1K0shsmW9G8eIq
XQtKzyjH0az+IBwH/648y6S6HkQzuQNIHpzw1FxeuDARPG3ykF6/qkCbrsaqTiHHW1f+PD/koMTc
r1fbuYxobt4Wh8ghCoHLCQZxjsKvQX37AhTR4D55d1qIrXWqpOZjlsWKY7huTZOPXrNaSO+68VTF
+DhnM1c6665CDE725UxC66QU+0ycWAN5ETRYI3sFIH4L5LntfNdvGFIrfHTDURN/X84qRpri6h5S
5/16pU4rVdtPwbrdZuT1rE16qxtf/YR7arWLFItG7nDUEeCfejbwC+yKtoP7zNHVgQY7ersBnEbW
2Cdp3p9LiEXeaBfxQXeSdgODDNtpgzM1p2EapEfVaW3m06Kl0WiLvzpMmGbgzsFOPVfJjjmrtfwh
IljPXGq+epDdrWszRuNUSLYVu8BdzMxPRrxK3zcZZzQn5B0RQg4BFJm974iHEAQwAGg8iQcCVuVa
M5DIjRDl5YlUPQaMzK+L71BxZQcUgGS93216+5b6B2Xq4uu6apFsf7ocDx00aD4muPMyoGm3kyJ5
JaTfQYbWcVZ8Ke+fJN8J3SSLvHh7gd54HG90gD6L5T6AWY9B5LIJzCXV6j4zr52xVkT1Mh8TFQ7A
m1qJLpeleudnIz32zvXxqfWls05nDXGzI9dqhtD6Kn+apSAqOMSytnX42J7ARtT4bEr5psjzx7+z
kZoBaBJiFRbo3KTbrd0zyf6VxZcmBX44mdzCd1WU29JKhWEFRmogG7n933HR8/q+gtRs/PacA/Fk
bQNxtUMGbXuHk+TUEYfAFgoG8MBeSnorWwBk30XAm2k3K/6l9jkhXh8e5qpOYY7n/B3mYum65tzG
PBMEhPzbc3gT7iYhsM9dK0DcHonrOpxDYiIHYBxllnzsHCECD8r/S9b9tSwuXJmX4j3GuyRj7fNy
M3FYC9ao9EkfLeZPj94SV4UdMcwPy6dZPnvi9EoEb7edryeJ/xoZLxGUpTdqzuwMqfNocG6uMKio
grqagl7e5xrrNiLFM6mYdMwUFCTKSzXMBIUBc4K9893oGrxAOrPoWVx7ihLF5FaJ/dJ2m/dDOaCW
hGR6NC/Tcv8A9Dv1X/Auif5lThA5xRVMUVqJvFLK6hyFMpeQjJBYiVWwTTgDoszsJpnLAwUjLbM8
GhnK6CjL0fXXDeT4LF/TgwGOfzsusCwy+QjTDBS4V94F0Wt5Kg1sI4aVu+2VsowjXnZoMiNNa2Z6
hQ0b9Q9xl7czJ4B/4w3uejsOR3QurLrGRgZvTUx+ZWmgx2U1+Gmn3XdDWNhDSa87OHIQ98lT8KBU
+wGbaz51FvMqE85Re9kok2h8v8QHxkjCA1oXEeMnjKaZf3A4RakdUrBeyytTrvGifMmH/LIx0GEQ
43xown5VOwIw5HOrug/Y/nACDBp0fMsb+tiNzU6oeThkp/t6eHXNXMRswam2N1hAPfpQNwS7TA24
6zMPlOj0UPunkywoXePmQjmrVzTpPN2CSfPxuaDBfP53wqsrwfmHHMOvrysolnFvhrlb6u/EGk33
Ob0TxZGThjMZ4fhjLeakMwncMpz4k0Sotr5FaboAL1PEOsS8sDT3WPySAsAYhKtsCPbE1jkrJZ+x
87xhEPpi0J+3+a4z7kBANGD4uEpoc9nYpxs9OcWMqTBcNGuDWByt4Utsb62nCuMo+nf1Vdz6u7Dv
zaxFaqt/dJ4X/shy3kxxymN4wKTHJWWDJZWWSD/2kl/2Z0laCX/eG6nOLQI8qNINipXVA54r28CX
FDDVQFAU+xJCzEDz99gi1rP4PdfCKDV3u/lSkl6Tys4A/ekSBPzDd6JUyLmMKfnyhdUdxBrFf/2d
A2I5JmPqO9vHnuGxxjmY7kij2eOpBl7PHnR83r8rQZPq90W0I5TSOxZe5AqG15MR2qCbBKd6XKT7
QYSjFCeYiClJfSjBBERFlhdNIkizYOYG0tXOEP4T9xMmRQQXeBRvJ8IgM5mjJAV3z66uVW8hW1pA
1mwNcaCI7E7DHjl9rpjGSCaIrXuUHemFIg7KvjNrOQeZZcz7YbPvBuds41QsSP/9+jqGkz6JLXUA
0XenypBYPp814whWmLFhoA/nTViV7mjEB7Mlnm9Xcdi0MeR99Icw2huGG6fVMcL9ifr069TzccRF
pvx+bWNu9PnPdNmjS9QdwT3j+CIOr0uVKY4yBkcGj8G9csQFwHL1gnb6mvm/ptrE83qvcnu99g+M
Wl8Pq6hKyoHzSZQABP2+KmhTMW09IFxQ7gJXlu/dT7Mx+2rGh4MH+rwKxnl7n5Qhp7P1v+O8WMgM
ibn7Y5JHySH5Q7Do6kdCIh+fvuT6NRBNgq01gxymnQyYs4tL1b1kj8m2br+g/Wg0u9kwKUzuq8XT
ag9f4JU+HfBI0Ey2w6C0nXzFCXpslraUOsnAxRwxIRwxC4cE9vlDOPP/EwsAv6dZiPLVOdFBTkYm
9KQymxVUkNmot8AEYX2XQXCHQeGjWBo+P8TkksSn0H9K0xeXQ34db4rkF05lxi3hxh1j/vkGS4uf
PR73pNNCz+hZLpeV4VR3gO+UJj8Hf2kDJNp6gQt4latf0fqu4N4JIOeYGC2kictq8mTedk+GoJ6u
DwxVbKh+GcXi7IssnXgO1s0+/Zt03r3E7Eil1QG3a1g+qP27sSXe+WJ4L7XU4lvOX3HsJcMLO5eg
IJ4kQiRuhzDcL+pqdeZVjJRbzrg2AbsXk1SBoCYnLOMkWOjEOR1TwBBVy+vJ9IcJ1p7h/R1ObUIv
t/iSunFnmQ+1AMYJGUFUL+JJf7uGwIYzhtPtxYH9RM9HzNIzM5iIz+TLeOeyjcu5fgB8826DyiTp
4vPX5rT2FjKExh21Q5CcXSTiLj9l6scte4i4QSfPgvxoHXXhZpuB9V/vtG5h+0dpHHb1N8OCOgzg
jzox7WGs0eQAdUu2c3jl5F564wVIVKmKb9k4r3/B2dA37mn8YXsPj5U6X6nR4JMQuszCUJBjM28Q
HUehACE4N/Gdz5vVoNOQmXoZL83YJJbT95lyPYQm01wDZNIlCRcX0l/qK/LYG8nHo1QwhLgJPgY3
SkoZ3P+ZKNUNnyKgUl6Q4j6p4FMBGb1VnKzFPSno0GR7I1jL4T0EsI3DlnyvO9xBwl+ujmMCv1YG
h34jWPEcho4vTcVXibKkiKqxy4IXxTCx8UkdfDTLY4E1hoRS1aPivZ3xR72XP1BBzlg7nWjmWRvy
YNEBgxSNWD7XFDS+Fe4UJllr0Feo62B28MM3fHVyaDvpD7aF3X3OX2KzTiP0cPbk6TqQDrfciZJy
muK9OkQNtgJM2ryzz27Jaa4aFCKOh6LLMceY8vfRHwCOBaqrO93EzTqfCT58MSt1mQo9qVyNmi8L
XL6YUwfjHMgQaWsofgEJYLi8fgeX8SF2DpXG20E9gNpovJCi42s+TuVDspiyy0yP7wWk68VacDwH
Pvsfjm0Y70sNgo/cXOCZ6+FBcUCg3pggs3UY5tKECCsjaR4rC1CbPqWcApfo1JkgEtyWuNtwZN9W
/EnbeIsJriw28iIoRwls8VkJruuUvOQGMusKl++R7ehWFn5DGftHbn8IxzjjBHusByOHQr8alsRp
yGsk2lqZ5nvmCqKnMWT3oW55trPRtfvxjm3m+HnIrB4aUYwVB7eXNvBH8ZNbsOyf1dUGFuEVXboi
UVYWb58iYXe04Sy2OYKMuaK9/4KwnJTBu91lfgcO2RHW0CSCYvWqqintQTaioIIoYa8PkfgcdIDc
tu9+y2NvBJMMP07ANUBkVtHs/Je0EMpn1rB/rE6o4ASRfpaBHUgTgMsMrDhK6wji/xQTqBOTbs+B
oOwGq0a0sueoiYHxiMXvh7atdGyCzk6F7TAHT/kimItUsIzSNmK7xTPRZ0oEINSlcO2aCxksTlWw
oM+otSkWiSovK8BooHgjigK/95InT5aNMMIEO+qc/D5wmD6UTy0gTRKvX0JRwf1AJlVMqETU/19J
e0B12aBe2Z44Tp5mDd70A0blY1QteS2t55fu48Q/JOp+kIntD5zWxvbBIHdZ6Pxg9wRVuPKi05QG
mFpbEb0vcU8Cscxogw23acE2B6YlfMWDCBaCo0n0cBj/NsNkrzpJNQ70yzUnKam0ux/5tTRfCCpL
kZkx7tqCuReeO6IgR6Kta50GLOuBWzhzyD3/Ed0vINNZeT/huH7VJRuVDq6ytoMZUC6YpiCWDwVh
x0xLtiC+P30dm1//oVKSyi+RbHhKV51TB+PHmdo5dqwO3sQXmGhdPOoyNd4SPu6T7UIkf6n0k2+y
kT7VmoS9ZFHAseFG3iijlvS2rvf3Cpsm6Pk+y+HsxpgfTHBb5L8S49qxAKIz/1t3o+Od/u1mivo2
XSNiPwCVbAFbxNEOYaSVv4gprHxHjUESBOFbHBEkOniZXzj5JwsOyh+DNGMxY7tkLj1wMRYDDp19
arJ0g3ZzBJPRffFONSkpUKT1lUVJJQTwtMGrwEZJjszS5Jj96Nernvo1DmZ4V6t9wiSo1yAJ1j4L
qr0M29nQqmvKk3nRVW/HlIc2YSXL9K/YSc62QNJolUJBleMM4fzspYy6FM+bMXjmeIhGP7ToIAHv
SNcSqIZOcTNZpW+cy9qnU2zxnGvJhgSuLPPh8FJP0R4lWPCObe8rzJeMor6ZkgvgKJJf2jpZ+/oF
kflWR6N30a1bMSO/8UOge4CuRoIcuTFwtJQDUUPnk6g2EJEkXPUZwONGxxd3+9qryMZi9UidFazD
my/0HxEYSGV8EBRzG0fu4VxNXsvEnEA3i1I91pDwT/XJRvlpj8q9lWvjoi64W2zZwkMU9Vt2bASv
0ucMrNo6KTgJd4PlZcLWy2WtnAoVKLfZrddggQDsI8qkp6w0y5zukRNrPnNiGEsQLlLFrz7fgbiF
aGh+ez7ruYKnxFz3OaJg6l0g4ahupxmo4owMBG24IIe0ZznZfjWGGfb+q8LpGRJasPoYYGdRuGGl
yAWnpLsXymSNa0PNynFKsJDC000yGgqZ1Eg+f5yVN3AKzDADzcvK8gZxikjJtOazec5RJhyTTBNk
cGNg3zYWEFRUjUjYPxt9r5DT9lzaS1TBpZ8V+Fwitao2HuWZtEHUQz6lFDcld5t3+OCqbFgJTZgG
QBU2BSmdcO6YTIgOTY+EfolyHhSN3pwht3d9FtZpXyZ6pKEf7zvHxmZwA+TXqeLw3qSM4jU8nOLE
n0ZcIBEaQSTPJwPfnREh2J+TrVN0IEwvIL1G+IMH7UmZU0ebjgsB1JQ37lNn/mPhgw7Mcez/u9aE
h7Xw9FmXsIgrvd8VoMCm0r2BhBMM0IBCL6lgd02iYxGwHrAqSkcwRC7H1dJcQWe5tbzpvPfSGTB7
KBuBmsYyD5eMtN3VRE1fnPhYfHm5KWc2c8B5BoQQ9zihBsTGp1BdSkeiE7y7fEKeswDWlLMUhyQd
YaLTdYr5JATuNw0mnXgqHq86lmsy1+104dmFmS1kHmu40u11o+qT3yFzATmeIpJ8BZUHGcUhv+wn
XdONuWET6v3f8hRfp9xWCK9kBO3mzr9rWmaYahuGdjQOFINcaBbDIRIB24Darg4tdZ+wKQ2GxXia
hjjQBigej5FX85bo0gbqEzTr1qpXTSTuAgsDtgund0XC4xUe92vDijeywwxrwE5vdiENjYcwU5v1
k4IaSq7x01lKnIvBfGqpjLJhXmdsLxpoG6phT95W0cZbBKh0yNnpnNN5bwiy4hpmDYVHN7NFqAj8
GNvvegMzBohhXZMb+hU7QPtAJA3EZI5bp31rVvLVDKQzMsYzVMdMVFW96f0zt7o3khh2tN2olOTW
68edrq/q5MMAGhnnnovjAZHpp8cdMLlVOLxVYMFgvPcaLHUf8x8UZCnSsOGT2sdhHzliQo1RPUXM
srC2sR6ZUkWc29BHhM9R7DeQCwBhgk35x7Rlv3DOotK7ff/pPOJmlJiXjRmvSETnmOFLDLoK+ypo
cvIQEK0u1lZkJMq4qgI56bNBldDBJ4yLA5CxXZGXt6X0zHGWaJ2dH+7mTxvFJVKNfX8I2TfIUN4c
Ek2vKG1hqyPA9ihCUQhxsVhBrA3SCW4goACXzDEg8KIWEzFrhUCfe09Ynm083hi6oORU1yDEijh9
Towm0Jis1qyML23pjDWHzdn7zKlx3u9Plss7LeQgmTJ0bGhkJ226wNVGztDJ2OWaKmTGK/ufYeFM
u5ExBOgoTv8WQqSkblkmcqN6rTk97Aw+t4j1Hcs6kbkrqXIvZoI8HyjDG4LAxzDaM3j0y23ovJh2
HvrsquO4fx0LFmJ9VR4Fvl6Z+mfcs4qKOqcjSYOY1y2p287Wrxptt6L6P3PlLXDzX2sURUBP1sDc
zeyq7l+Qc8IW1+vNWx/ni649w+0SFW5ZGM3ksTgBtCcjd3G9AoQks9Hf5WlGgjcXZD4GSC0a1kZc
Ed7msxH9KesyEJhwisuOyBOkn+VIqIj0QnY/v4qH1hdZPbpfOABTXvtXTCPp5dTEDx8bOwxTP1wH
sYTaTIZ4/Kv2glAU53x9AxNT2IMAkYB7J/+M8C03ONELv2Kzq3dzzg4Fz3RG1qKySLzEMocH85hE
Dp0Uy8n8ZTIxLP49F2PixN5GNEJ5Zl0mkFo7gDz2egoCCqDUn+7BjLC/gvWmqnFwO42Zuz1YNzRa
O1gjTIoTjvl8z940+4/wq/YIDE/pJGDhx1KYCABnynoq6bwGxKY9Fwl7JNQVLsYE5i0W+gcO33SK
X7WhP0enO4bPANZtX4urriOhC++c2jyhIYnQreOI6x7tICnUqhEOzddUZJEyVC+NPWw65slmrUsu
9EBw4ZaNZUb61eJlbSHmdRMtzWlTwtpo07kRgKkazmP4wyHgftqOGxKR6JjLtRvAudsh70Vhn3H0
YExcZo8nUNDsBQYtEm0V1PAq3SWkf52ufDgtl7AqAGM97Xa6n0RcFVyIlVF7q8B+g2jkuIltO3KR
eyyYmS7FLJzdZR1Eb8Le/3AeAEVSJTYDy36Kxy4bJe/7P6zo/j2EfchUd0DlkFfmDCvgIdy9+a4L
ISR3A14eJVlHyXEQMcTPbAp14n3dxzxGRehIG/5RQySKqZe10IepMe1wc1SuQ3TPWJGt5nk7YxPg
IPJMIAu12ejKIc7D/JCHlPVXXZ7SlssC6F2Rnuytd8RiaT5eNHf3bbpLxfzCLLDPYFPlDBJh4E4j
lx2o/vF9Y8YUMyGSiHnEz2CXg2faDjAIZCTnRX179tYagKQcZQbMNtDYRC1a9EbsKY6J2Dn0Y5D5
Y68rngE7NwA9y6JMDT15VQIRIRDLHqi9Zrz3KacyoCM7jIn+ujei8jKe/dEhaK3WSbg3ll96peZ4
/KKZilrgZ0IZw41yko2fp2nMBdCrIdrnxl5MRdbXUIzhLxbQvJryhqhWRLkrh412Nfx+KJZPgUgV
k8SNhDdDu3ZTTsBL0CKOUbwZIBRi0NQBzhWUvXpaOubZQPUQQGpjHYkLE29d7xFY65pdIptdJh9q
+I2sno5Kiyy4ElTTJ86J0LCwRvKALmpkqwc2W36gFM0Ut68UFKvq3mtLyEEApD3tJMeWFWdozFAI
SauL0mFjvPz+yJqdQoHpMifweS6Y33OLk5NGbiKYrdmBROwTHJ3skkpGdFnfaySN+5ADEahyaLOf
wpkvJrv0Ixee8g4HXrln80sKYJczKsBSMUFEwmbiXEUaV7FdGgkmcxFoHUAh4M9xSHChcTvVM0J7
hmV03jZJwHomp77BdIagi02fPl2j7fBdmKN3hvNMOz6BXl4J6gNZP/gDRg18p+Ny5zJGMTXOqHxz
P34oZB+gcIb6Zo8LAa5n58RK06xZQZwrm/f0Fe5WhqQaTnan9rTUtKCUyAVawvSuF3VDSCtUrPZn
hMhqgcp/5U6aJLX9N4C8C8A81vSVa1K4eS9amSziWUcDwB4/rZyoZB29D6hxwdWuNE1WtKSSLt9S
phCuUb9VI+j+b11XJSKCteLcHBE+rSFrGeK4epB4GUihYndFlDtm1ocmWJNeBG3G82WqAeXqzcD9
qpgwhMGPz68o5BJiic2+epCIFmfM/WOBZUKowAPjOAwG3fQDJD0fw9SVy7qgAGJxPeZElqpBduK1
oVeKHCmlhDj8HZLXGXo8S3qyNpc/65JCQEmdr0Wu0DCBCcriKtmuE5uXrNc6j4BajFVcP4jJ6ATB
9HVpf4HffVitPyXV1b+y1BCZEOeVmVjeDwSxViGO/PqhARO5A6IrnEIlSUXsPsKAl1LBi7kGQxX6
oSATzlAUh4gBTfUQT3NVFSRM+SBgTDJEOTV7gwbNGSjZag0S1Ut5I+sUh0edvFxVQjJ6j3vshoEK
PgWnODz3wJIRjG6B0abAENh139uvx/3WmYxSaPQFsmdg+gySN1UqTW04DbifToj/WfYmV6ZU0yzG
LWBFfILR3Kxw2vY5zbHd8M2TKxDGDYD6vurkgfN41z+Ys2gZhiEXN2BngiAaZM1DPGrl0q2/S2UO
9NwXXloPjbRZYV216L8JR4DWApicKR4GgXjimrDN8CCoVj41yKIQlKA8l0N3q8ryACSFHvBn7p2C
DXjeq2yUBG3bl2TqUHuy8c+k5M1kbf/iGqDaidp4r3i61a7olu08ufeO+CvRdX8B3bLoO3wqpJrg
UOB/kTnnX9Hb67SvUfCbNHcygUKoUTxrn9cznILfD/ePDojcirvWBeCw5dlHdd8DSGMOiy8RBota
CODp8o5lylIVPRuvEWCfL+PksHre4K6QoquS0fcs0dHUpSgmG5RPJAFwkQjP5X5T3fagGJQLSZU0
sMMcJO0kFEPf81rzFtcoGKOmdNbV1Ccq/lYejM5xDai3pCuVnLcbbtj2/cBJF/WXP38MSCeg+19Z
p3PTr4o9ktZmV4T3kmu1C0wdwMfTo2BwQGIukmEFf8oC91CGIGC38yy55l15ZAIDfF7xCZ1bLvzv
vy7eKa2FA3aYoTDHd7glJIxh4OLTbRPWjAthFoqEGgEx4FnJNr0Q3a8XHTo2vgsjDmNLyOjevXsS
ACvo4ure/5DeQNCiANMu16b6sRNO94lcQcxdZaYZPcE7zPeLJbVJpln4NqWhz6VCztk/KfaDrFzG
pEitC0EhwFXzOf8RnssU8KeznA4JBK9Y+y3o+Ft1I8lUzLPdQUO7RxUR5AYmbqnsCQmqe2MXOmAs
oFflouPWcN7jhydoXlROCRTfRVHZ0aio7ljbyICDChswsUeQAFRnXaVnY1lvYFPimgMnW5s3Mnpy
YCN+yp4pHrVjpJKuRyQLtx0PesiYgfiR6677r3JO0WGuOBzcIgVH6Hte84VXwaXRZI4Mc8+78yf7
TN6YbTuh7TwaINJRiLGVwgPQxgAyclNbArNeRSGqrT7SGSU5dEzR8FmCv6EAyWoDc7smhsk9ttDJ
RWbG1iLixyxx1Y2v6guupTfH2wzdD1ylhijTU3A0aktHhI+RgErcmIx4dIgvmfmNZdT5313dSZYp
szIUY35SujOmhuj4Famd+At3wWZ2nB8A+aYmT8Ai4TBXaH0ywoAeQMdl0lcTtlKZTIK6EqVyPKqY
v6bGPOWq1dO/1r/RRqV6BOBkYPklGqtWYxxMHO/nHj9H8kqO0eKTW+lwrKOfNvU0op2uRrqdoZLP
l21+VUBY+ouohpZ8IdGWsMYe0bf8+D5PnAdBc0kLNYNXavymvdHJwUqdj+DHCxaUabq7FlwiusUt
Km0N1Npe6qv4AKHYjx27a3ktBkmZsnpYyry+EYJ6HMTKbb2RmM2Pf+tp9PJW5dFNTiALP/6uTsJt
gV3vv6sUVyKa0i6jrgUoSet3kPiEi1v0nNkd3/cJEr89cS6/hcVt6Z6l4C5SByPPLXQ6Khgt901i
xb0wt7X8bxpw6233Od8oZRBzGzDymASaGVCWb7vs+w6bEsbwBmqTK1v/yBjTjjqS8lptFuB/ZN6S
NjHhZJeznFKfc2QU0Qj8E3CHegEPBJM3H762pnsGigyv+cdKYykxTIu+046H0mYs113+vZg0t2JH
ijfucS6qYFZdIaEUi6GVvCElGB0pBR3oaB7oLFZ+pEFninMtn3YXsMiOyrAc808l/fdrO4W25ssj
NHZT/e0pTnWkQ+gnafqWLXHPPtv6HBMDhWS62Wyn4+v7/Dn5foZ1jyHfjZalt7l0SIGF8lCqTudV
91y0vtTNOe3tG8iTiTOFaD6FyQP9kuaVvnqvAgigNDqicdYZyxORfV+G0jp+FgAMBM3h7g3+TXuv
l+s3fuWLmrriA39pLIx7JiTPm1aVwVANcl0dp+e3ZsTBxTppnro8Pdr4z7e84jsaXVk89Vjcau4y
olY4d5nHkaoDG7udfdPQ5JwQQNbUD449dOgH91n9iDs2DsuLnlmiM4V2bFp6N8JTiYS7oD6/vpn4
PPswL5NTVTcr582+C9j0jjZ9Uk6SxbyOEov5LCIbTvlh00G6mrmPG04uOLwGy6VzrE/TBWicohA9
siAW3Vix3rN58u3HKyeLxIzAuuUHFmhJYTBqrBltCxx4D2c4MADBIvntYnznmOrprhHkc6NlJAOl
T8Kf+F2ijsDykKbod267jZgnDPW8DSM4M5voGXgjz4nN55MVbZa4GQa6R/ASTJa1ulZgLNGPwRm1
pyiRA0Y0pzDhjhvkCiThe0qscktU7fYa+kcWyHJ7qCOMPbvYKz1VQEJFdPcTs7RbhhSReSWa65zQ
bdjwJDqykPnyyQOi0uC07yXLXcd0eTgwmKpeRv9q/8TzGTVAkMXlmvcAX6tQUUzir447EUmoMUHQ
R3pC/Iygoy5E2ReSy0Vcno4ztBihoMtUgidvx2XqMcmZRYkTBJ4WBz62u808W8gQiSc1cPFZrCge
6VxeaPCTL2VfvmpjyjoAbREyKWyjkRKFGu6o4Vd8ecoDmTcvStQerlEPdYR2xUkTU/bCW/u/CAXe
qb9Vp/DzhA5SiFsUeC5ORppursum2jA92D6OtCvymFTkWklNlB0DRp6IaqeP4lOPkEv2WTx9545Q
OtYDJCd5FZ2GT64y7tv4lgBJ2+if0dQKrJDr8j6nYDonzS49Kk+9iK7yHZUrXZkPY4/sg1k8EVdy
1QJlw9g1D9bDSNtd0D2ylKAUTUUXO9whMsj7LnBymFo32tTOQ9b5+nF6DV4f1oad/xpyBQLMknJs
XgH12ltXCMe3Zp91EsWHv+eb3B9cUtHTxx9b1CjAcor2Z6BGuqq4SRaHfdZN2LxoLWR3cquuFbVG
j3282IdkWwCdD+9SjWFSbhaIWl9z8bwmyNlIOmhTxluOuJd1r4NyVEDloaDTOX6MQpdOTKl5YcLt
8NVeirwzXfAyTTir7osvm4pl7Jb5E+IVwah6nOQuy9ELtrIMAN8bQTkntACGOlJL0dLml/Z0aKj1
A5+qZjG9wBgiJbMiKVkXNmxjBFyDhT8uOdia/RGQsTJzgPTaBEapX/ngeb8BmXKxSjCREzdfuWSm
zzt6+ki2VwkrYHwuclz8LQZ0MP4VfyDCxeD2iwE2BYhaOVsrdghulKM2/sCuCWRAOl4x6p8Pef7l
I7t2mDPqtnQqmVyk6KGdyuQrH8I10iNgBAip8Hy8pH8wcYozy6b7BasQT9WiEUxt9exYrnN+nXZ6
vWzdKiGCeglMYpgyrUQZDpLgMqVrlOKhdniq0xvkOkvusXFMBob+3i0+2Ftqlxm++hI4LIgr7QVf
5kXusCJ3duNIKOYHHcQnhsJlgdPpPrUjTtlATmCYbUQt/BDh/bVc061Z1cK/xinUzU4Nlwqwd6qu
RpUsqeQi5LKd3JIpUHINqFtoCtGZ+zWdjYmpirTRuClLf+uySol7qMMXTdxk4PSTJRMLlbCHevXP
DM0fleSID/kH/X8C2icwthLl+T7zVFgleH6w0AdwrOQ/ketl+OZERXGiHXaABWhN8m5nCNpYqLjb
g3g4G+DKXx2poOiW/cantXnAz2EiXzXJwX5Y/c9oYOT4y679OPThLwKpz2TuX/Jt+hEgPicGifbr
Ieplf4PiXM8rCRS2c+FQchOE4m0SlQ3718qPFGHpaKuuDrt5BRRkYhwwNtt17PZnbhXK2vddqDGq
6HIYwvHITxUoFdlF2mrBb01AZNEiwPJOQScgwnD3FxWpeNtJQKUfqSbGI/Wdn8/IhZMG63+ieE3Z
HsBj6Hia8K1avi70UvBoOdm6eyx72cNubc1shfOfmmr1eSeNIe6WxxAgBdCidudbiSlP8PgquVpb
uR9C4o4POJ2aFHXSTqxwoo8CF4m+d8NOUNNTLVWU2IM0VGuQVc24Dd6fPclgWRnC3OQ3QFtoqvtU
Govgh7L12kixVrLbft4CS4tHd2kIc/fu+vPyiateitCxRYf2UIHB7n13SuCROVgDcfnS3Dj0WUuX
qVocdoKaD9MpR/ftrPdyKQXGWuIMQCpCC3UtSKj49+IX91e6jXSb35N9j9D3rIm9LwP6TcF3rFVO
RvlOgFZpVOYA4JaPnKj6ag9NqQt/Zqsm/jSrEI/kUM8ckWQjdbs7C1aXfEOA5xNhi2KrZBcs/lxq
AbSddpcqrf4hd+nVRsqQ+O0kWCTO6dKlgvblseus+MqpRST4EzvL6YMyVwJ09w/+homVU+R5yX1N
mzBrQ1GzVA8CsY9lmgjFGNP8H4xaAwlsNY/IHp0lwSlm6zDOTITon+KSONWXDL0NX4E/mt364vdy
veJ52nlS3bMXLFMa5v5+vn+nFSNwDE1Ctugs3S+v0cWDZ//lHFwrELa8Svu0uQAaTJhY38Zd0u8i
oMx4+TTZI4VLjIIO1SdNtKJDMuO0ZpvCqMpQmCM0NF+8UaMEg8F0LQEnKWXkLkZd6MOo4gW8cVln
0WhJSzD7YBSUXhrCaMEF1VjlwmT1cCtne+LrDor+fuYcFZlSAhAASoIDLSGsHOi0zrBtiSW9UrFb
EphqzY3HbVHN8y8LKos6IgNOjMV22U4yMgHLlcIu2NmxZSfI/cFFjekYB+wbvBM3s6eZuVsP7gK2
/7qTVk/Aboa5FmGP8ZSzkJ4T1378+w2oi1UVohGvLl9c8O5UOO3bhSjxPsE7oiIR1dT3K+vG3fvk
P2QePD0VjfKrpJLFotxJmQM6segT+o5i92fTbmQJ5avIPITgIVFpGskMjaM97iWQcTULoHnggV3m
Jpf2hkcko7Wzje9N8ZEiuvgZL9UVCm6OrnGzKVQuS8Fd14SqTLdElAngjgfoXbBZo0GrNv3mcd+v
N8sHAgxp/uSboNtA+gURuWvdwbpE9Idm3aGoyYTtP/ozcYMh9R1u7/arlBe9ewDoxjbZfw380ysx
JJW50gfpRK186GPeWixitDQJOssfxTn8Um4kPnVjJAaShnQORDE573B4T9FOQgC2MQ6lYgGH5xDf
/ArUdizueajHoXYbCblOrLp5IK2TOtanHKuPz1juMSoPak+OcmcbV1eRqwFYFxH2qbJQ2ufOTkQB
1ya6bKBuAbepM6LtoL9dAIpyyWQoQP2Fx+GZTU+xrAnptoBC+O5Wrb0Y8lg7yh0/yiU6nR7yO3La
tDrHF/LrA6WmW6ew8Fup7hvdjoeTNE7d8ykefljvfqFaGkYOsUH/QL4h7fgZIrKBhKAIFH4TF1m+
wVGN+p7Qxg6Ohxr8C+uzp4Gd7FYRWG9lPpSZnzWE5UOnwLjhWACDZTbyaRMa+fEfpW2MkI6PhCDI
8Bu3fF7UC52jttScq45prBBmQ9GSRp6566dbsvDAgctuSCQqAS7ga+6jvjZKFoEV7QLJuzF5ZYaH
VPgY3XNaWFG7rayWypZgofcxzOQIQyusIVbEq63GZ2+m6DgR+xgaJSTmyRzhrLmc5XK6tRaoWhas
B6wYWIV2SA2/8JS7Zz1vOQ2d411fXFyV7T61dr2WSxdHvKYTvb1P0PR+//boh9iu69UlIvoQhlHM
fSPDHl3BtV1JNx/S4CiTsETu2BQMXxVBpw5qdKjul/o/LVht/su4PGvFbEc1srmQ3xiHklEj4h+k
vKdr2i7e2DCy8GdBqKTANW6X8/oRK8rZW2uKilLTh9q+sxd1Ki+ylj2YwFvMXHBsd/cF35jNHkTt
9zwKKf5bDj3lCibwjM+vruo5MCOX6LzuVfgmnjE3AACwcM2Jbcdij6j9jhhYPswa2u3Nkwy4eklA
29eWGkzgs1ASQ2z2yrW+P6Q+lKaEOlstyZrBtVcg+CoMAKJ2EphGCClRjyZpOYeWti4lwObuQ+vG
tDXSpXYHJc3Lre1QEAlUqZy0R4ruK5EJSWvKZVVD2cEEQWRYPUNYQsPDiCwPhFnunamWnoxi/XzB
B5ljFMXjVWCmCp3lhdw1OfW/5cNvfVHWo/Xm5MDlMJULNWqQe/Z2G/ibLT0PdzOMjerXj3isHJ7/
TrPCo5nvMjgiJoCxWOdo26zj4/oVsFIVDOF4QU9Ng67kw5P1eJX20oGohiPKQObwJsx33msmyfr2
BwOOxCvS/ltBAUNm1cAYH1uvkZN0q71vRWstq2cVQPedNSFsESiHspvF+D/sQj0zuMllu8gg0G15
G3ZhT7wGoaMkZ0JDFw7ZM3JprdkqPlmB19pGnNs3ruSlT8+JUdIml4/bhyEzhGK8g/JRDikPNXJ2
DcZ55DMwOojTSzPet0GQ3brflqN+dJiUvoKvt8nAml0YuqlKe4l3qc5orUOSYPNh55mzyqsHZyZ6
xviWbkH8HlTIUbTpSYMjrFbQW6xKMNuNu53o4isG4sk6YA90PGTPqBgYKWyT3/GLowPVWvcXi9+s
1+lfzw0I+LUnc+m2bFySxJ7W+jGgFChXdGfl93DPCsp2FWLq/OUWz8lcjOxDySAlfa51C5DxmjKW
rFD3N9jSpIsdCUJyZWsorb3hNA7oY8Tl5jtkoCrvOy4QRks8Jijnftk5ydYklt1G7UbPCQ1U0h7Z
MECKVHDQ+hfIKZxqImN3UvfgSe6JbticD3IgvCLF683I/K017WUkScuWHe3lZ6s9P8iQ2IoSZfZ+
gQbOQSYNHMbBNZCNfLMobV5RRBbeqvU9f3v52LddpVY8NGZsmxKVTW/9G1g5v/bf6WAXLLd1xmBO
RRhflMTlW7Fx/pQj6EDXj4N/D0OYpeYtzdw1/lr9z/qe+ehp/+OjEh2wt+IlzzFkFPBBnOXCHmOx
b1x0v/x+Tx51XJ0jhdibxDKebWUZIwDk+OK+CnlRL/s3hOvpXCR+jzIS4AVTSpu/z1v/zq84BCv4
JRXrWa8V9RsBFPZ43kTc5jXPgOjzLKZVxMAA/YusNylW5udvJDsn01P/lRLTujo0qLHd19AX+VEF
wmk3yXRa1PUCy9IAdYxRP4flO2MDaxVyiJNWJ+Y0tdeUpxmPXBt2GN77vNkrsKoWr8uO1ueB8tCx
+Dnwk2k84gUfhfu+NMQlxla1U41+ogu/QTZKq5q1vCaT0RsJzXB8LuZ3zHL/9zoJSY2T+ypzhGDH
7VFbSmy1qvZvAmUI4Q2zrxxGwT3+TLDA4nh1WFV1I75BYc9rZ+mEGDIlpWxggi4/kvKca6ArRoQF
NYiUdGH3wCVFFyudbCxw1Ho072Khgo610cZB/kem8Fv1rD4gTHAO8dObRRf43pF7j33w3NphpCJ4
z9a25TAN6ckygNniOKEDjpK2CUmvk+UUq0XNEyqbw1sthJLPoX5THu4xB3E/vcwqwV71VouZWnxn
Qg+4AoDrRaHYyv7xEj6hlB1R+EU1G7AOso8A91eD14d3nIcsDGgvkKmokx1UWd9/xIP3tLnMERc6
hb0N2NdiriHH1wGMOpGmeb4sNxuYIzXfsv+8rgWFsAfPEoAOvn+FnmOF73AeFskjb/QbAK03dI06
G2dlooY4TCZuua7suYFa/jVEAPAVD0v97T1OhgsogfjfXSM8k58fjh3uWDYXaDiNTEcM/NX5EQiF
rT1vc+hVa4umltuwSyjQwcyYW2Uw4gDDr55WI2HqU0FPv8Bm4Q0vSPjPZ/wU1W0wwC8YjXVBzvtj
Vs6EIQlTpolRv5byHA/PbHGUZaY/XFTFsrxzoU/lHHBw0LMGr8jxb25BXXM/qc6bNSctm8e+aF1g
/++3DeMwQx+9IIlyQaDPfmPOkZF8eezg9aFF+j7XEstkPyqjKL9MYyGJIZuL0NwHYTrwPAycEzFl
V7QK9CJUCnABjvqI7IdBNa6ukYdwpU2d9HR7hMfkZzBgK/rQa8JYueuuHe3NpLfhZzwktEARMLxo
r2+m8uSiUoSgdxWalh9GZfwb7SqeyYtbX6MIyziJ8c3Mr7Qm+eM6voXpM+MdDZu9EAyvan8ssFEG
adpZT7ul9IeI5SBj1uihRuaRgvdSbJ+NAZ93sAGpdcdiOf4EkQ/i3VC8Mk6t6bjVFbidTY4JsSI5
QFOgcrI7v9/NreSXej1mrINpOju9UWVY9NDTjzF+XAsvSpNkuXfLHBIz1avV3ynUvHgblS23wb7s
x+U2IQjNHBGSQZ5kJo9IY8CXN/gnHDIzcTU8OzpeP/qdvceS0Gie6aUK9P9iTkgtIMc2u2OO0/hZ
gVcGNTcc2ht+WyE101rvDmaAQ0/xnu6OGM9qsmMmR7CRsQPLZ7vjGbjWfbmFit55OCsy+SRudIS5
xSCflBEVtXjPxXIThm+NGKOv0WDVyvZd2oQUqUCJzs4f5MGZ3Zm98h0ROlgcQbolP6MYWzmk5Oq1
4pQtv+5hqAIysuJX4kP/HZpylcta0Obxp8FIjFM6bV/xHsXhUmoRUE5/KHO53uHMdofpX1MN+Q5G
Pr2iV9MAprokVt8QntdUyJybPGRmwNa4p4ZwRrlRtgDOhrm/aXIsZQYV2mGnheeb9KRLx3pWGX8c
X3BdQR51y0xMz3QSySlEvQ+OROGjSYdwTCOluHqDHUG4OSxsoyt/yBm48QQY8aUkIVDI2JbgNYMf
HluNnjw+aFzdfEqvtHmoN8/9un/60PwJi00jSdjGO49vgQNhmCDbcwGAUOhW+zUJiDvJchHtIemY
9ypde/d43lcIt0e/qxWuBJNxPsXJm07z1SxFBNTG856/nlT4Hh+dqcPH69fnKa5NOSq+gKk14RmZ
SVETYX05czSDll6pT7LorvYkgEFkCkq1rA7BqxpOvVt49FQM5BNYkkT6OZ1l8ThS+uXu7sSdOfaz
av922JtkIV03+LnqWCiOWXNkeGEbKIDqUmCl+omaxmhJTcLDvvc1n8tnOL4CqePiKxh+lpU69yTu
DtCB7l0q3mtsINv3NXYN2748hSYH4mPVO0vwGJ8Jv8zlLyNCNMWkcAoSvAoFZ7G4qnGFd/LJM/Ip
/8JAfRfX7ogCmXfFR2X53Z75MV6bA6717II/xdoXhsg2YMJOnDUBZ0nikH6XlKlg2+gWw4x73/VX
JcQOP9v40QQrI2IZggSvcsU8WeRxAvijh8yZj55qsekEv+mWdv5FrvRrqe3KRt4wWzRgZioDq72f
ZBfihpGtKQeOa05PlIEej0A88sQdv2YwS7FdynWlu5WXXoSqqulC9wYxDC41ecXvwl/g/10d1c6M
Y6CepWpeKxyZZavSC/uSxw/OiU1tzT0PAMtIryFmbASRr50zemQp+gYyVDXN2TBQb3Wt7xx8nzdl
xa7ISGs5lSPrkHgrDihMyQEvhAJLqnbmYY0ji/EGOIswj9OdPH3yWUvviyLimiK2CDbVZ2O+y1Hp
h03X3sg4k1KUovXpvtBqFHiU2X+XFhDzFLp1x0yO9UMjXQCQGsp2l5MweZUi8mm7YT8FUobMN5BZ
Ld0z4cr3MpmQ8+UmEIOUIqC0eSdBeTvlKUV1oi7DGzvsYO9XZsYAG84DLl036M72dkcp+UGY5Uzl
cWxgbFstzI32433LYQeysTRZHbLoPbBlTA5hnkhzSU9eJT+pWFo+graFCEF852q3HoSlqT0MRJvE
ZUirzvCq2vGEaZl9TKmsfbeurNAN267HKcveu50NJnG+j8LuDyC7xoGLulUFgc7xzQOt1XGY+uv+
c2rlbL3omyCjd93l3kF4z0vdX1btMMBaPywSNPvFJ3a1NGcPTuhVZEpmN6yYvwXVvwZKIyv9DSfE
tmbCE779WTIM6aibAwuBTi6dx5g8aHKW7CMRaODi1SPdkwtDUx6FCRU9BPdXwo7XlV3N3+8/Tuz0
z+z2RuFdt4nRjHmXaU6bGnVbpdlv2bYgS6bnbF+RN15h5N1pBN2GYk4FPVVnusSzhcVf9Krg9+g6
djCr1VwtiWkMLODuJf6gP+ZzwkCw9xD76GcCM5NPxKcTitKNgzUj5gkFe//r3P7WNWyo6LxTKxO1
Wik/E1GT0GZbDBoQvSpl0fhvUjyQY6h0sp179vtGYqYK0Ud6k0yO54guyoL+Z5anwpwVbHAtKD/R
X15rP74ZLdda4IUQXSL1ErWltyt7ogqTO30owCKJNhW4eGPQy7n1HMPu5DsAhIv9DL808OtNLnqO
xXWVWK5dSOk0JoZOkgoTOp7pUgfaH8uiU7Yr0ceSqUZnddOgewpzO+7/Ay18RwQvuU+/G0nRC4su
jLDYG0mm3blZYNxzasjz5DxJG+irDenOU/0V4QuTbcsHVL+rBJDqmBhy2XNdlpGFW9oaSa98TLK9
mpxkKHOnz27FNvIyc4HhW1XNlMwXmB4oYa+cuDcIBsxv7KgbSMMeACxebxhGUbW+aJmdQ1tG2PbS
N8lNAYYvuW+nDl7oWS4XEph9GoyVX9zbm3bbMJwBDy/Hq8W0xLM5cC5m6+8fafFVJ0tAF7p87H99
crzhvSvesRrVKum20BRtO/dw7iwfmD1cbg5SGTg3Uad1GfKoYMWZZvmqhk8T1lCz+FyWHw0YjvP7
oYCbxppFBExlWxyCrozqBxXRM+2mZXhBpC6vKTFYMGJAki9pH0G1wdVapsWAPAEefEnfN7/0XIPy
L8YKXFo9Se4eX3s6lJcr/On3GZjR2AE5a3orEGibjBLbb1uc5c4+TjmJkh82NWxgTfh0nEttT9oZ
WafPgXdGiwf7qiqgEfnJZ55yBU5eKCvbt5OZQX4/WTxQbR/88CanyOAPZDyXiFXQ9QBqPaQKRIW9
aQu9SZapMfy4p1G/hfFlfse4LfHwNPSfB1Xre0/a5C8waPD1ltZJQuSetr9xuINqfRhIy2pCPmL8
2+yihQHo/hfxqFafTMKRQHCJjfggkDY47AeMMLDmXPgOfaCMMPw5GiZid8aQDqxIHaxL51fURffn
20lXU64TUN0+qgdpkpuyVd5ns/hLr3E51BTR3nwDBCwHHpNyQ08PjoP/StyeXzjyPIJJwgiWRftC
QMXBmNCTPExPr8TxsCPPH0dWdLny4fKky/LGjlFa3+BWVKtWJ52TkTk8UBitxhd/91rTo+uGlnMg
VOcAbyG92alMWkWrz3GXdYBRUnJayo0l0+MUt428F1n0GWWkrxxvf7Q6jF+tgHovnUK0tNxnzTMH
wOo04LoCPcfiUiei/ArxNxfW8GxvytnnEfrpIFWts+BSDJKjPyyLXyDGWWE1C3IjKqD8UXewDNDm
+VumrB9VSUHTbQgoZZLgWPet6yz0gSYCkz20XHYS55Pecw0R7ZjSFWMSjQ9evZSzqLRpMHLdMgnl
E4g+fKGWKNkc6MVDtw+2x7IzzHV6rHtFAsh+21PrygF/l47IVh46nQeQGjdCtD+E4Mvu2IbFw02j
Ckwk6+fcu1YoX5Vsx2LbJdlxqrSCyG63ZimoUQvIfAurN8Mvr99jxYFT9a3xHNopRVP47beKSG93
FIwo2wbcrGg3vJu7mIBQ1SwsBJs8uaOP5Yhk9SIoWAOnDmqmILKhx7NfsiuhRlcbDlp9ZxNZNIGu
Hwr8gySCiawJ+QmbIGHwrpwmlX7lvrcVs42Yggm/CPYdYvQrlaEB/WpBGNewXf5WOOL9JHKCW9ZF
FXQUQ6zfOi1sEvf6aPEkMmwpXPzKRYdxI4S8TrS2f14XGZVnzAp7EUosLsZLsotsWbJmjF2G3f5Q
RlQoA63d7VWt05V0p0gLEloeYDoBFC3GOvLPSp0+zgG4PfhPP3gIejTwVdin+HmjGa0gpw+XW2pL
7i5eDTQdFW7xWwLhLTu5HvyE74ajfLGhY1IG/N/i4Zbh7uisY79sRnPV2U/MOXUSq8XGATGCOqYE
ZsiYEppNqnSeIgqalXTBN9I+UVk5N2N5HhJIlGxX6EYwagxOlriohnYy2MiXbWqG2wwyhod/0hfR
IedcioIJo5UUEJKb+5MmCT6BD95Y5nWNF4BpJNW5zjX8+UwjK30jHejX2aFKHvKJAxE2dp6o81RX
5pnLbdpA0ra0gAv+8OljKuwF7NhedI+NunFMUzeVtnxUoPgJFtZ9WEZgJ+1YWZg8KZV6fSwmFcbQ
Tc0r/d9mh3mODVim2qbc7x1nJzuRWmTVFSfHtnqaMTJ/Lc7frQlt2NLL/H0PShB7Lt65vmCicSaj
3+K4G7rAQ36OUvKNYAK6vylibmNV82I/bnkTQANEZumn06i+3dysDhOXAu/LMoSpTCTgkXskgjGg
AMcchZufI/ItYBJ1dEwXRNjkmy7rrboPT4wcOHUipbFtoLZW8MHtm1wKv1+G1WMvCwgOg8djqH2n
U9RfKgxai1AgHSTMuAPBZCVN5W4ADmrYzUZhq9cPiR9teqUqwJxiwDvrPBDy6hPceHzcfMEp5PUB
CdqF3fhwV7etL/mlUZEARCWXDkL8xYwYS6wVkeV4S75pdQPzFv054FL76nQ8waxDyif3S4OWdNUe
6AYPH26X10m0TZF1VuiYz6L9c84xGqJKrGAFTwAqQ4kYb6i60Jd1kOlS5klqNPJ2kHBf15xeJsNV
yomYqEDJTlvI7b1cbZnx7+qUyu/HNF+SaI3K88/r0DJmoh2ahcOqcrqXFftDnTSdEbQHZzyXA79u
Oac12U4zplBeRCmfHeECE90IBkhR0vKfIQKEcZ7G1WcwAzg8ZKmL57O7+E9IhwvmfYFP3Js5uCpO
yQWvWiUTxF0+2abaWn0ZEGY43S8Pe6UdGsbZdvm15D/S9Z0jEum4qwD/LVoX2rFW/dQhScvHKxY5
O/GGSr+36zEEUs04aCdez1uY9BTxMPbBoImf9PFx2NTO+l4n6SMx0rw+RKaKFlG2w0lWDWfZZfRu
Avu/FGGl/ck0Gq0wTkNvRW7QSIRUYTZcTpL76AJ/noi0s2Ty8OU4jguCeGRmtvDzWXIuiqKvw14/
a+zj2wtmNiSkCivw3DmpQ0D37VQnwFpa0MECIBnvfSCa90csGmwYUUubjvYkWbsjH4In97gwO487
E9qVEasel2rGGKFjNOCFGe/Y4b1hBFOASL3/osda0OLQMoARdQHjfDWvZGyPAkBE5SLRmiVCdIpH
R8YPwg+EMqUA6v+IbU0u4DI3zQ2UhQBZvVcjw1vjphsDFBV75tCvus4LRWtBJi+DSXa+1Fw6Zdf0
cPIOKZC54LxnqlLI0o4Np9r3xEqsWbok3+3oosH5bhwb2a1dsUZUPvCoWthzr+eqoczD+Xqjm80U
Gof8D9TvVXG1I/R8xVTBQJD6HehNhKMeAEqWmDfVByXhXr7u6ciRHoUt6vYCCJxtHXSMCLPa8AeQ
C7uS7EfgkepnR+JeSzOcpXRw5ygFdFaKr8KxExuJf0h3OSx0l6VMB+AvU4M9kH7bM7ZPDvML0FBi
qO8tPe1G41M1bnuPvHEYavz+HMmRCtsB+Er2wFWQSN+lR5AROfVdYBSju9+d0V9Bp+vepLIxe9gh
quZmpzzmhqenst99QurNvV5IMSJYQjmlMd3SrXKCd89V+BxgEv2vD63NdsEd05VeIBclx+PMUQKU
VzsgI/CkpVrgDgx8r8MxrzihTjPQUZgrnf6CfbQ1LiCnrZtNpid9WaWs/rEP0vkuluFjhZjvC42m
Jy2tdVVsiNLBHctxtk4vMidFzgOPkmMipLQ6GvRLZFmpmh6uxZPz1KZCr9Y5FCIoMRNP9XFp7vxg
ATg92C/l6EJcP54HtKmjH0Kr2clHyNOnE1Ofkw6CFieLof8dTskN2ppZzmB3Y4YmJI7Zy6ZibK65
9wpw7/4WBMwDiKmz4fDx8tPXrYOE/6MFBXKnIB8z5vZhMR3cI4COuqhTMPcYzjVcd+YLQyhSB0V5
nIaMY5ZTx42r8UrB3K8/s5O2ZsmKpvW/Y5dCokgIfi5jWOurH0suoyxklZp3U5PaGI5UYLcYJjms
WnNpxPOFP7kD7KpVKz6yaN4cW1oIpVZFHvoTD8caI48M9kF+7p0MbFn3CrRRp3KnGzu3gLCoXtsE
8nBo0ZnHSDvryLZFw05XkLhIYDqgFgYS6jqPNeoq+fOOPv2AC6RY3+sipo01mifMdrUj/aLwr9cS
8ZoMOTAzyRyvbicQtIku92FPTgFiqoHOudUSO1b1pcvfPU6uQDsX8ix3nxVt94JFB0UO97jpE8c8
Miv+NY5sh+JRuPo1J/a6hQjCRN0k4hENdSwTsuuJin9liG8hFpVROOc9nsYwvad7RONN4jAaOFr+
FbZgimcp7XMwcUfn4iS2Iv5MEQhW8V98GSuBmf04zTyzZsFmW0KnslPqtvLAqkTDIm3jbuJ8aYfd
rhQV1nNnriVYBISUCkuwsjT39wMUtPw7+L1nVUvQnp8sEfUP0/ZabJte+Qpr0aG9d7gWScV2LETQ
iEoa3IczB5dDYCRKtjG/O8mm8H8naUWuJyC0w007IBGvM1jjBjmL3Hv5tM/vFIV+ycYBzozVISCL
pQbw9Aec/5CzSR+xdVglxn8nI5pkJUoYVIydFzL7MnC0eH6FTT9fEYcPGGrm4Leybu3gLfO3fp8s
pgg9YnPLyveKdGezELaoT3uK71/Wj4xA6/YvPRwNgwqKSlfvSATq7lIC+eqEbKASyZcz21w+XUbm
hF4G77RKvOq+P73VPfQ0Cw5z7Zi7/1FOE2tsO7utr/Nm1JrpTCTuCSRS7+CaLuvr+D8GsLt86kiC
hDXWJ5COYTXmxmn0KAFiggXttXjwVsqOMMhk+LUC/AfnyU5cpDzeseiPBzodnK2ovBv8lfNKjGBJ
rsc459SVifhK23wTpbsTvf5sSnjgJqmu7GPJsMk89KZ3ikDcBi7owuXuYhhliWPkd4EUV461uyzS
XMmdc/PQm23wIjcuYaY2Z4u+mti+r/OT56XpA1wEh6r5XyLGMxha81nNDLlYchHws4ryrfyCptcu
1oxPSBSl6DejvVhXVSMw4I+MzNCvQzWhfpKzpnb8VLk9G5Rtb61vD3V0gZ1lHBlDU7NsjKm6fvud
2O3KgNtko6LGAGC7+zi/fJ2SHeVAbiBvS+oNuC55IvYtfiUUFvp+xq7aLlGc7Rav/aXvoxHKsMYX
2V1N+hsrnoyEVh5bB2PA3WCFSSmSc/HXlbGwvl2hbdncfa0QH5aONXnp/ljGPczX17oK+Y9mVEY1
y/LbncTSVADZseNfW4JHm6Q4LxwsVEHO9jZ9BH2XZDA+nNZ1DvaJthARVsbnsNWVNu7LTukEkm17
ccEsBD87xIrR2paLWi919/a//R9TuPtVFYIhbLrmPLHE/weqRjQCENFOaxAo0bUp92HRBB0203JI
PiQsyetS3lM3Aivt0eDb7UjnSo27wzeUIrC1Ni54DSOqjo42oOBIC4Lphx3zoxn/j1XYT9GJ9zoQ
fWvlvONneWrnTutRH9YeGUbyQAm537ThqpQpV6P7Y0NfuanGptAODR0iVGxTRggXKEhI1OlSkpek
ZMXOstY1eURXNAsUPFGcDvX1nws1QpmKSBar32WgunkiTo3TGHPthx63m9RaDdQ+zi+wIGKWEECh
gwdDxchdFRzSoSg1MmFIcDr2lc3qkgJMo6LAR7xDvO3y8ad80ALYTtmQIJQnrrTO4Eaw8CHKNa96
kTBSpVhu8zGTwGDxrHl+3hFjSeQ41UxTezZ2N5dR4SrVgu/u3v/eh3IbR15lX4suO6XqdVvIVkJL
r6xRrqVAnp+cndtIpb0jaOxmAEKmWUtQCeNXMEIq5FeoJPUq10rIWcwRIjDBPJVd3wzeAycoWme5
fa+xkAvP3tShiVhyrwGQVow9AlGi+knPCYs0n8b1DCWkvHHxIE76dbDCUlblIYSHIUTuG4ZXD3gX
BTKxyoiFedC2g/wiHddTPgXsvCK1vRgMJG0mJc87xk7c1QZ8S+re8pjY51qVDieCUdXkU0QuN4B/
4DJ7FwwKXh5MYXy8PZqleXF05A39vWYYJZePIKUu+9FjYmJVIG/7LFr1SWaIW8cHasQ9wZtm5vku
wi4rcI6U1ClQoDF6RS2OScHNEUEXU7XlbAVLemOMxzvJqN2p6AgRNufDrkKz75DWqGvxNPba3bX8
7rv9SknEYLEN9JbOWYwFdvDTUTMS6uM5N4z0NxkQg8hlC2B6OMB0JIY69lbGmjhG1KejuszBsPdY
yCkAzGdMbe0qUsMOPj/f7ST07lP+NRKkW1H/hfF/d+BL+wZQ4b//2SSqHE8Otfwl9xUhA5MJU21I
Gx8y3JAbvOncOAvAo1HYb3Uro4ciiSJU41Civc/irr6l0QlTxr7SpXFXl6ft+ptoD0VWCqSZtsBu
+xsrSy2h406FzvhI9xOFLQOZW1Y61y5HryPPw8W2vEvwfDEsCrkmu0JRBAFNZd0T8prTW89HBb63
0nVvs8IUfBAIyhNweC5EMZM7TIeBxit8h9jn5YmxK90idIT3e31Uw2mX/1zoV0Y2k0K/GT9li4yA
ztKjA88ER7ZrGCGaoT1CQ3jW9kxsdoKcRliKI0HA7Jbawx7PEdpBviYaMeq1rbmHvhN3YILnDT+7
MtluXf/oHu48JqGiLp+fAR5NAmdabcie8hRuCk3gbPrq3Dzvvka6Dhewhz4C9A1pE/5Ht2TZuSMK
SHdj7ERY2zKVhGovSxVnohhDQvSfgfYXtLWZooNYZWdFXJnYzKJYex9tCLyYYVE9XyDi+ibPrHCH
z5ttw5kmm8c+oNqXq8frvEhRMJ/DehuXHkVf3gNkfH3fk6VCWtWgJ6TfnTpSuRafZKJFLE+u+g85
lQCHbTwGLcKKNZ1ev/sFJw+L2GLvZeAfmfgsKvavFr8fAguX74ZBiQFpiIFAZhT4uCf9qhbTU7Im
HB0pZ4O6zgtz1U9pc5IEH8GS1IHcxYysDjETxjh7Q2uQGf5v8Rnj1CPWzPPEcOiFz4Ns+Yot9ksp
o1THgQDrC+nGPoevl7kOdb4C4g4VeAKHyMuU4b0ctGWIulncKMcRDNJoLgeAPnXe+/42OIl4yZcD
xVPDYh2FGkYqXmSdstzKFxXFZHFmXEMCw7h8pWfhZoswR/tcP4Jq+3VkzgUOTzGEvLAzf7vxv5qM
H/QMzYYhd5LtGhlAlCepHrK3ASrMKUE0CMfo+5okyh0mYN9yJs72FncTsaJjk32hiOtLN9dHjV29
exZp/PenxH1xrPg3HsjWxmSxUleXLRfCqrcC6rzsPo4LNKTRU8beKaUQjSFt9ao4QSSK2khEYF3W
6P+OVuaRL03NYyozUP03z7WPYYXJ3u1XsVpyO09TLx4gASc8QUP7AuMCnuKii9m6N+Ms3Exc5n7c
D1elVLtXXKAibnUTdD5ECJPdfehy/vjnbR1fn7uWh7k0X9GM89gqeQYPSaQaCybYrgbawyEg4UAu
8hdlvONHWQwJ6IYc+bQc254LkAR3McqurhNX/kRfURX9uoE4K/ectlg4I1D9cc0cQmO7YInxB6lc
pmHb+KsIIOQkf3wIe85DjYdm/w9fGLPU045bONEIiGJa+9p11W8t1XJTvP9uQwvUxyYwBhEQwqXY
H6iUro4YUz1GooSE9heADI3w038ccWsyO72iGwEVO3CFTJTvZw4NpwfuTZ0NzL9U2a9l/fsN9WTb
6PWMQaWm2Scbem5Sy1tSDXb9tDcmwP3EpVYT+sOtrzDFoKKIxxNqWmO8THx0n9/Edl2nXbXkF3Wq
z0L/qtgReklofD7B6PyBaf1jU+8kKKM7298XnpGYIFH6U+TBesMy870cUq9BSQ23ZSg8fA9KSPV2
+cN+rvWcg6TC7larL0lJz3ka53fmWoSgOa/tPy/Ed8MsATy2qeDhdtHz4QkEockHh2u4v07E15Qr
XfZsL5dQLw2wkY8nGTZ4d0QdPMAh6CaPeLMjMb3mfrM+hrFbPgoLa/Z0/riPwZpTdZ3Q8opTABOi
+VKwFKN3n8foO92+6dezL9YpRN8mjLPZMzdpQ2ELLgD6CKDJV/2YRsrc3a2YaiMLcewAAobhYTM9
wyC68T9gmQY6W0unEtWW4Twlg4m1a/MmY5PY8VMY+n3w03YEbiN/UWZGuHsckrmV8FfX7Uv9tggq
GZ8Li/1tfrpW038gO0KrcphShv8MV7BRCanwT/GrYQRjSuIPZA9HW+WYbrk0pPwLXg9xW/VstZtW
VcrgRuybCW6LgyBEDrc6ux3gV4L7PITZ2ba1OdAUuZ2qqxZ/60vKu6yce4n484LUVsN2PrfEfMXp
T8ab/ERqklyNPJx49WFi3jAPaQj+q+w/9cj0X0F4+Zy8X3uRxZjyOEs1x3LBlnf70fSKN6egLJg2
TY8MBcVq9RLT/n0Db7wXGW/7u52XYyxteylxTd4WzR/RusJjs4yZplgecdq7NaStS0xQbhVSMmwP
PxdxI5TET85o0xfIDdmZnJmxFJZ8sDwEaHWIml4GrA+zTwkZ9dwgyKw6RwGNLYX7BVcbQiZmWwMK
ulmQc4k9Xad8JYJJ+LvV4iVqmyqj+lbUqZHTD4SVLjp9ZrHPcHgTk6sObxddTDrRkO2MakgQ6Re5
AyatEFs4iS60uXwdgFmwa1e+nKkKGDKvcPgKLeQ/0OqwICWZRYE5bz0WWZksZq6qqRdM55UHxNiE
4vt3UedQbVRNk61e+HAvIyE+uF5PeBujt4kMPLiJXNJDN5AJOrQROyKn+BUnCUeNyxgO1+uJXKEN
wSEaal9HCOAJrKoWeQs2sCvEa3ma0ENTEdrSaPHCO/5RvWsrQ0jK7yW0bHZfAPwJyL8tiOB52iQM
B5Hz706nsRtv2xPCtbH6+SD4nqU3zlB+BD98BuFU4iS/3CyzZi1q9x7j4u0Z+OR38QHKXV7VCqW8
l7NzuxwX8Nzi7L8Ia2TslHyTQKshMo2A0LeQhBRSDQcgPOBtrfrNuIEGbhLkJDs5z1/t1YvyMb1b
jAcXX0LBFEMrkneJ0HebrgklXWyufU9BzPQsx2KGuNsvoazfWMewEwdXrV5E/V3CTn2jNfkMGIwn
o0LryEi7Xm/tzzkGj74eyj3He3kiy2zivA+XFB28a+cZDQGKcW43V3Yqpzc4ZcJMktBW4Kuidwa3
0Yo9BGJIbfMQXM2hCD5D2gpm9Y8bLI8I6WxeQiSJgL0hh50zlqY19R/9k8cBVQcNRz7QlBlC1j84
4/wd13MUupIRkM5bYR7t3WA3I22KEj35xg+DXnuwzpgkwkJliYrBLNaCt4hKiAvXsfb3JFJ3b0j+
3IE6Ke/SVaORDY75OxkJx9HC28oG+dsUb9WTm/tm195mFe3x2A1IAx13fwIdZu+et+j8ejsPQMco
X91bAHfQCfRlh9hr2NtRSdX+BHm1cuat+2xVTn2fayvRXUX7/U+JRzoLP0KyOpYFiw1fzyiRRMTk
UBH2qd+7gu09a/gsP5dJMleXhP3eXvPZC+Cih+Y2vHJa9UbWzQv95gNboQUv5ONKKM5kmb0jhYDW
LjgwP/5mxcE8JFSevhVhxQKJAaAzC1DFZGGH0wXYaC9t+pC3o8Z4ne9ug4h8sULHj8c5raizBX1x
rgQlWkxdTiGn7118Yj9NXT7JSCROllG8riXkgQsudFlEVBfR7NTkfdIqLSsjMtS5XDmw9DwvxAVU
oqjjbLmG/5OYL3CCZVpO6B+8w3nUhVPXZRMx8Lc2LZB8bsQ0OVX9F/yvExK2Ab9SFVYcI83pZPea
ABHTXrUfAZn2P7spNxxvmiJf9NANkzWapi1ub9c69s+eu0j4NKRqI1hGLyIPtYLuDbS7RS2iF5Yc
aF2Y/ynab0/vWxIImb2ooXAP3KaorQTadORVNEqHN0wU1oWoCxbamR5IY8GlebsYyS3z7VZ/4+be
PahDXp5m+dAdIoO0zLLmA0WfpkDAoYLcx0KVi7ojRmzdi57U8/Z9LKyAIiqliRn9neTE/9bLWK0B
jbCNgUMF6xso4sdK1TFP9kylc6TmADk5kg6x/FmTjx85Bwqq4nK4kQJ/nLgUEsl0U1W63q61HGOh
dXsPcMK+z8ovm9jpUH4pM1g4t2R+AhFEyboZMeENp/sR7P878ZxEhH1CGzGfszu2yeB7LiXHCCaJ
cQN32DJZQd1VddlW2Yhq6T58PPFhzA3lQQIbfi768zpCcaQw/mCLmxr2tCTFky3Kr7jrUE4S4861
6Y5ZCNspt5lN/QDdxlg5VvwnbBmCQT7lx1wjYZVouJSZ5nRJNArY0jJcueWOv+LJ5EmhIU3/JUDp
p0AgJhDiBfiFTRqbUaGqlLzjUWt8hGpMEnu9yptPaN+P6lHf2Umz+vGoYFl6L5FksYo2Yo0ZZ390
cRDmFiRs31yJHq1/grYmBJ3Alo9Vf9mZ6LRW22NKqB/kaidSPVnK+ztLmv2GoC4Q+NCawNNw2nxi
bMGjMFqopqyhzjYVbZpm1NEe7VpJXc/VS/O3stLYzqmidDmVgS12sYEG5MyMx+F87nOGwAy8vnr7
kvnYHJeW2JQND8IfSG/u7/JxwVp8I3PvTtaPCe8+Jc7T8zWWloUXVqiVma0whmZAUBRqUNTO8pLc
1sXmJKZG108jEr3Y/zjHzR4d2pPJ7ijbcozZoWdVYFy/pSq9LrReX86vTmNw8zORSCI3GFbUkvhl
GefdIavaMYTrwLYnzHf0f5sFvW5m8a58p79C4l+2pE/GIUghrp/WFbV/swlTpppz7EwAhscU6vDg
i2bw9BV0oDq8HyZQUDLnn/9PKmIFitybVNURlBm1n8qi/WEb4GyzOf3uWE6+9SDbvQwtpIIVImWJ
BQWtFp9q8eIFIpHqh9/C3puEgWtX6oQtCmo3uohVbc9+a7QbwAeV+1t7yr76zetJrTZ4Zfk/HOHz
DHjR8VallHdkyT3xw/LxRA00obcinGOuOzrelqwJqPAC6Yq6PzNKfixleh15cdT2AcNjBWqpprwI
R1w41814lD2fUNYdumA6ObQYWpUB07xFxnpsoQzO6shGc55ii/rDFnwA1UmwGw+aQj5w0rvHGbdj
N8+ArnD/BjsKYjDuL9R3AB1C1aUeVlHXFDWHKxcoGvtFpLqkAmWdsbOY22DCwVqedLUZOhWcdg9e
aKonNlO8jEtvTyTFhBUkj3VJAq8L256DOr5Ao4RzGs5AXORHANQKCpimA7FrLjDgLAGddQJrD+sZ
3K5krWZoTDM4jhHOIMo6DuPh/L0aSlh0M7ZZ2MBdcQOsTFc/geRa39M9qZIPY0820q8I/y8EBY9f
JBKlPZ1XvGWcYANnRbAuc0kcanCnDuZ/3zravixMCQPRv3ThXsiE0yJVBP5dSUzKDxPzlUfZnihV
Vhto3MYt106vnZZc/eCP4WnXreQQEFN2AcLQn/eCveEQElqaNaVYceHwjdCa9pveIUlm4htCXE9i
Dc34CIwXjzimOH1QhZZy9yViZoF4rk08nleEtZq6D41lmhpe1UL3yCe+GKkV6roKTiuj8Zp5TpU6
Dq3RlDMuWDCoQ9zM3/gLqFB00pdL/f2w5pyjbj+OzluAGzmwRgk0UDn3227b8vPr9mTfbyaPZnk0
o8dQggE8pUy91UvYX2I0giuzrbDlC56m4IT/ikNruqgvYxXKwI4cXL33Vd1/O7qCUJOOOl7aTcpE
VRmx1ifqI5O38n4TtmXznwxagCNsU0wYUmpoYggTqDi1yPrJ0/UZUvDhh8r//oUWHzDHWeREK2j6
utfZZWXEB369+G0DaZHVSYVqKDjU58iQiMuckfkVf9ISt+HSMosAcFkXjKpvLejZE5ZsvDOLiuA1
+jq55itkqtxnYD+6yOcHKFAs9YXsvqCO3XJEgydRGSPMY9sGcvWfLLhtf9LjYURdWNXHlRWXziTD
ix6qkhr7/pi823P1pNQiNFZ5MEghwDDCzbuezgwbJHE6tEXZLeUrOXyTP0+D6ekJ4Sz1jQh/cc9F
+u16a/GlaRc0pOSeD44Hqi/bUKVHkCcIpTPAydMYRzY4X4Fju/l++scOnBbaWCYCiPh/bF8MncTU
jCoJGcC5YAuwuMs2Klx2YujAbeJYMBkMvSqbYZe///ajvrM7kuAPULlPiiHnQY/imI2hmefCtf6B
DXNnIcQGSRcQjrrywAfh8hyoRDiyiQr/ZRULlPDtozrcKMKFDQmu2oJHaQEQOKSD0o4CsfE51KbK
BhpXernpXi+EKqvj14KYYYIVdAa8FuXBWEOVf6ZDbYgAqdc+OQVEjkNGQJhPgGjY9j27Szw2/WNw
GmUCfhq1MTrLuUYssgmZafnbE+GS0Hb/FIDDrHi1ZYksh01ISVQglQaz0dYAzFs9Tw+hLbDxeqRv
2BWDNlrSdHkiWI6rM6t+Nb//h+gBMJ3FMs1VI1MjmXfnUTXvrHfQojGSg/qu41Y33U/EeJFu0zMd
jO9iG4Qd5tG3VLxQGlH/n2e3m7us9caP/j5z2kF/NU6pl3W2m7B9qZqAhFHJGDHHd1ojClnv1344
7yxXHkiDm5P6JEroJSJE9899gLCulcC1IAFZuYz/3N9qoGlvvj4A5duqT5BFLK8HjojzlVquP2Ih
6AzS5qDUe5xGRzftwagSK+/WzZ/o1iWige/vkk42OknNsRWb1niYuAS4MT96VBnRB4D1TAl/wzOI
pfjB0uquefW6KkF3zbbhPnIfXZuzbT38mwrAhl0itKDiHIJvYu6kLVhNxm45iK0wwV3Zdz7r5ZIG
YA9w2YghU47/E953nV/cQ83Kuz7GVZ34qJDUHHcSU/d/ZPySH7B1+a213hQLb/hici82WUXES7c8
25lGCiMDTXAA4M7/f/cQRUjtMLT+OTnUXVxD2t9arujkV/hBN80eNscfjQrC7ZA35ovE26QGCkT6
WJG8ZaRJgPukKNmFm2TlUefFAo2NSstjvxBEJXV7zgzvWS0tDfc/uSUnnxU86TtEEpm/xaglT/8F
ZF1tRNm5JrMnffefsKmmuoXGeQ/WMJnh5QUCSoJKVO5OiJa5rhikQqGxhnxjy694RPc4+UVlmu+/
VPi5l6R8BohyGaVwLWIQdVgQhWqLb1hDsFKOWlyQFCYscwocJWalxi0UH41s90Cyu0LEJiFMkDrk
6vfM3b6CYdZAZcaVn6W/ss3gsnEw+mgJp1hFPl0RjHqB0aOkUsOuvZRYRASM4cZpncag4l56QCAW
uuXFhu8tUzMqW8m+sy1Txg6pHKOWT3ArvreVUUc0Uqyvf0oTqhcHuK70FbndObOHa7pDssTkcuU5
oquraUvB/S0oyelXQwixlZWGDYCVDj5FYXTR0CQ6DAY+OSjSPN6R4IzdQ5OQ1lApn3BDURKH8BxL
/R2rCfy/oc46fZ4FQaI5SLLFUCCIcUEb158wVDCEbiW0LkES6BWz4UhNCcWqCLkWWnbJwdoeB87m
jHKGYQUDJuNFtpikkz6FlKbXBi0gDcfY5YIJH34uxrcgRoGlIx+ZrqQaT1LVzEtskB2ytiZX8Ipt
CQdNaf9Z+X2zhv2N2oDJ051x+eCVgada7p7He6ViflGnuZqXzpH0/Ax2PGm4hPkebMbsPRcwDjzH
k1QHmFkh/2E0o9Myx1Wh/kZRCjWUEYhpPlnOyN+Qip1wiRXoPgJjR+4OO4vFSrTwbjn5fHjcpU2v
9SUtqBs9vXYeRxpJvawzk573KMRqm9WoVxq/t6tUsWoTiP3qW7giu8vGJhPvBL4nETPPAtPgrNfU
iedeCdcmJzKeUM/PLF63Au2Z1ETWzKgzdK1GHvoCqW4YQc62Rm9UEfdEg1t8P8pQrEk6y2ucDGPw
7M/pvrKs5nIDWUO9n4Z4xxwupGiVFwk4oa/UMxVEcLlCjD5UN0k1PIxlAvrt9Hsn8HxjQrFMxRDh
3/9ayXXrYmNg/IJ1UzG163kNtUEhWX4+c1EeeY4ny0MhMb01tvLVB8vQynDXGWR0M+mifSBNi6jG
gQf/wWPvb7+kT5jBUcBvsMl6YZ7kXVdt03DLIAu+9/e+aELK5Mqw/wXDZO/2JHG0Ml52Vv3PQVrQ
2zs5pSiEwd/iAGV7nGHgmQgylV+Vv/KxYotDJrgXIuKHBu6BahpcVcp+gjcN8SOwh8Arr0UT91DD
xNcw3Xd8Z0tNRjGWb1PWN1byR1QJDrS2IM6zDYPkrJ0DQF5G5jP6UxND9W1Yox7qMxHrisLreY2A
2yzYWXwm5/jzj50AFk7CC6WI2tlJ1dbetGpygjsZ9X75gG7YV9AzZdD4CFujLhRDXX55Cxo05Zky
AxiqJ0zZEVsuGnx3nNOAF6i9DtVttMDxwy1R+X+0zDE704SKxa7US+/hV/otzOedla3ax9nlBsl7
oN1Rir1qc2YnQPcwleWg0e+gpHn6guVJZFEj5ifIZqvNutnNDdTPfxnL4BKllnaF0ZvsWLBOCTpH
N+I+TK1fwpRf3ogGkm0SfkyhD1tYnGFBAzsTOxFBfAyM8olpTPgR3x1ILPdcdZnSgcVPecdDtqJk
uBsj5ILIMJpASovpHeyBwblc6sqZlb6oUafGjFwzcKoK/koc5AHHhSxTQeIkQkJlDfg0U/I1sZLt
HLaWG9iYmngnHidiB1DbjZBNU4KDg10uPTqMOwlPy0IEVImDGA67V79iB6mtDZYgQrw6jaBpMW+i
qy6fED0iSzN+wzo/UNw8Fi2ZtMIw/X8zwHTyccSvCy1hZT8PpwhtRdJ8F7+honN7eTc6Ebh0Lu6i
u4V7CVadVN1MGz//Sfwyk7xhpZqIIJI6J8kaePxoVRYNagBzeHPgDqgQstAiHWitLpIDEV4oAzdy
ikRw1qW0Ibu5YnNZW4EvJcjuYfjsbEhxjwfRLKZIi5dRoIxVkaSt888IulIOBp9SHpF4xYOSn9Ih
D32GC/jlf8jxJQSCsf2hkAFG1zUfF38lJJKpooZ5iG2F499vy/1F3hbZKktWvO33+kPPx+u60XZp
Wtt+GR1QXO+vO3iWloL06beN7aEt/qxBw6qbNNNAZ4TveYMezQmvkBZS1Jmy2ZG/4k8RFBu8QHqV
8r1TcBH4nyDHiryP4DlI+L9j2QeuXishM+LHm1NP+gkp+N8MP5Tu9uZaZJFCTGqw8MLzI/V9Ad1D
EyYmwGT5T3iSP78IUthY7wTt0Gzh7nFosAG65bpLXHN+L/8fWdgGmiPFe5dTRlBXFIaF05N6iHJm
C/13qf4YA8kLQsoFjE7WXqRs2JMiNcWgOrB+zdenkpYVArTBDSVpA6MKELj87Q3fKwVUgqrgEfG/
uPSlqjFxgu0aR0TC02zpaGn2YzWMLR8sS/pTrCS10xQonK4lnK6xYpyGv6w4+PWv7CKadiLO0HcM
45WqYCqqmJICxVXV07QqXHX7FH3JkK0nJlDe694fn4R6Zbynf7Leksa/9puPsSbqGv0e1BOr8lsN
2t43ExFNm4ys3/tqQZXKSeddVLF7TxD44uSpr+N9LK5yFVsBgtWpmRvCQkPEybYE7dkpEgb8gdH2
BBajVMmPdSci9epNTxwZPW4xwZFbznvPYS06Ukqzoiw3RUNeIvOZ9Dm9W3ERY0ZCT/Unl8b4lT83
PODkMKsNN3GsZNykdSohwFKRcAWEvBAztIAYPJ9v82nHYThD4GTyaaMPA42teJGjS21l4B+dCYoe
LlWEJRBpGnQW905mCq8/nbqrcL6kTxq/WL+aeeFb0zW09DAE+GITLCKwmZsYKigxh2+4f90iBBig
aCd+UuzmCun8K04a8aIxTudscnhGGATqxArNeR48rzz+Og1IxPsur69D9nGy7zXcJDcaM8leucwO
5j82vBCQU1nyyiEmh6lO0eEE8CumsQ4Fo+X2yegYVfN6CedGXYckOePfS3Va94aWqqMkACho3r37
FDHf6etShx1uSkQ5fxe2zSnKfO4XgnOuLYbL+gfoIfJE3buQIkRJcd5Wk2Uru9cKAC+y8u+76C2l
elWp9LCjRqbQbqeRHmHWETgjmGJdxhHmMkhGXLi/O2JEULkW0UcZhDo86ZMlggJPqazIA48Kaub5
llAzMy90uHVPb3Q3ogKXdwrr0lXyCP3p/2R8nF8o6YFYoga3ekW47+MxdVqm8W+u3MOobBhUteJk
7eY/oBl+qOLq1WNNIGCSg/ufPmMdpPvhllKS94siddOehbWD7MFob9STXi3GfY/jU+FfsogPBUmU
HYX45TAmULR2laocGaKLd8hmdkWMRJPZ5b6esO4ydEGJBWYWSLucM/eEAEm31jnBfPJqy1rkcWlB
lVgWPt5cIRne9axQ2tZTmk8yI60l7JDFaYK9EUAXkfwEgS46WUqqIWIWW61dOtsoFdE+iZPj1Vty
YSXdVDugU+yEabSD/xmeJ0XFNqmXDihRjd66nF1FYklNfBo01sOAZ2N3I3Rfi8AKZHxTXrOdAijj
TEqB6wKrbD4r5/wa93P+ZzKwbhEoqM2EmISzoxfGjh+bIG+m/m05lsvpJmld90qAAJ3kUxvkTJut
MgHHUNJc2a8FlW56hTjajsubyMjudsOzY8W7pegXceU2N1HuoE/WM59ueC4SRZXrCPe4sNJ/6/hV
zTpuUi4cKx2mk6V9mnN9rugmp0QuqgQtEGu59MkibJuiE4xj4q8V3l2Q6+huSwXUauc1+HjmfFAl
y0YZHiQCaXmU4+ONtR4iQ74Fo25yf6dplmNPBJZmN/43EsjoUEutnaP4ku3lRN3Qosz+oi51j0YS
l6NQeWYUCeek9ewGNTiolknqTq59AWTYTBsAl/yVpUGOniAoBXzoa5aWiDIy+n5uzlOv0mtVwhd9
KFRSSKx3BV3JWks3La+7YaNSfD+gM2NEZ75t6C2wAZ2HRmm1sECos8ng4FVBhQRUlWjXDD1RK3+g
BxuWwBvuizJVJGAq6tz0O90E0S2ImstO45TOqN4io2UGfd1t/Q4fuObafchjE2ffmi061GsbZys6
AHs48M9w+1XfUK0BK9NUd+Z0lBjCFMtXSwNHGXHmTPTkekGQ3uhR9ELeT3rN18iExjQr6Zyb/GIH
UKh8R1rTY7rDhMyqRQ9GVkikrsxI9l8efzkRv0bapBa0j9BBFxJyzwk+NTVNIYxlKWNn+knZ6B31
opEJ5w28ALcpBTV2k4cZEIbm8FYj61bSXd41swRqZwcTqC+zDFs4MMrHu1OG4b0RMbGXh8sKsikk
gcYG05OVafI80uEzmaTATmTJzUyH4viNu+eCXfEXHkmwwwWNdke00mk+98Q/QTDuM8nyEGL6wvpU
ufIhX62xPjZ1yAwiEq2DEz4BQ/CaVDEZowXFcL/uMc/kyDSCuwvmPSAHddhXN2Mytzue7wb0wYTA
jIEjY6WAqreMb/2JQ67JtA+M5aAkrxnJrmCAFtgV5NGdouU5zcCG9H+hftLlABukM0gfwVJx8jby
c1KOaF6WVO/ItbYd8qWMDYsGgVSYnGtDlJHtaK5BIpOQV2ExOkhRmZ25Iv2zb9nP7nN7o2NZRnMf
QkfO+fKUpjHyzfdyYak9TaKTCQW00zUIjyniITwfu7LJJsMSROEj6Bs/Vavu+gQet7TdjAe/4TBs
XblJiXSxu/2FyQzWADgOjEEnwJsd9FCDaqfgl2EWwlo6u+uyNGzIF0BpQAFXSPCSfdN7tz4WDaey
8fkkkscp8RLOImUy9vu3yQWm2vW30aKb/KGVcxDyToeJMrjcvpRhCFZWYnFbjnveC/k0GKf1M4kb
RM1+wMAkKVVp2UVv+Hj+R4Zf1UrTjMcoun2EBgDiBRy/pu0qIlrmVjyrd8D44jGG7ZSKpN28C7VR
lfcp/J370vVdofY8n0eHwsjBxUBouMZZq9EApvXtb6Hfc09Th9i/elQCq03YGTz7vQsphs7Yx8nf
1+x3y9Alg8Q28kkUcMw7H8+KGU06Wo0GRBaw9j6BfKC3PEkiCr+aDOl8JC7BfFfrTyTRODLTsAVX
EPW3GAzTAVaffP8kMFXPO9Lau8saMqArSU1A0HmjSn1CGSQwjux9tZL1pqbl29/I0CIFo6PV6h/C
0wOPNCv/FGZolqg5k6VpDKGXPzA+akFraoX5Kett44hAc8W+7iHYPZ+T5jAIHLe47E7T+hj4qb+k
pbjw0Yz7LJuDaoKRrVOGNKqUxZldQdNEXx/LenppL5QLv2LxsatI5iugZEW2s0V9rbLqtgfkngf6
eNkevvFSKEur1iMzXQ5Djv6Qvn466vsCJVgf5CWMBPZ7IezNoBMa2k+hNLZ4+X7Z3DrKSyqjpZem
uELqVc2JlL0KYc7VbmcWuP2ditGz8Ma5p2fzqnuvWZCimt3bksb/FpFsJm7SXSo8PVyXrS4SMCuN
iHb+uTEgkZNSAwU5Iu9GL3h4p8g1DgcbUU+HKVPo3zibVJdAcfGhNkTjNJf9Ungyq/0PuxGlViRm
OGE3c8U7vFzQ2wSWyLADHu3cfw16VLUuaSyEFoAoGwnpTPEFOY+9fUT7K3XA+3967s+GF9ls6upZ
lY520oTlwBFukbFa66xyk8SrMJmt4bfYlwDKyKY8s+jEHaXffUOx2IMG4HUse3+t7SHOcqYF44oa
h+CbUG/93HEwoP3oZHpifOPGlnT6JRjftqEvGWhUOFY7zzl88VB/URh1Y/UFekMJUYuwv0lbU14j
L2CHcbaojLxggKWSOk9UKrVg2RpIAqMFcdvbZ6Pdc5KbjoG9fHllkrj35bUH7bv9ZUUcB9QDfuHr
W2XXLvIeHoXOp0Z7qcsZUR/oLbgIZGendaLNrcHv5Mfp2xD1yT77HZmuYZ8IzrebCRBPhTh9DCuC
thQBZ9J9OBXValcqOFgw07UK2pWZLUysMY2ShlVK1sMzZislbgknMxWV/x78vXKITqKhjvf70Zkm
8M2ci/k6JQ7FXzBVV6rGXoO2ayE78ZPfTtm325M5rPysyUTyQhXd1ZbinzboatYREsB6DHzFMSkr
FuZ4qqdmJp2JBdTupCPBetkn4rar0Wdu8QtWTEIeBCminWvMBeA5OC4zWAXA9U2urYlB18ozx07b
YI6ee5GHvVtZxl/aW8YbgUUgEETYBRSAhbgi0lIFCMYiIuT0cC/WLzeMSk/Qv8BPcvH6r32jneW0
z79RKD+ModmcWk6xlAsYaGgaAZ3QLJeqQ1vZbrR0TqYPX9rr7WUqBnpKtWMrQ9Nr7rz/RVus+qzj
NFcy3Tp75CU4LS4cgRIAryZKb6PfOcnsenD+VMlGoruATW6k7x/uE66msswsjPXve5Z9IwXMTthi
C2ypU6VbU/P7vTCOH29FxeHEEUsWMjLPk/zkbjo42PDXSt0xNTuhzWukkd5oNtInDmlYJFCsQgNw
fzb2K1KQekRq56nWBgrTjLau6E9r8CpOwvZW3yXz6q5/MSQKySVGkT09HIMgBxHT4bUykW8XUdae
c5tChRn7LFRd8CqXhPj3AQHZA4w3ymGb3z0VhqVtq7pN0w99ktyR7b/pUvuElzDPaBt+cEWMhTdr
R0MQ1e1vLbIy7D84w9sOmilvf5tFuyatKQc9UTLDc3bpfLrGfYt5voMbhgF1CC8QG/WA5l5ru2Rg
wxAre4J+TgxUgNpg76hs/vFNzoORevMy5PdxaSPg8GyltePfW3MD8he18IHGSIyhMTIRhiWrw8Ag
++EFMW0DMF3XTDRcSXb40l1Q16uAZJ1B+l7lBlhR773RBKkOQmF3CcUNUrbi7bhqNSUaF+0ONplv
NRXXVN/gbTwyjbnrmrzT7xQgyov9EOJ3HVJqWqjFUkTbzdqqcTQ7zJMh8Z3r7YLVUuCEDdRkUwKn
0pSO7Ui8/WSRDWQI4xqA+IFDgPWztKODMpHRgjOUkIMl+T+8IC5RIZP21BCqDpNBOec5gq+3Y1HB
QUMAm9glV9pa1lISqRjhELutp7z9sTPcWuuB3hTEWPd2Njp5+PfsxnijCBAkenqNKUaosyVsEN8e
ESFlpq3N2JmNGKKfp1gchbaawWqRo9HKqTAYAHZr7JUmi27KzrjS8IWxAM9P+5evmR3UHUoj8U6d
uFO2q+jEFABhl00oXpa6N8C5yM6gB6zxKeaWwRerr5itEj3HsKwQUxVkyjFX4Wuqyzz2xfAt4Fqw
qoIeEYMkQheIXqlsYbnV6PLxzwFlBwM2ceY1nnn1u9Jg0MP40CSI3dZtahwsuRA96RyO3NBIZ4Is
G7J3CTQeUyb/O2IMC8xVZtO8cLLOn0iKGyzSvLE6fYzEckLlS/K5g4JZ44XvmINrE6rsmzJR/9aa
KCOEf0ZmYEhMkNWAbB0EbMB/PhbbvqrYPXSJ7Aa5Vui7TnLwetL9hdVIHDfThcVTAsn5oLn2TtN4
2CLO9cEp3eeQeRMpZUvOpdRsZQB4zag+9vSsdYg9SyvjWLy7aTBJSLr8pxOS6HstF1vlZSP9yvhE
+oKM15qpmBn4y6gyHEfuw2BXaG7oMVZgFlADJVFGULVO/uZJsktBG54vkIEXDoSkuFLDZIM2I/k0
mQHN84fvvSodn7G9s5wvLMIVwYLlqQEbz65/at4HuiAR4arLcGTIqtepTzixKjskKXsAuSI04ai3
azj2b9pO39jzMYhVm/lK6xCpDJOeg9P8H5HbfBYzRsCWZqhWHsVUBk+/sbT3rjfc51hbkQDBggIV
ELyonHPLZWQkaIK5HcbuOOEqbTWWVOL+DeVItfm+lr2GhKnPx5c/92Tu1By6I7vNWZomXcj7i+8T
KULhRndDSRjyre7fw/u2sgMm6e8eoRG60ltPG7cLNFbabbMgaB6VdT1gigTZ44iGYWVoCmMSHJSu
pk9iepdgwZ3DWrxa9FdI03Pbf7YoU3vto3HhHzhW8hU/kVQ1gv/1Nv/r10BIqO7URnMVBPwVglKj
z4gE85FosoitVP6ieIj0WyR6sj1HULLbOv0QwBCstavKUcepebE7d3/PBtRJJsI1NLUvWOppJ+Ut
iCCbCg0Msrskhy6f3D8B3OmBp+mIJGMMLv2p3Pz0e8aAxd4HVdvO1hgplaZk572bg1hI6r7SeiOA
6FD0DTPbqyv3K5LBsJ5Oo/Np6+aWYfbBgyG9CwN6p7RZNNTstmzYxvbpK2Q7672++e4HHmd6EirO
94/u80Vckgjrk4q8cdxcCT8Gv/6b3xmB9nuZKPSQXSIzO3y08o+rcfavGOslGj6ebQzeL1U60FK8
YlGdZdXb19U7psKZWrOd+o+NV8ryyG3sAoXtgpwyJ9wPHV0QpO+/71foDDSKEKpZSklP63uB/UED
5hlveehlh6rapocr+e4S+adxOzMLclB/uiMk0r6JI/Ey3CzM5CrPJNJ208jOzqy702rBpyJ24eHU
Hklo2zy9Xpf0QXvxtNDDi6EpLw2y7E0OeUb/FG6ePCGSw4on2+jDVpNKPyrvpfyfn2oLeZMuMBEZ
HO6L42JQOXNBCqbyACv4k+B3JRq0XinYDlMZ+DlM/Cx1+xLRUcCLlWVWPq4Oa1ghjJ+SZ2TPgwKP
3O0hgnJiaFnzh2t3ePoF+V5UKO2jde1DDNvPe5ALp+rhlkKK81YigYyWJ24PJQ4ZY/coA+1XX4Ui
i5SCfFZHjD9rxJNcBnnMZ7LveNAIbOgUHUbAZXKRJIZ0XJmjes4VMnNGGprROpZ4x4Hr+3tcpcBo
EFTpTw3QMi0EdS7EN2R7rWSA1rj6vLVWK/AeQPWNcNZ/9h1VHTzdZkhwc0Yt1DUg2aFWbQJJ+sAC
2iXFZu7q7KK5B26jBPQHB7WtBzsg8Bs1gFyEvg6ych373daOXdu14Cl8FtqX2YBWGNgGDvXgpm+J
2S/wreL2vXGVbSD69jzyAXlhQhbWj3OirVhlvvx4btJpPRl17cxPvmSNXegudJAqy6CyhP67YmS1
FTWPtWgkGRXdqA1Powt9+HY89qeIJjr4gDvSFqi7LA7voSvjWvw9xDvg7ITI8Jf/zEisFxVsZYj5
yZEI/DjnB9hAF6BO+f/LXUoou+7xf50RxzZS/6UeV4Hy1KGPLqOq4HhNHBIjZsDOgzzeaGMGsLGt
MyvaK11izdjFoCDpG12f+4DkrXgVnpaKyQifrkpSml+XmPHeTKggLeAMGa/WIJj1x1p93UPQWEJz
2g/I1BCTWlxgYrlsI677Uz3R17CV1Qq+cEgHwcILG3BO17y6Sd97UovwpX98BvhjA2eWYL6t50rS
9P9K/4teUiK+sqawzpbrqHmdj7RLL0PqAys4PF13QM9g0C4TbasB488FQgeZINgkA2+lwg4xJdMr
KPi3YSa/9KCqsUASARpNfsDSCDdoJZSvh9i/OkivzLVnn7UhjTczawzTauxkfsTzRQCSnt30Cqmc
3HuegwBa5yrv581+elsH1xSfmbUELGXV0OLfecsI2BD9gUv4KA9j7LBgDB0voBjiWhI5oE2HzNfr
NrCXTE9zC6PN69teuXHEOSB1pDjX32/W/Xwj0f7yD3Wx25WvQF1k5kY0lRZ2ndNIjseWylTkE2zv
CLeH9OK2Ns5a8oSs9F9Zi6Hk+UmTiKyt/SvBN8ZVy4wyrZOv98GiyvJ2c8F4ncql/usnuUPBu3Gn
dzaaP3nbANHLUEu6zTfCqaiGQNwmmNkAnrrVOOQdkSxQnFKzvm+jC1JD4sPeZUAGygFfd/NWKyJ8
4Ew/RCnKE2+HFEQX6GjmeynEC8NsEKGWuX2TzaRSMRNc7eCA582ldgbvcKDpnXh0xkOxVGQ8wpLg
HnWkJZSIh+/oVtM427f2i40yLPnCUmsnS7dDUKIsPbP0kpn1g7AORjP54NfQHuXavODmzPUh/WcE
QuFEDpFzQE378k4TYmSB6qG0N2dXIOqAM52fZjmGmLQ3vchns7J07o8P1rpZ6KRN/u/BvR3gj5hl
pDeeLWVUWf+LCEnHordIN0hMvKqdGe8zOitl059vRu8E5z+Dkx8ZCX1vcoMG0x8PBP6hIKAHBLI7
WYL+SspwUWlwEMuJU80TPoI9iC76WWE72zqGDtercd4r95jJGkul8yCaARCVgfuIjWQFMrnz3OyC
OXrlBuYPvL/40c1R8b/IjnDlHF/YVT1lYkxuEg6pmyWIbQZ9jksJ/O+X5JoAQp8wZ4i/VINVgPZ9
OEetqtmzZm9IK0xRqvmRlD8q/zQserPfzvCzhYa1P6mO+ZisdC3YLyh4QGLopry9+8TSfUp0QbWl
BZVGJJ+jLFwGV0sZsDAYAu5QIR3j7zN1Gy+xmAuBSTs+LlmEl6yEzCqCmUNZWJ++HnUGtnxt0rSI
adktRRoYGv3Y4l247BPru+txGDFbp0i/uA20Bf3sQ1v1s03i4n8bdYvSd3JZSXsx2dfaWSiis/y9
eZ+RPz6PgaKZQUzC44JPiaufixzCx4zvOoVsNEyktU7bS1rRf1ndfVqKn2fgTpIJnx/3ZXDIac76
krB36A8d151yR2oqSUNDkXwZB8dslBtydkiAPB3e+kT6rjTJeLaut/e9fMWxqI4IIS1/yYlhTZdm
r++TG9s+NoMn5ZZcdIdPP7cvXWQZ0KGok0Jmd7NxCZwiVOAfpRUNiLr1fDo8z/wM51HkBwggf0tI
ZFOWjgFy3wodLRjrQU0Gx5vO/TXkzywn5/T/Xsyf4zFpnGhHAKTT3QyovxvBYVLjtEihnfztRhKO
xLVBFq2EKf7fecnsZSGpJSk0QgnS4gBwTUfNTNFk5UgEE9YEzaoZEO6u5O+fVQQ8ULB0TWs/W58+
LdATD9LZTplfI/2zr2Au6HTlNPba+T2mSxD2sG9WQfYFrE/VOiBjlBVhVz/psTfCt4miTdsXsOLR
A1nwdZKdSHv8eF9df+7YryMzfAWacqv2GiYqvmtQQ1XUewq09mKWYZsxD3Q3Zc4b1va0C9kpvuIG
4PuJoyRXNYoW39QnALdsbMjCsGvFu+waezSSWvYmdYmhKSR1p6jx/ngMksorwiVQpixE7A1EEP9k
dvVuyBZLt+a3fhtIVjbOEKBU5tmzxCaInwyKpHG1W6StoQ0q/61pCNJNzsiUARkB0sb5uQTJfrT0
oBp2Q4a2jc2fSp8kbLEFAMOdt7GlKhUGeJ9xiRRNe2lFUlYHg0fYzQqS5ottyfDi9e5Ye4bqlzxr
15nKDu23FxUE8T2KkOKNuwzQSBVv1x89M1vJtFOmQndYUNpdb+uhIe4Gqh0I/qglJw1nCC+KV2mb
zGV9GTNCzOgdhWkeu4s4SZ1Pmv9N6T5KrhxpyeQnNi2nMN42s/tGjhAIDzgu9Pfn+2TbbJbcktQK
tLJqWckkkMCTaUqR3x3+oTrrnqeKeEhUQx+AZlUZtxIDkuN9Z9cw7CZPKQmVQ+iUL/R4bKTllpd2
jP0D+uBwBvuIJNpkpe3cK3HHypi1N7hQAE2TY/fqsGusnw4xLgq3uMs9s0fRKxAMvXtfs9EDbfCB
bMJI5PX160pzeQhwTFXP+s2Szukojlw4LE1chmPtaNY/CzB3R9JrOSuAzSNQpEtD8a0KLTLRuKHC
yDAeCFB+rAJj02tgMpJrs9eGpcO753PsyamLZy0QstA25qG1Qc6nkpaD3jPsEBOFQp09IGIwU9JZ
fHFelGz7kRFxQ9Q31N+C1x+09Io2k7Upx/AxY73YNjUk1NYQDAKwUYtn4ux03UFaqg+mddmxgGOe
u8zQ8ZU/OV20S8gynIsp8acuSM2ECZ7rzz26CmSenLDfmrVfAcBfSHRWseLJBDNsB5Zcqh5fEV1t
IsJn97TsNtPzwezimrr4MpNYXjev1xt6NBXayTcZZ4YH85+natEsjHfvtg1aUnbcYXHjN4QEe8Hy
KJAJFV7lr6/J1Xq+i6WV5CajsSICszy3W6Jstdg06zkydXvtB8ffEk1gjJH2ECfbhStcfTtMXaTF
xTlVbtNZhtWW5uhgJ1Sal8JAAkAGAflJbIjNjwyU0RUIpm4c1rGuRA0Vm+Km+l78qTtZy2LzUA3b
EngJBht0pngszlMsJSEtAN68+cPkreH01ywDhMpWTq5kxU2Tzox82EaaVV56yPkcm+9WYvIDT1Jy
Uo+WIpxnEwX3enwPqs+xWKq+ns17zRG/0h+G1kd0CwlZpAtjTcwQB8gC3JU9iCsk/Am0F2/r7lEO
cauS3drVULEW1QaIiKga2jMyyFI4IMpM5iPH/mxfx1ibAdhvOJwgZj6VXwwf9cLcHMKVSpASwYE9
OWswT7YpfUICiZcE0OxsczcZ6OqGpHHcZ2CXxEhc40BDZWz27rLIunSw/fSfaA70DcsiisMGUtw8
+1wT+ifpch5ck6hH52Zpufyq8GYkNvqoxk/Q3s1D56m2T8b1UCJMO4ZAmEQFWlunCl0gNVtcSSyS
8XuCKkSHfx8Dfu4p5hlX/FHSWWMM1ON+g25tpS8j3Ov0u2ijnBAMZ5G8qHduv3GFu4BWyN6z/ge5
Qr0pcXAnJ10w5MzQZPgX7OkmFGCcit32EKO2fN57ic1QdaTEhep1Udy5huWgURI3HSUM4KUlPhwx
Q7juar8IujGxjXYAoxBJEzExMrkm9YmbV2XgLIgWJYQ8DLyG4WwaXRAmSRRLuVkhFB6HLxswWCbt
9HuxDJzMN5xqLKFzwvrDw+GUU/QQjqYUsc++aEuPevrtXM5g7oqLHBlspfPeNOgiUritESpFGZpk
vZxU6xbqTi/S8U5PyHEUjUGhuEskh7+2Bnqv5WgRCB2LDvaimaITGt00AdQ6wkqTXozB6wt4G9vj
NpfoQ/GC5NI6fjsexbdmvl9Db4QMa5RD38glLvLtF4lq1btrddzTXTmADtrIpeU71ARm+guSQBCa
ztxehUJwdWSHACUoYL3M3Zo2AlCKdO9ymIzy95PLq8e+A/R4PF7Z4liDyjPqyCNUwAM6lQ+zv+Z4
wF8aqv/PDNjW5H0EODqBZTrVvsS6Z2snb8nXuRoUyLayFeHN9EF8Irq/81YiePWqtfPxL9dzIeh4
ZvCBlduGKdDZFCRLiAqWedMLr9wlmc1X7WIc1tuJtOSC2tmwLQTHLV3uoOtZLPH9O4ZIVHl1g2ip
/4EMraSAcTFRWfzd4ysKnQuYT33DKL7USc4aJxSh2fi36h6wRGun77daSJvJouTWNUMnF9oJ3uXq
DDkh3VmoKjcM8VYsJcdByEvMJvSPb0Y9ozuzZxzIguU0HWvPdv/+Y0Jg9wdKx0Wm0VB5A8LmR3W2
lIjoGA04O6EHgBN/mLFPMmUlgU3tlc24qi1YnqFsDMrdG4ORiT4adqECZYeiCNJsJwtcUVMrgScm
mMjX3+V8yoX9+rN14RmB0fXH7USpl5jSTsInZkSAPkc+rpi3nFHe6j8UeIPMA/Q652WpFCPUL/w5
FdFf+7BbGvTlgbPfPqqiODMizOB0SLLpd/euD1BsznqDXzgJddZmRs4U2HXMSvh21sA9wTALXmtO
sEO1qByueqwqb6/wu4tSWn6GioNBhP5hxow8EMQPzJsvbLDMCIPItibEHIIcxs1AWihfjK2IA32O
aePWConeUUFqNFzy84/31Qi0p1F6aEqMddDtUKn9T+wJb5v8WgbJzr1wsJKo8nsixki5vnXUQzp/
B+v0hoV0ZyHmrO8lQ1DecRvPWTQ1fCT/MN2ncIteHAIXqoB3sJlYDxFynjh4uGIPNSnXSkugytqd
hYfXe8jayIaxcFPsyBJmIki6eRGID1YTrESccUgmf+6KqLUQsAMWdzNYG12CUAkyxwTer0MtGDwX
GYcncD69cwNilI/jeRlppQ9xQbhYcMtUs4OHa5AnvXfUHrile++V0SYpbYkVIWDPSn7EVExMJMkg
kxvO1CwvuzLMRT8DheXj+aukF8DBDvmt3utrunrkumMbS62vLR7JfIn+FANXVUMkWEAHSKI3yNsI
d+BW2kIrk7CjchwrSuUvd7oriu4LeGK036bcJefXgcSs+sRa07CrmXjzJf9pGXu1EO2GPlGDNs++
fTMDnR7XDIcsdt1CAszLaL9uBQlaFqGZHjVXf+HJryQW3hTbUAd+hLEjQLXDbuT/+WrUdvBIrnOi
MXfjxv1IZc0qY6f0yhBeIOyjPB+vHPua853GqEKU22JFPbbDqtX7eBdQY9NPDf208uJG2f0V5hC9
fa8BHxfYTRK/bfXBxf/0yMpVztIecxDj2P45x1qDOQ1IMczHlaxZMIzM7YRN7WGX9YrYIocaEwPY
XOuH23HFSGv6QbzXVNrJVdfMvq5CAFagUGvyKzTf9dg8pZ1593T+i20OGO9wioHCwbeY5SkM4Pd/
7zbYRg2PxeJbwQC8KLsflJIm2/9W72XZZoJZlcACASSlSntEj4Adyww2o8jVLFJ1uE2x+95dO8r4
no8ReRV7gy/wO8GA/rJec3r8ZdpW61SmeQzaa0v1M9V/LVrW4IaCtXiUT0IWM8pIAE6RW5OWyzPY
3cm+7wh9i0p0aNYyjiS2Uc7+0soDKB84o2JroIo7u94cwWX5XWqTRpSYvYAk9bt2PB9x0s57VekL
ByYY+H2qqvOVj75Hm3Hhx6CvI5r5kSSF1OD+N8dCo7kw6ALO4y+ww/wWm4fb8Ytpl052HmFcEBDB
8XDGyJTmU5PdJpr2uRLG5Op0twWL4L7K6G96oRu/go7A8eP/pUqUdV1rRyK4VEk9P8/DzZGDr9LI
wkkpcmAnuMgXshq7WfGkXSQMzdbIvUhp9prg0wGipKj3UI/uOny8FGjPHfE4ayc8a9Dh0xttm2Un
VaSlAdE8qb06XN1eiwcsWlXPf9PL6ee5ycu4H3IFlIuI3YUqqZDvVckK8ZTh+ikHXlmjY7ajrBho
3EfFuWKIpyGTIzOdcag0PyEiJsYsXBXX6BTVeG+oYH0SU2N9rrXqDnNWZ9ODNHUVGDWN7OzEOz2y
3b6YppFXj9EkorcTDq3hmNuId1ZqTlpF1cExJzar5YLt+CJDVXeaSXemtue9ivR1iMvGHqFf3isV
RRGChOFoeNsp4/rPWsqGgTk7Ep7PBiLBFCjR70urIW+JJz5XTVcl5KzJLgAOIEOPUayggQm/CDJD
MgTOGFYXu4wppUvbHi/691f2reywNb4FnqPQtGqDu0PLmESVT9ePUrxjkLJa+CzcoCXALVx80h42
ERVi1vqKNbWu1yo8GwpkKtpJu1rMGEYZa1ORj4hdFY/UaOtIA8bV0Isv1tVUTEKHuZddD4qdil7p
f5aJdQu5d/A5wnIUc5EeHuNFKsZnO8SiCPw3KCp6ECee4wdFe1N1Gr38EaOtZ833NWDfs8E1Oqi3
kH2oYL/LAX+bYAugzBU0MkZVv/V+cB2vXsrMIo8fISd0xrcLL5GVxOigTmiyWOf2+UciXgU9RU1K
mEQmLs3onkjdYS/wI8W92ebGaMOgPhr3O/U+EMpKANPJWpC8nOPkdmNFZfX/NCbR1hQbvYUriTiH
4kbZhdTXueKvehTbqYx7yxuqj+RiOEFgqSGRRNl2Trkfrb+lmZGB3q5v644lmZp9JRVqN5vfl/TP
8+CJC3Lz0cN38ymsm27i1MMDI9ZnSOcRP4yLjPyL+/rEP9BHF/LSEV5c3UNNiRP6oK2xTTfnxq/P
RI73p+X3kPpXTLY7COl/8VoS4hCmMTVgHDRe0go4y16Bu4W1HG3pO+Yei7ywJEZ6KF1561ftho5n
8Ws2YQkUTn4zbleXLtUFWU9JVfi7bAcfGcCE3mVHYinUnDh4AIWF+hFQhMCtLm20TE7u7+WWDKlN
Ty5ztOQR6fNCFDeg1PjTY+84Q8VCtZmx7sCJ5T5eayA1DTYfBSJxIvNv9q9VhDK+L0/bxNFehTlv
dj65vc2CzahuxJ7Us6xfYSj8fJroOwZpev4SgNDZ8XlwIhChtxgCFgGl62+2WnWrbFnuNlXkqOtE
S8Kg/DhOJ6doDwxQQlC0X6QWRTQ2hr7meSL7iTwgeHu0LWKGo0rSFtTtL71+yyNDyyeIUe6gqei3
4cilkdGnGcnmfepfqtefxQCi3AmqM+WgaT0FJTa6wLA0QcI2pw13uED9xT2c6YVPSrQFaYmjIq9p
kRgWrHKHCtwZDf0gLcgNNfNxiAqz/GyGkOKt2NXrI87xSblMuuAKiXbuBKz0f3WXVvOMijFwcsDg
xvvfMpu+KG0etBm3oylNPxdl3Kc88od0VhBZN2hHxMEcVZ5y/FMmrfm0/6xZuyFtt9j7Bhzsg/4b
CcsCzj/qRANkJYQg2m6WjagoC/dowEVfN4eslp8Ykb+ywKHev0W2r8XT0A1ENcaQ/ImhI8amcydF
zZ5vXbeZnEXEUe73+EiSVfj4tVypqb0SjV4adKFOD1PSK0dHV1EBNQi01BbdzKeqa8ivWDjq9s6H
CiaS5JtVxo+Yrz/JRnOioskAf9hvHyWI36PqQykAaSmCWpfDwBedkODqU/zeOvrcS5VOBBEGZfcN
CJ6evLilEqgKjt/WaHhQJZmKqh1y+YP0GFNyPIxEjwfx4d5xPvIt3+S7pBzT0GoR/AsVfeDQEG1k
JXETVMW/BT2ykM3P40vEeRoyFHBXE/hexJNOESrkAhmIbQAEQ1QwgA4riGe8egHIL+ZrfG0VzSHN
E43+dOfKdttUyB3xGPFJolCkWCT7+ove+8P6OCkUkw1zvjOlAl0MttvKk/f3Ibr4oNfuXdPLc0sP
Vet8HZ+b5wXOPO7X6gYbqHCFTOTbYx4aFa/fpSxYjL7KzWV3M8n0XHywjcUiB+FhOUuWcYG3JUh7
w0RNMFafYksa0il6DhyCVarzulL+Vql3OizpE+VKeoE76UMclR0jOW0CBdlSlS81vdqgjQBp2O6p
Lq0CPzOTufW9UoEBx5FQmQFMKrm7BIHp242Dj5u6psJRlq5HlPTs8SKiA125t5750JDU1rcU3gSe
/FgQy8X5wfXQJSvbue8+rxIwWqhnfv/FAMeJfcWLXIWjwLYC8IJIIOx0hFLUrDocQJA037zLGSx1
jx04dnSTr/WOPoQNY1evBu/8R8mq8mkTiRqx/Wp/fU7Khe1inJJrqmeMJdp+MuE2HMhSAB3FTbKE
bicDi5Tn3mwfU/duCThzWtj03DI4eqOTV1vznCGCfLha/6fWmNlFc9H2HD/Sg0wIcDCg9qQZeOIx
vnQkhY3bN8fiUn+2o55ZPme/fl9gkgQvFCvU+jRWrrcTEMC6kLoj5EppVtcqvrN2KrLLTJ3laZy2
hO1K0zR1x3CnYdnjn22McHw6g0Qpwgrcjagx32uWTWpX6BuiZFpk0e7sSE33UJo0K6JLPcj4ikjz
V7OpKuL8oYoe0LD2i74vNEfN5t6K6wfKhzrct8kt4qe1ym+G0gpvuKMcFxpoOzMIvUwHVpw+hOhX
aKdA137leJhx5Sn5o9cNLhCQBfkbL4kD827+HlowtWCulBJHVLfJVcUtpeks0UfGbEqjlOymqP26
U7p9BL9urej1XR8/lSaKqnWQSd5fHy+1qjUJBgDR5KSeEEQd9i5P1YPU8n39/osFgacdWgM4Nbsd
UVn7K1BsiadFPBbsNXMA/hrT9Wu0ctMnx5w7BjQZ58096InAQ54e3/Gj8uEAi8Rqn54WSK05oblP
FnGP+Tq2z1Gs/9fg7Ps6VM5u061VPOtvBV4QM5jPRp0H9CzFdEoxYMAqHNPh+hZ/tVZNoCHe7BG4
ZsZq0YPADqi80Le3ZgvHJRG/iEav7Ywx/hNMmqr3rpcCHeyyUx/5Wy6ymD7EPlgdfFzvtvMbffX2
u2Uw9804oqu9PW3FJio05lp1a2tgl0nR48TjwDCZTf48uXD0glirEgTof8MQ1W5pl59zUXhNeoGZ
heWE78+L3EoWAeTYevt+L7Q8WEBu+drA+EkaMLljZCp92UZGvEy2/+S6tvjgAXgQvj3o6q3fQdlv
uHgtm32S9nLG6E4qwsEZTvGIOLZ8M5y6hgCx/ueSKmPLgKL7grVJTiniSV1UH+X/5UFPQE0kTVsB
wC/jfPzUAIinTjjP8dMPHBfaz2VuXVLPfQKLZvs+w1Sk2X/Wl6Xz+8d56D999588PQMVGtYoogpv
TZ5Efk/8Xe/11G36VMbELtAi6Q/NpvWip8FG6QzvEw3HK8oeR517liBU8Sczn5pxOGrH1690F8rv
MkeTMnxE9J1bmTVS13fsdC4eK/ZgupCSI+JL6pCUpOwNoMSHWgtczIaNAHVBiREIbhyqd+3q3IDP
yyVYQfGiWIlwi9zS/u3fSPQYDZXRy3PMJCovk+oqEYMGxW3TG7G/1DFdsLvptU6pa+F2cvhy/qk+
IvQ0URUwx791sDOt31DHoKNe5XuWTglvIpWPkK0A+bMtKn8KzLfXZe/6lT01EGHPYHMvE8vDpFz+
lWri6vKGtJ19y33JrzVvLpNaiq+GJ5nPYPILTbeQUa2ybSlL0VpiofjgmrooUJfZcN3Yw5yH/LvG
hGPjdIWxyXOqMSigq6V4LPJez5FpqymyytdLYaEkma12wZyS9lkq9KE/5hiIzVR5Tj8lMsfu/Rao
MZDIYzQ1y7l5CMelkjIvrTA3pCM3Aw2hy9L7FMU7p5CAwE+um+zDBKfhDo37aWHl4A8ON3hg/SMB
nSamLs8lQTInW4OCLpTZTJcQQJZQcr0TUXy90B+NHl+BUzDh7RfnsJzT2AULPvHXfj2wA1Wi5U1l
NEPUiDvv3QiJnk3HEHp3pGkvuxhhQyUbdbYyr3hJi7/Y5Z+CuQs3O5q3s5VdEJecKHV38cLGAs8+
QQlkTwH2eGONZF0+5tL1u79C01ZzlXwAbKsDm00R+syjmTdLV7ekbPa5yCiv1j+LnGYgvIOsA3hp
nfmZYUwv9Cw8ibQusVD3a29Hxp2BkdQ/KfGU6Bq3ylAViAGUM8tH9sPpnaHgiYOW7E7tasKqzynI
lEg0a4ealZIePAkcFmYlhRi+NYT8K/mFKbJA59GzdJEgV+knAqyqny59vVur8k749RNCcJVhu9R9
/2l3ky8Akl2cZfltphfHz3yzZRsrtXhLny9YDectpxZKnYgsmV9y37EzoqQVgH8/U0DTs4JJMv2b
G+tZcUK253c31DBq7vbwY5D0CVSWCfdd6zGUg2kZQfjATUwIoxRlraBNBMRNWD+ifq3Jp8ZF5C9z
WTKuKxY3JUMpC7+n+czv55SWfbg34bxZZtxFG4GA25ubRWn8jpUYSr3kHrOC6OHbEYLcpiSzzncT
RTZY6qfC4aRQZQ2jVublD4y+ibmwirKNeQ9vdbM3f4ekl7kjjw6IHoUpGA/ZpjSUrNFuOo0HhkXx
T67zUK2Mw5GU6W4bgjkJbCocnfC9BubrCbqDjcXzaYPSebls3xueVcjJrPWrQQuZB1Cgn0lD3eHK
gT/6/vE2y+v3PzJArxkCR6VqHgX+vw6q6WxenIoS6TaOws4zLxw6Ubh0DVKfNb7b4zfg7fnkAzC5
f3Uu/HdBz+FogCqY0hMAoLblY5ho3zG8RnxasZHFcqt1F1hztyuXsfjR58os7qsmkkwd9CKlfGJg
8cQ7c2PQ16XMVEOn6utgrWoBKOmk6oQD0VtZrKR5UzmgBucCzB/W8QMsirkz2c2TH86EfSpQp03K
g5KsGuT5StM9GDn1CnXquoLC3EW7jiXDAkb7x2vjCqwmE7QEX6ul1PaGZWhm6s8XMwrR5OFmzRvE
u5t/zRkPtiNVJiv7angxNYqzAue+pczkobbZvYIDjoQsVCxqpQi6LQWy5bvFpMchjJREN2JMxLd3
Xamk0ibnaGHdp9EVbcPDF7pcpTI3MUoHlpDlsYcbEgQVnaEsWLfMZshXB+v4uYbte/imHabrXejP
qH+Duu8eZE1V6u53EY3HQHSpdnc893H09xHVoDC2Q5jJXjRTWQfs7QmsqTl58oGKnTitd0eRfP1G
A+dDO55njjFboqpzQRypHu1nNW3Ft1hA6Ju8cSapnd+YTV1kzYW9qiWAWDBVmvteeB+1TBotsggW
8mC/Gnaj2Dm+TEj3S2w9monbmWUp0eAXXk815XXZAp694awBskl9iG6umW5Q1SNoTyooKFWYnaOE
+XlnwffxAiUu9kqzg///HiyEjO7/ROFeryNLHyxj9i8GXqWr1z739rrgzKzJS87Gg8x0MOnf3H7S
JLNanjRRkiHevVSVLoFWd0m+84Th42TqyAgGunaRQDDEQRjGIc/m3rKVmsZssFva18NCjWivNkdf
zFsfpI/BjfK+7ucOfxfCbXJ6qxylYrf/kwNRrpHMH/7H6sN9Jh82xKiQCKZDuWzYpJDNrF34mxPJ
TzbVKfH4XWHcDk/SQLHqgdU05DqsToiPrX53qSSkblCwu/FoAEfZCPMaVrNaDd5rxYm7OcJwGIQ8
1owyuRYdJaSH4l5aVxg9c/NsNHaVG45S4zqtY/TKQAlJUe+IF3U3+FmcBuZ8u5hgnXt8pi1T6CLt
LE2Jh7CHWrouHMiNqU+SJsHKDafMd0cdMFfTQExjwNb+rpSUp+tclSYhaJ8IlBxnp0EYB/aTveOx
EOAXKYVbdZCsiPgKd8qDsaNNuzYCSKOdD6ZOKsO6AZZn8h4YgJSAtOj2VB6t7Oi63iDsJQc3Crvl
4y3ZxS+S0N9FCmecilj6fEGImfwyJZLDYSIHXh+bHlukb0tYrPvBXoa3a+bn+STYeFSZ2BukP/2c
1Nj3HzKPH9e6Drz61xi0cmCMiK0w58R/VurEqGTpeyrGoqAxm039JBVal8/2WeDY4OqKtZx1ITHS
8j+RYuzh0rV3ZsW3XCC4hU5LZREuTHqAlYsCYWPb3001Ch7UucXdLs2VK2Lzcan1F4Lw1BsScDJt
RcS893DK0Pw+HZKzPoN48yJgc//Eko+kvXNitqhQ+E5viVQ0Li4VPghrQo341GreEBEycWQhZc+8
8Vt5WuJORtVyOthBUPHePDg97hYAMzCc/hPSePDKejvTWh+N2tmPjt6sGPtl8sODDVMmdl/soqL3
1RbuGQL+3Fgjwks6r80LJuBH6xDiOT1zxBxxKX0/PxegX7B2Llwuy2xoVaZCHm2G+bPivX4xWFyj
NQ+oD/mJAUbIz8yPQDz1fYyQ55/UwksUvwh5mwNrn2VUGmDMpp9owvcA+FIrWbkApUu1NQH3OpOZ
NjJ6R/4VP6Hr1Cee3yJNclGCbigMyRgKSjpRNYtoYECEFGrEuIyCWsiupbn0qgpKFoxZzmS0T7DJ
PGK+ap+oZUlMYqL5hSb6CMz2Yke/+jZOYiJvaW6lCIq3HpxuZSGJPrMJy2OkX7hmqqUjUm8NWlqs
2xDAfCdOWkQ36BZP5xd78/u0ZvOEij/EMQexdAOXdxKXpaJNNZ79TMQb3HHhqjxP+XfnUGSjIjZ8
7BDX6GUuT2khsfdPMKbRrdc3Ueee4Er1ggKpmasT4FdntlLoS6oWJzYHTpsfuU61yOGr3dfHn+Y2
SlQzMsaZ7UYmDjz6jTYl29bHbXuvYLsteCVKLNC/yi0aLzmT+3Rjv5SDnBmW3nJ/zqXCf3XwE9kf
JSnc8PErcE6NQe4C7ok31ZhWdvzJXcsegD2r1ZnTKZLtTVSXwrQ43E9QBUMWfqbzbDMeASasbEtX
9iUtD5lJYIsqlkfFWvHhMnxHPszDj/t2U0XlsgeUxqA1pO4bek4msDfiPyXmr1JXkm6LkpXh6HLy
aMh4xbRvVKX7wlQgYeJ/C0zW1BNIZXZR4/qz034DxhmIfi86d/I7m8ZEznhHnNllcc0qmviAz7fq
PZCM0mO1EJEKhGntl0aM9U1DJbQlZVyoHQyw1Ajj3rdBZ3j+DCnotnpOjRnJ4Z1taQ17VGlWElHj
SWETOFNZd68DaIhy3ijTvkO9dZfVShDdMuIrgBjkEe1bhPHA9vWmMuhJDBnppSm6iCTLuFYYKmJS
SPai2ND8tqZ4QxRMO14EiVSZ+Y4dMnYTlwH/lzWkoJAnBsEjL1+Csf246/KX9x6E0+p/H3KUaona
CvIkbSxxcVqm0ggnRvLbEPwBs/uiC+mbntoAc2VpYU6nJEKJgWeqxNBv3goeTenMIR22ySRLYCuV
tQa96B47x/AFhp7spGWO87uPNTQTwbkMovC059NHl0oM6rx0ThlPdkAJBt5T/FwdmFhq26p9CAW8
faGhgq7kmfq9On1KQVTvALIbJDkxC+lwIimzPBIW4Q4RFuYQFGsuSb8XW5jYXvI+DshMyjtbwJzP
enXVl8spnL22AgeQ0VREKnD6w5jBOscF5Uj4c+WvRL6rQclTZNr1Ggjiotp/g2wfvpFNUgGaEI+3
5beWXY6gzJXJPhAZ0+uEECxode3gIMaz1AFjNBOtTaRgqH1nOc7bPKYcZFYusnZOVlk2k1eGGcpi
ebdHVhXcraT57NtoEUYxoTucEZbvPrqQYZODLnVGyhoNZ1JFUgfhdyEhY5gYYC6ksWiVgWMrOb7z
u04o7HTVLHESp9nxYIdVc5yrsQ3u/txaqqGRXdJxcoKnP+Eu5HoEijVzK8wk8p2BhhbjUt3xl9Vt
tsWxLZ37DW56oKoWijLpIAFq3LrSQ1m6sH9Y/IcQBK8k9RHtrcS/yTjo+FAxrJ2QEanuewrs45+9
MfgSzCl5PGF4YF7f/B/ZZ+2kANkvN0OsgjP+Y8CnbcDU7zXCAUk8vVDUOwty5bki44sCO92M1jem
1aUTtNXU/RCd6g1QN6HshGmGEt/1gEKXCa68HEgD3Nk/AXP+nqE88kvICzxSAia4Um5vIJmfP5VJ
KAs9ma75ognAc2kfrBnnjmHiV6aXpeQzNePQhskeb7WFf1LzP/QwC3yeVrnB0lyYfWr17grRqzSg
uOtL+JzPQNa/HSkYrUqWs8yXrBRlviKlKqVc4Nl2XADrC8yuLAQTaWtBUjwE4BV5OcjIpB47TLIX
SDAemQTvu7yTsWg4stX3dGiLwHGPYmBVX1m9sGZ5ju/2dRx+lwMZ2B+7eQ7Yvyt36JJwuVgLXc/c
+Au3RgfB6UNx2s81nCma7stJsk9q+gLO7QscBchh8qRMHjVcKmnC0xKHKLAi4ijQR11PscXC3CG1
KQbKY4tyZwSNysBIcvCVl0wDpQGveUQG5BdxN9/rqZ2L9X6RAGPJntFZPwbG1VVOPX13uh2lYAvG
xff6pLCJNNZyK57H2EFOwx2EXwKozNXui3qDMkV/tKv2OYMyYV9e4alOsQx1wKhRUjYnks9ox+gL
UA2jTRKawE3t2F6XL6+39QGrvk4lemqG6m3+iya41ORMa2CR1sBuszGjV/UoV9e1PbXim7YGLrcn
KzsakAh7AMTDPML5TBa9OPj4KL/fLdyvK9OOosOuM+cpGj2SCfanA0Scb6J+/tFNQff50nR5qiPs
i3yKuKMZe+W5qaUCh8hom2l+RsxVi6ggJc2SWDL2FOoN5ka8LDoAejSfCnygqx6v7BhqTtg+YhJ3
XT1XmrwMGcjglb+m17PQglin1y5LD6g0uzGqjDXVMTb/l8g0dMlD9RcYCHyH5fP8xkoJkN9lnVO0
z9QE7srgThk0ud/YCV6SoZdPqmy70W3bacWS99Bgea2/yYOvHAqYJ1saUqg3K381evFbz6fT0LrE
fwALzPzau1zpWjF/x9NurajkBtz6ZyspufTklWRSGJf37hYM5+PJDU9xj/lKK4MF+8fe1W4P+r9a
sr2hwXrXjCgwRAn+aj6p9r5Oz81/CgL3TFk3m4MPe2QuNMtUGxJt8mZsruyMaXVc++RrbNXdgogs
SftZiHRjMxlleiQlXJMj8lYA7CTWeH+VHmBpEh6yvEx3K5L+7aEEJD7rRm+VcxnFS09cfAaKinWZ
SaN93I46PwnBn5tlHKeNea4Hi/WyTqtSmTIlqDhTHAZfVTlwjTxlvvHmtB+H6EksvqmSXeTImReb
M/avVnTj6JzfTCpGmf8sWrAevKCqLO1B4U0kbDPQ2A/BG3CA/wkW/MMAk+5RI5ZAYiXphMCqrtN6
i712BYY4cFbhw5w0wOP5Q2GdYvUmuWjIe3bU1UMD0bQyNVfH0ofQ+dXKS1tdyNkSp9ptMfXlGSqO
5hFe1rsaXedzpwHceSzIapYZwB1f0ri+X4FBSxPcYS/JVgO/YHdOWNY4EOz196J7i/E1hOlbMvBU
qB1IYXkQrDYzwKeCig/5enuNlHp9pyxcha4cmSlKUTdFJIh1hOilEvNKdqW0l8bal8fq83hU+wJJ
Hg+op9dL5sbdzMHN6FZGne0+nKmiQIIissBrVd2uXzVUrhEDqisyAew8/FH/k41urz7sQVEKOAbn
E8Ft3dYAn1Rgrr3VprxJ+rgzIhPJNOCLt5rTj7OcporvDrtDaj55di4r8XYGpgp6cLc4MpekW9+s
I+5HmUR0S5mZQ+WCtlhi4Em0B3t8YuDqlxjyNCgaKFZe+2DL1s/trwdiM6CJm3s3e8uz+nNrUiFZ
xfz9nBoRxDLokhefZ46i+E0WzZGDuIl/SRUpkUxyFfZqzMH7OO9uIVXpZelCAz5pJMrD1xavmB0R
QADCcM1jtS9EAilE4DC/d76CDHB+9CfOsdWo59z+yejQ36tXRhlwfapGcXSEbmsrWVvHR6uXS5c1
9G68mrrPjhimsbo9YPmAXAaCBi7CaCa9KQ6rE87MPMe4afyKSJqUMKlHgQle/39AZnVET8jWUO9Q
09cdOMDJ2+d34MsLeH6rV0m5pMA+A0iNb3pX+m3e+sgVUXURxXvrgF85EsLqvbtqeM5uaGJiliMz
bZLhv6LSx5uJ2GFbvY7B9kfFyFb9NhEuEyiZmWCLp5BHGNOBWujEfzfvh5HAMhDRUyG4Uo+dbKKF
gjV1Php8cZck2snZiEWIsyXx04rwuaP5zERw/ymN2hQRFZkp+BC6vEfM65TDcfvxIjgrduE6Bra8
0M+WaC+4NDrJFjzNcudta/hcTn9j0aJr17iAPyFqjHtwoRY3pJemnrvLiWeNOd9AxEG+n7t8o2Jm
v1cXbBSM3gFchKWRPV1mKZbeF3GqhjfttvDGyvIYTNWxZoNb/inq1Z2/o1pdnr49pTJVLbYHRu4r
2nKs6GptPcHcNJYZ551E5MbsMHhle3VPdBqsGYp81i75gE8/serq0K0Fg0WpQ70Ifpi7efrBw7zI
49wsLtfBCWyvfN4cieZqutfrpoyD7mbMV6Idlgy9H42k9f8An+0lKFyRa6d7JS994rwZ2MS1nx4p
S+2O7kkyAvJEc3UsR/XpuSt1FRoSOImK/AMGkirlBTk4HJlry0hr2kwQbCcUNMVpdGfXIsjT7BJ0
qQviiKBgjXjIB9je/WqZsQ7NEQEu9TMULjAhRIY4JFwXMMccLXoZ4e+vTfdh+GeOmu0cN3hWccCj
5PkILR6F2QJI/jw/Se+lDULI/OB3+ogT81BicqSAogm9ESftT7apNbFegrtARSrQylyc5Do3VZAC
eQNQZyad0sZVqMa4NZI+Gzbg0ZQ8WV2zREjMPtaViGy+l1JghDQUQaLAP21WTG6hZM2TRhED/aE8
ASWxxxwia9lJsj9MW4F+uSqo1TT9vgAndRju6sGC5zvb4vI4IR4MtzBwEB3MhvLm589pAN/0kImk
hq3V3NP7vPD32KPhe1tbXg47+uaYqXX+P93/iiG2XNr2qdq9qxYyhqNyzEg5k779Ui86GZSuKhFO
q40i7JSjeH2qLZlMvlcpOR3dZWmo0IE7c+iNgVRJ86MznlgRO3VHBKT7Lg/dUxfnw46SVP1IgfiM
QXRSMNgHgW854xvfAl9IGTcBCpl5rpVzKgtGWhJAT2yxyFfiKgFmLTK8aSVf2Y5iMVh7NCA5O/XE
FtG0W+LkYPioQIRI1vTjtUWu05fDpueQkj3FGB07mmFM2uDQCLeBqtRZ5rs7Ye3sOOZOaNztoKzj
xjmXfRyRrO/SJl6mIrESRG9v2Fp9g3ShUVeldSPKhtef2hrNcvQsCaKZMx6woUh9FYHuBG8URgqf
o0wfWk2IgbjL5p4FpgqshqdY7c/ZDgsXmKO4KWcjN/Z9vzYJRTjQNDnh4RSI1j9cpUBOCVjVRp6H
hEfppvZeLcNf/AUp/PRZtMewtZPQHrHE0R3u4BCYYElmx5UCZi2wD3STRnytO0T+vevr7cFAQUyu
8fPDkndzRbzGLTTnpkjRQQszdg2dcqyJ7lQdtPVeMKQzlnt9bAyu1C3EjpBeNiymEmb8S3YnHR7t
vWhaNjUNwge9fNIOndHAy3HiHRXwyYRotfHOb5gRyMH9oHA316V/0t9H2vW4lgFZHuAbm1/Cd25A
md9IsRuFakZncjlbHqPsbBPlnuPVmKAWJ8Aed0yRPxpa7BZ1sonFxmBeNL0kDn2f2Qfx74IB9YqS
tv3KIRoZ09lKj/yFNaw+ULovyffTuLtGHakA9UEFYX68OF+z6quS3Om6AU8al1zg5MJ5j0Rxh8oV
Wyfs+HrJqN6RzDuvQl5GIgByOW+x04JqZwmPrp1GHVW56xgIH0xrYf5DBD7l9epmg9AGVt+0xcVZ
CfoLXxIB3zY6oVnloSCqTq2+7Fpi4a6mpK+0BUxujSbeJW0n0aQ9R8l/KhrBGO3ZhzJUA9mlEceK
zmIFtidre7Iv643tDgEV1nmuFbZAcfNOZcZ9T1l6jlMgUPDXoz7EJAqks/R1zRwOIlIPxXzkUPhu
lI94ruvk/f7ved4+Hz3bcU3nOL+e1jNfr0tdYLtOIFpFX2Ms4zl0zBQnvgVnMWJ1MXgAgI72m7Br
Xz/DssHlhPstdBxYE47iIWDLh60dCsCzCyQGd72V+JSWhBjGuGCfb93gTDH0c9EVtFPff6ZFYEfb
YLzA0rDIyfF68wah5+a0qqm41NxX0y9til4DJ7su/BCsPC+er9KBDmICwEyFnam0a50uchoMi0Yk
jkrljGXIf3ay4SaUph9Nlw2GhB9v+5HJjxFVAV5BtbtpxtmxYzT6NQlehuie9OX5MUrV2WRyFxfE
/3rw6VU/JeOQ/8j+eQJ0DmXOinW2FUZSs3GKdvzzEeHaKcGXQZQWCyxflez4bk++GbqvqmYvWb+I
J5QSlRm6PJB8nKQsrT9zOaLLJmMTT4l6gM4GBKFyGKuTbJ4hUX49PYsh6fZjWBGnm54/yEyI0CQe
14edjdvN9AhmAr3TJx+Si8GJxemTmmz1tFeBE3zo8yt0mVUGx/GEa81rGSqXUQV8rs7QNS9BrJwa
CwtJ7dWyxLbkx6Hcepz8ZULKi0pGMTgUoMWAtF7qk66kOp7v0USDqd8cE5E6/atPfhnN/0cNLjTE
xna94XdmbfMwlKsqseXbeRECtSgmUKdfyHiij8NJ1AkjqDCzYpXDH8NTViXgYUbc1nqZr4Sy04in
z/ju+DC7haWdO4jHVZhmzLIUXjvHxBJRbvpNVeqB3/TAuL1hb+8NLwRbo/k/vW4pwUj/TgCkcE17
yWZ9NNh9riXPi/mweSvkjUoezI1qE7nDnPeeDQOAPbH+YmZS9tQNIZFP7iIcszxz8KQmEqTzZ0o2
w3pqd3hXg01TSLNOcdtAK8/SADhTuIPy4AfWI2T7Cy4X3NEOGXLs6EmyvAkOFRzWIJcbaWuTVtKA
J7zAEUwBrsMfuxUBctMhsX3/acgSo0cumrEScB3WFAEmtvDZKgv/mYsth4+RvbwlC1s8nE+KjDXh
vp1ujW0dz9jUkCzgVA20GHcJg1knse07nqCJDb1DEK4klbt0zboZfbgnzZ96XSFXVpW1iDsoP+PX
Sqy5xuRvzauR/ZNEqUTM8CKSiaTkoIv7WjbBHhyqYQEKzqRGsLby++aLNrndGaA7Gw2lhRqVF4tz
Cpa5qacV0ryQ++3zS9fXBwB1txm30FbYJ/qFXOwW/hIt6tQA0AwryevSNiFsQ621qEU83fGZoFiJ
bcJZ/GjtgayaXiew5rYb0oRAgnlcmHEXj72kukBwuwfjZwuRRmJHnr/2r8+baGez2dkEEgXuUzfd
4Lssmxjd/cpTB4L4pSLJaA+2qJAFsfQLrNwMSf35W1IM84muN/+nP6eeLmA5/fwg4BMEJNfSwJeL
f7gNN0ozeA7DtC3PuLjVi5hd5wald6KMmq8r0GzsPneyIjbV/ZobGI94MQ2VWmby107e1lg0HqyE
KffPak43+aoqAqvpiSGlMbpKi7k5ICSd87sK3YM2xXJo8vZn/MiY0MQuzH1ySI3u5Nv1krSCpbN0
twcCdgO4wf5qTGUYsMK13awMAwuxKp/TyHyNi7aTEDEyvaXGzVT3Z1+0Rak/fPIm5tvkwklX73Pw
XTZXNzWX2mpaY7DNv/HS7XRANFMS4hR3sZWdxmn9NJsTv7rgsfXD+0iEhi8g1j/2sqeENQmD0HbL
5aGMeONYL6Sz+l/AguWi0Lrv23bS9T/kpr8EwK+v8rshWanrwYyNiYsK8ypM1mcrK7AJto8nGubp
p9OXYopMuPcDMWhbhYZw+gYefQ0ruO6Ev9xjhu17KKgGwn6Ylo6bT3W4209OG2vuS8fnWsg62f/b
gIjNEyPjs9Flv3VSt+E6ByfNQr2Pmx0aM8Uo26Mn3xSBn1yRSZgxN/r+JN1+XmrY1tNwyOm+wPEk
YElfEdPh50oFa035dSY1yOquecFCz1WOKCScD3fU63o725wrYgjLcEFP3fC/eLb5WGOcB2QZa0ml
JmW/ceahL5dgu/cPvo23AR5caMARhUpZ8yxLFp5TsdmJUWklWLchNtlAFvHISZUjRpt8BCdLlmSB
SFaGzgomlzzNdZIUrVqQNWz4hfIRc49rMy+9Odbfl0BRx/5wdbSMB80KX0y5qDKFuNCeZMkZwoIg
opMJ/zHLavBWuLMVO7GSbB1kBozz04ummpbTzL8KUgcYpj0hh3dGNB5FGARhxGJ8IO8bkgVVNCkg
Kl5jwdkIVgzd7Yh0NyX/EZANCDen0IADG7eeiqj5HagFBKnTSbqvPaVQb7Nd+btvgAUjRFNjYkBK
LY2LhsCV+qMW+PE+gSJG6jBv2Af9yixtIKOWfQmx9efBSthwj1DGxQoHWCZLOvvqdANldIqkYBDW
RQBo6RZXP9a058rKWnUSnmnLr8/yoS10iVg1imkaAnaPB8Db7SPqS4voDTnTtSe+2mP/dyjbYc1B
vq0ao5CnKCrzOq5pV9IjFQHjbRS3tLSp6bVyhbfBDxGQM1BQvMYJuGFsLFIsPv49HGL3E7POuZST
YV5l7LH7vXXG6N2p3d9EPK0S6NU685I0SKmHBt00vtq0tNZ1qtnm6WmRoOnMPjI6hL9gCMurgvQw
UAQJN+s0Ww4LI0arV6PmHBoa/GjktnjKdWIz10ASdAiLaTlVFapYCPTu/6dYKUoyRZHB+4xgQKhO
qlHIPMx+bSrYlyh1LaAaHe+x32C1g7SlQ1AFHy+0tfr1EpW623daGEO9zDUxcs1mcjVLhgBYh3Ao
QLNzV0Pje3JpLbzKFR0bTU7KkYXmmNFLzMWug10GD+cOYqRgtoUIRfvQYGyMsHwLdmKb4l4X6DIJ
PNCHfYqBM0Gcr+F/URvAXkNcMaIDEaEO/r1pJJpwBKZh4iVl46qYDexHzhQNuo3RS1lSwy/uYP9M
5mym353UBVG6tDHgzYv383s9xLBvSQbnQa0q7O5CDwiRJznSPgH5E2cao528D68OnZTuOOmQdPI0
1zkC5egyXwd7jy0RmDfihppEWsOEsxtSmNqAQZU/EEo9gyqCjJFr9EZgqJTY2silHDUhr7qvqBF6
N0Fgb/ToNFyu0NmKqlZesHIeUEDLWN18eqYYCRUO9OXUzEGFyJ65CyXiVZ1yE22XFjyRnINVZwY3
eqXK0kjO/PyemzZI6F8ATu7SZf+4/3Hc8LtOiXxBt4t82HPTeTXY2OyZh8RKSNTyv4AuINBanHr8
bvtN/gM7MzxhEIhFCsDEfe3fdDTW8WFT/9o637HOUmB69FkIK7MLmxSZX0z51Vwv/tw2g7zmoYsc
H7qbCW4KnqoiZRakxDi3WIe7m6p3JHD9gqGYxjq10+4WPSwpfHMvOatC1PLy2KVorlpC4ZoE3qKt
fG+lNfeM2lJ3xXYKUQgmkTxs6zc8iOOZienm5xkbXB8J9Kk+uVf5k6oZMEkG0hdf+yQkspAeVaiS
BCflWpxlq+h/WukFZ3GdJRjn8WRR5JcGP01mvNVhURbmb/ETPapHL97jTYUsTpihyp1apVahl2EU
0RwU2VxpvJ3++OOD2WNdASb1N6YEwP4sbSVXVV1jLz5AFCT30qT7j+bzlhUanDsDJYUJo6JcCzqL
z98IyUw7KW0OhL5eNoBhOLiZEVhL5rKZGA8s9aAF2ajtiWHAnsEjvP4CvNaqC2LNfACsgu0a3bzS
vTgN+CGyevOoJipwKxhb7rFtwcOV4HwzkA4ehwqrqj2WRHhzGz9+URvc0s4soAxmZr0iFEjEsR2q
z8KeSAlyECmD1c0bt/eN3XBss26VR9AFVBO3BiQyJO5zsX7+pn0MnX+tc0s4HQ7R3bEwfhpUAKSC
EW+0vvk6aBEFpQCrjKIIpXdy6jxTRXVH0T6ODjRh649KOXps04uoJHj2bfzndMld9iNlkqBUUaii
BWe4vXfKA6RVqYUd8+la5s786JUJFR1eNL/Z9jmhVsJdLcbynYXNSaQd/FrRzWZ7Uz1o3kVt25HN
dOFAp9Oyeoev21kuLI1sl5PoYHyR77384KSDmMCbroeKeQzMvcR493msfaPPlMCywXOP4n08y8Jf
ilRj/4WClRUT9JDiAF3Rh/a8pnauPJ2EDJTDoxCitTyRjeuu35rK4ll52iyUxdUVFZGOs8920suq
QYs9Aj09/yYZdjxTWzIlylL6qeM8Rm29rv+LSbx7FDizT9oUoBwBAMznWqgS9Ba1tLIvrTO0MhEl
nCwwJmYLrJZvrXQgNIWf7hNMgRn+b1OIbh/UmR5IJfViNeJS+fdBu5lqIpjk5t9D+DUR6TV+F+fB
7+V+qSoJg/lRhKS0edM2zO/zLHR6XJemrE0D4OK4NFosXebJ4Bb7t5W+jsF2A6kFxFCxru0kdwbH
LNKk3DMQ2ATH0e9Mpi6jkpsXb8e7pz9rDk+I6/7hrPtgMu4+byTSjfxKVCNhzjFITzpgNZqK31Xy
9x6YPIkjxu3w0ttrKqgGitgmbkFA1xpCHyz3l10Sl3g4pWxfZDv67652doFQSpjZzyjlbNb7+PIM
RPYFrSbojNbYX3TUlHniPse78s+RTBJ2JaKb8UQKu7SFtDjAMYe9kz/SqDEyAO/rK0P8RRkP+Ben
KnhXZj/waE05zdoCXL8wYGcVJw73R3z9CoSkAzEOT1GM+tlRE9rze4QIZwMlbGPeKrDgDlQAxOsj
f9BBOiA0VlXPGbGI4c6gEXOrlICMdODUXZLpaXS4jEUvdkBWvD9UwlgY0UUhRjuommSyT6Ys3JlY
XAnCtImpITtYd4QvtF2iOTyQ3cIWJn4DIeFksWGDtcicH8vdqpOpkbdCRvQuwLYP3CNakq8zUBpf
WsEGAY8hFQNCmR0Y15yUZ1Py1ThacOPzZzKHlUKK3mctMP4oWTleHdf2IWNlE07frWgbHTgTZKxO
fMrnyFwcIU/zeuNNP31kvSsGCCK3AGdUr0P/N4z9iu9TBTzI1q2PXIH7pM9HtFHtClYjk+vYbC81
3xwcv51wxTh2Ukke2fOiF5xbtQ+Y+Tv8UcquJDw9gkpJ+yk17AvOIY8uM2kqps4yj3s1tnPFS7RM
aJqGO39USi4YPP4DgDpd0YYeVat8dqTZ9cclnBkPHPW708HfaM2awB08UqZZgNLPPqmC0/YRvXeN
R0kMaMq/0kErklakuRTC75LHhGpc1MxqfmpZr9KhJzhqOO8mPdVYTaJ4p7Qj54Z7/wiHmVDl9OBI
hVCvvWh4RAcy9Y0ofjL+QUms+FonniuoSr1O9CEb14G99hpo0feE8Y3oX5b1Z8dmE3TcBbqhT9E/
W0uC1Yr2JNZ4aYYArxlXpJeq/dvIY7sCvo+HOWWtzZiJcsdyDn8Cp8CSA1iW1jatvp4OFTwG31xV
1RvPABTXmQQ/MwWwDGFsb9oyr31eLJsmhRHmU3PdvpMMqQCL22eR4eyq3930MHa64jWKcllZRS38
i/M93Y/aqzu+JU72TGOyjVkP0Yrj/qICgoJAkqs6xWkQJrlT4SB0AKexzBzTZAdjoyD86opK++pI
eAr+6WH10gmuN/clIbVb2D0ZrqtNACMHwyxJMq0t1CO4JrfJG5qqmCiR+ZNuca2T4MZtXVrBIQW4
j+rpV6Ws4ZF8tpiDVG9npWOqVDSpBrGRZUm05LnFGivqtuFMPbgoOhXJvqOqM/ifLzHtI3/Jrl3L
FG/rsD/twpUNbZZilO5gZdMPwjFTWac4E3rVVxZw1xLVqvZpiWJZYMsDfnoD8yCB+2+yHEdQ+b3J
wSX6VLkNHUmI49dKC9bWJwCfAwzgS3ANsnWwIN284TO/sq6PkFZ2i+XpKMsbuywlAC+bGv5zgg/k
WxksONNT9sewrCLAzv7kxgbaBhPfKbicP9g9E77f3g8vrov9b4yZQAwyry7ISFPuVGnMMUFaktu7
e5izHKZP8PauqXZPQIZn2IGPlWYyZVhtQgk2PIw0szYe/2YkWStUFSWduwAeKUON23YStsas/SWX
zJ1g8IK/bJe8yCkBIkma7mA00o6Vvo9MY5B4K0JHJDsKBwF5k92E6unX2aPlU0bMnbvYZVHcdcur
aM2AZTz8SxL2gtnhXFs6J3uzcpFF8NmPIJYLUp0CVq79KyPKYWTr+sh0E3EAxLZi5XLpAZ641eVz
DthoE1vEZDunbZbltAVe4iZj5L0fUGLrTwAnVbDgXTtdRTbmCsjqyC+6OL8kdJld0PoaDzUOdP/9
791H3LC4DZsllhb9PAxqEE8dTPy5K9R7MVT+5JiMxFUCiEsXDDLIQcnSjI7SXwdqLulEp0cbLdTm
cF6HK2zA5infD1vuoWsmvNO0vDr+mt+rBhOcHZYr+5RYzzlopO7/a+26DA/ve7pHEMqXYFzgIfZz
m3Zt9Omt6Enswki1lHoTlpHCJzR3e/Fk/G7iq3lqOr7s6QKw85zSc2RNKA9DWYLKAJ3YWgMIn56K
TOGUZFXp7HSb+sfJbdFOiJV/rLdRHzVLno/OLJGE2Mb59ur37y79A4rIKtpX76Vsvhdx56H85od/
wiIk0N8Pw2z/6MYtoU0A61s50wR4+wVIXo++V1v2GJLW0+H193pWLB2h69jiv+U9gz92e2ND85Ek
fn7z1mJVqbY1jqx9e2g9dOuGjuZeKVb/m7uVC9UEQ9sQZwfIiJwOQxKGdMv9rtiQh02rNipcgbjn
NSfAvIr4Pd/x16Hp6Wc2lJR6+3sBY4BVmHYqv+Ak+tdiWHplPxBpmse4ipd4nqoFfhP/rz2Otpcu
zRFjH2qQDwDt56GQ4RGIQXw7l5ygBYE9nHqaKvGKjoQwQ8VsndiwIU+eGu+wqJr6OWGftO3kL4MR
lMtmKIaUthj5YCEG8ZQFmlrfjas5UGGXhze+OtQnf/Z87B/+jE/P9Z98JXeNIcqyG0s/xYvQpNeS
KQdtAaEUcOVSYk9X+i2L5qjV5SG0P3heebZAutzYcV9BS4xwn9O9zo9Fja6bTyhKrxHu0DCM8vvx
pLvqiWZ9czeNKyw9WluFVMU92bsXS4N+ifNH9N9wf5uphTrO5G/5Gr4eSDq7Cy/iKAOf0RODagal
KAfy1lIa3RFfabgUpjGHAc3yDSRCS6jnix5YmTjTflbojPQZWdI+I0hLCAoJwtd8xbm1BeK1oEGM
Y+nJUzG+FhWFR4pKeSOAINvwYvSGkyk7DBk+oqn2OrdG8qOWJlSgivvUqHTkTwQrUrC5wScDYcdQ
OIXIcKLomjZrD2PoUSJPWnx0cDMIf3E18aamHt7QrlkcBqZcXkhdXGLxM+WJhMvGMJdCJRnO+O92
FC+zuhswNCwEED7XiifSEyQTjKNxJuAI+0ScDauZbKMQhTFwzN1rW5dE3xmUTZEBDi5+5hhj16z9
9iNvpOyMXkxLwB/BzgumUiOcsj31YyhfB0+gMqUUGdwLUpLD+88awlqZKk2p3vZ47TLH3wyhsCoL
tqZUW5sBhHj6uApiFCY5/MFN4Ih0rcV3PSIsx8D4gPEhOkFOzJem7FoWRfIOrmV4BmvOwDO7gc4b
opWkV0J2CWe3VHJneYgqsavpcOWHD5NTSzdtmkTFMSkzeplBlto+dP/liXMjSXReTEphlgMFvtDS
/VMP8fSqlkNngDtOEsCINBs6e6lriRn4ovaXMnqyY9uJrepNdxRp98CkgonjHxnVKks/klMUpxHM
XgkQCwJXRnmJgPaCo3PLq1AxBebiJrcNI/5XrDjx2O8O0ZZb+1306p/OVHK46nMYaaRr26AHap2y
rRh3Rlj4OQ5rGvQadHSLLb4DHZjfRkJha/WsBUlZZU0CnG9HiiPR9K/clRfszY2azpfZlqR4/i1h
BrW434CxyDrXoRDA+CCK11Gxidh9r0qsCQbbZ+SiXrRkPFvvFM+6Bdy21ZIOIIH+FmJESIiwhCiv
0WJnWSfZ+CKvlrfFFYsETMIJEGcamZiM895324J3LZTWNZYnJ93V3ahAqRIUmHfel1ifPt3U47HD
Tk22xEgHEfEBp51jCF5pvp1JK8dpp350vjZWg0Pbc+bqSsut1Cfc7mmi4Snsn6FkCZnQU3wDsIM4
ENiGvWd3WcUUchcnLhiwUebh8tz0tE/4i+iAney3fFxseIbHy42OA/TjWtMqxcLPlO7LxRbBqdPX
faFlBf25YEUeI6V8ShrdQmuL8nAVxqgMU9wLSE2QNGruFTb3WtmNkCL2shjr2shusGriFVIfJdD2
3UlzR/bVnU0IddJ1Uii911F1LabaBvxqJFNf/SZVORppYFmizmpuokNM4OEcbJHvyo0erH27j8sT
Ch9aQ/42/NUZUh9hFdnGuUqLn6fGCPsjPwxVQhGLijuCr+lhujIdbWVeeQedDTrYByF67PZHfSx9
xG9SjDjlRxltVcIT/SSvsE3ByAka7Y+tGX9w6jL1k+CSaTv8X1gg+HidBiMr+eYGJY8SQAYgbFb3
FwIOi4LeKMWNeJUEr3XAH9ABhTcSGVAm9sRhozSVz9ZM8etQgZLc2jIax38LpdTt2lvTUo7Cx/1E
g64PuJ1B11x3tNyTbgZ/6smObRDOFxCRVu/kGWUzNsfawfUuT0PnZL2he9kH//DpoRJJ5VDyUNwK
51m/VPG0p4olpSlKK5GuAJzS+mwn7xS5B2515jIyoBoJS6jEO0BIqscnz958zi6Dm34wIkXEVCzt
ptOU5U1oY8RU1dpQxG+ibJbo5T+qVT9+34m4fzxF64I5IUzCCJe5fY3nJ111m5rnhExPL11nSRme
qH2o8XnfFLwmuNd/n2Xt9QCv8bQ3F80qA77Rz4U9tI137fmfi58DGTz65BuQo9gfFNVJtss4HV8u
gvTB5gBvLplK/rItWiwOPHN0baqv9vVg168q1WS3ebOblaDHOjX8A9zbudEQjTg69VP4JX413K6U
p5c2+CksRE384NB9alMLACmImSFn7MPd+mrAgegbk2eEkh2IgldYQKhgryoEOM7KUooZ4qfoN8/H
bx5nrPhW5nj1oVGHxiP00GbwwSY1+TpDt13YlPAjY6PiHCpPyxrP1devDciLgIDuVgbGIq8nXgIx
Nu6qNIuBFCb1pQlI22emV1j+vPBKHUaxKXtSvpuv5fiLvTR3GWSusUoTJqRXuADwR8VgkUcDDmiW
jbd+xhqHvdLB/NFANFGj87UH4iTDbaU55TRqVh6oTR3n/mVuzzymcNUrYI7+bROsG3jdnc8mJmQD
1th4Snn9N110VZAwrChBoGvWkD7lFwEXCex1w8ZVY4jQuM6DKbSKIO7p6CsMz8/k/BGarstvnJEr
KpJl9piYTWWM8zZ73bFJPjxs3NEaML3CRlh+o/nWXkoIoFPvsRekgsUlClxKIHyr6BDuxMOpIKJ+
v8u9oTGhfdsBBS4De7SdqcmSsS5SRvIIhzv3IZOyeySSApe1qVxPZePLCRcvdJ7yCT94ZkfS40+6
+VZPk8SpSJI2ZSW/oGb0uN1lHHMG0uHIZEW2BdSAAYSuJ7HwcDx9frh3TYfOx4NCG0i8wWCnLT+b
dIaIW//Bo+9z0zN+P7C1oQ1n3c/h+Fd41GV10XYBv1IT079dGi31CcWx6nAfG+6zEg8Q2jstVUgR
KAwVreoAIrlPW1oC4tZzEW9YuIMHTT7R/3fdWG5cubMiFqopqLKMOrDf8IOm/YrW5S+p17Uv2X4K
ofkVd4+YSedErtV5f+I9Crjr5xHL9BB1jgTg4bucHTYIXhLM+MkZIhTCJ+B+TWn3YXb6KPxSwSNu
I3W18qp9j9eyQC8iIqD6AstXurknxZku4M67AobJqYpjEgepgenHcDzDuwLB0bneiS3aYqYg8AK+
HPhkJvQDHMIFNVjDJ4WLdSd2JytdSaaFdTu/+m/Qop/AVGIY6/BByVFVVYljQ3jyrg7ih7bxsuHO
yiI8MsOo6/UTbAP2zD1I/7hFaYOaWMtTe8jFgrQqGIb0Jzd7ATczJ3x2vYVAhZCAlKpIuzc4FkgE
0cIOqmIHyOXRVct4ZCXr9Y0BuvK+0wpl/yX3m+JWjWeMNl/YTiTxZb4QID3PlRITETs23H4HBFBR
RApMNNt5XnP918WC8BrieymE5aJQwKxEr8E0Vw15X+U5/NsHXoKs0NIkPJcMO9bjpe1ypJGV4vtf
RUrDH1C2tWF2yLI2GMRKGZ6pxtvOgF63LlLNHLObWbVcbngGSD9sSKEPS0yqPg5aDHuSRzUUM6kD
ps9jzFNWmPpNuSs2X4LzpF9OlQmwah7fONTPmfCOKSsyqtGaaNHugKrPmvIp3ImUnQ534V05f7Pp
4AEJzN25s4i9Zlha6tKAMWY23din8hvupwoVFh1QizbUKQnilU1InSNzeuZKaT3wk4FE8PgSjjHR
NwQ78nd94LKJBcCW0TOwmO/rVWOo0k7Z3Iwv0gqrC+dJjQU/wc9QSkPhZ/XssOFPOSVHE3p8FxzG
fjnCm1c7LxxO/Rm+lmSXMFjd1WFXgyi3cSlv8QySrsEW5kBlhvLD6hL7xknvr3Y9++maE8djB9FG
EdTq/2rFtZajx0SlHh163W5MnnTq41yU69Yj2xEo/Fv9Do4GOCatQZmHvSXweKbDFoYU70dI4TE3
JNAZ9WZ4HmPzIU09uXhy+lWw/nBCxV7MzSGW7gjKZw5q9dpD3i2UdisQoH9STKlbwlvMO5HYdN+1
DkntWoEV182tPGi32Bm19lpEiOyoKOkPw3gCKsUcFnaoGDpH0tMHfsUbzE7aT1LTTCexXNUJ0XIH
9CqmlNkSXMNImyMx0LWOzj23DvD5EbQnZ1GUZXb0v0MrVtl1+uQ+UHElRjj1KP3eY6XP0/2yuOpR
6o5Rd1rdOYmu+tao0eiA9hOUfD0jW/WlE22XFwhaylIjvarTGpQT+ESF6od275sQaFaJ/raLDerc
O0rXpEIUaUFzQxk5Hn1qHTysJ+VSUc70uU4qoyZwdbYMx7+YoepgBWmVSpstnw1LeOYJ8YaaGYAD
ef4eXH1HYu3HNAlaShpy4zEu/t8TdY/eDiRoobtThDbMJNnRp5TB9F9DoPh+cdvfE18oUVOT54u8
AgiImLDy0Dflaw303frhHNIfcIc7S7JKtcT+Lsq12jTZhBLfah1t+jpeqlYT8AltZustc1j/XXbn
LHudcLBoG+E6IEhkPmC6/ogygz5k5wddy0SM5rBsssneFYHJH3B6ZgJK5L1L1XOGd0mLMzK08tRL
w8TmcvVEZxvsti3qAKEMplhXtQw5bOfUaPSGdG4K4hWau+B20Z5za1wqZDEqVVpYJ5YFwaM61D2m
h6fUqzPGc5warzBGtYoza9bIehIg/Zsrxu8eD37NXZHEKPfS/qn3K3OvqAx5iDdeYMuophd/daKe
/fnsLFLq9AmUuiAU+sFh2pLuT4GhgHRn28zhiFunIXLzvWAiuRApcErrOaonp6hWIqRttGPywlN/
E6YhtG9DbFGzrOtg611+k9Rfil+zytWblBghVJwDrjq84499g7+JgAsfIfb/s0Qn98HdxuTbPs+p
YqKWBFdo4Qn4HduYrmTylvGPqiRsOUjmNorhZyr2yb/gddy+Xh3lkzcfZ/HD1bgXtgCTdsKmXju1
k8mHYhHkdFLHD8xBEkys51miVCpmAqug671TqgYl9iC2ygzLcH0Os+j4mWCvjjRGG5LBtaIAoFYX
9bJVtNhkygJyYCnRMw7vR4eRM38G/TbIthUD6gEjA+/PXGyUmZpwEJdKsoes20/OvlIAthSg3WPt
FIA4956cejBhpLg4RGfSkdKaPxNFT5m7d8m8Jt22ZxCv11gnJ4LWNAjdU/ZGKZ6Q5FNcw0bZczEO
sK7YTmO3CkKxBX3BgbS+ddWu5BPCZB7OgUdP8fVgC0Zt6FwvXBl9Fi0AB9r49JQtrbLXqYZWSmG3
l2lqIXnWYPPh1tp8GLiMJTNInLRrnvyQFjqkOOLcTQFU5qUzckSzqRoTdTd/TZpSgq6zRV4o+e2O
bQoK72vBQUCX1yh//YCaCqck0lAS7BbG6pIBk/GYfk/VEkeJ/MZWadN62NEAPekhT0uid7XQ25fy
BoP6YS0HECX6EN0jiWhY6C61bR6DrhRxvIh/dbRLMNQXWnT/8EqFOgFWO3bAMzCf0+pfSuMoNnsN
ToL1pTon4lbqLLuT/h4KqNib4UxeafhgV2ucWTkxWM6sTCYRwzRxpn5zv5WDUmbnlfEcLsVs0JAS
kN+wd1tDTbiE5UBl3gmspzrWAwV4iNXYo3AaXkkbLVbS+V2ONosKW4y0UU1NY5fADmpAMi0FMn4Q
vajin3QOLrj/Dzu9kBlgSjl+e7hfENMz1bBZa+1H7QOe3e0p3SKrw1a1fr6yt56ehCtss6x/pVMM
8OkRZzRr4ObGHfh5o5DP1qTm2W1k4eLXRt9VNe3VofxEvrb6DXK5oxjZATREidlhUNBEZPWkBCVl
VpSItkisibwEinmFvuwmtEg2qNAI7HdGd4iqn6xCyOJ5Pz7GG/+izre2daohDpBgY95ZyIwPjztL
nOuhTBiKYzmTZnygjOAMWXm3Y7NBpUHrkCBpbB8tj5yUul1KVYupa5Ak8IT9y63ddOtfpEcoAUD4
jiAZlU/PQ7LcVnD2JAoLlMmkngi3EyzvU/1+3eaxYq0Sw68SQE0a5ILF+/s8Q4ESAk11onuesEQQ
Dxjv9+OiJs6najmuJ8pMI094a0yd2Ic5BcFDr4ykurMAJYUbcu/xfER3LdbPBPEUqHH1cl84jA56
uAg3/MKWeLfE41wZ01pC/2o4x9ETqXCicmEgt38fcfuJHHBsnz60K3EvLGoCfjVtaiwRqkfYacCW
WexkZOCGCoyUUHg88EdsoHYD70bnEpG+gWd1VkK8pazdw19vl6Z82RxKDfc6dmVZnvtToT2zRfeW
2QET9l+FTCgEdnuGtbhyeVcQE0LMr7KtadBVxmIgTuBLxBQFe7snEelrEdXzB1KLE8hPkUb8EPq4
s9eN5np5Mct3/OvKbGfzfF3eCDYe3TTby3dM6BZJEh6KxkV6EJFH/bbUUF/nXHQ2GgOYDbtA7/5W
Tiq5tWSjkRySIqHlHs16iXw9joGjSfe6hH+2YyMTOo/3CPoXJMZoCnO5BdiIbY4KBMyj2rC8h7kJ
LvfO+76fXMo1sVn+gjz2i6gMebjgMp2lNSOPhoDTX5kriz2D37/phxtyuhbqVMCHhmaRN7TdUtSa
oCI87o3etgQS6ap+BE4BsBm1XUvBFYoTBWOKURccEDeU0UyVBQkzxYbdAITRDZhBtJqFbX3Yhfhr
0bW4mSoVoc0lCzxZrCpo9fNyEWbcDa+mcKWUkL3MkuFM70zu4qTeCsLo/FA1pTVaPXl4Va/e0TCC
yQpwkO/Ka/aJ/rFmmqWCgTynTFNZjb/8/fsX4WSDBN3axukj2heae1Ru/VyAlNfwpxzpLt8+mzi1
dyQg00ssiK/FumZ0UmKCU/1NgPimofEB1IdNWWyi1XyHjOo7mujpDf7+J8162PHUtiXTIixS+is8
HFo7xaD2UIXSDbRV7L9x202WTxC7alJumnTHRGLxTBz4TfGPtHAgpVBRzOMVkeZsll3mZ0fNHUpW
kuN5wovPCgvyIcJFeEMVh38/U68lqaJ1PCrCq6+pOoDLT2zTTRSKhkIJDPUD7qSwrxFqhwHyb32H
RaLvg/lGo8D4VBlnp7TgdJkTneDgY9pMTRUO9Fh4ae4qUn1Nj95oIKAatRNUXx+JeeJIhKx9xhtT
DanqFlXXMKq6xiIUrMonBq3wXMGTpOYvX/Uwb0uN7v+IhHQN23gG7YvhQdAzAw6qFvl2qxUz74Gp
Qpu2HaUE6VhGma3jYuPlwU4DaXNoI7dZkdW717KisH+bQxvP9fZikfezySO3daUNdXj/JyO5y27r
QPoVW4gIuKiO4EcA1lN+qOUVge8Gs+ioEx1VAGTRDaTrksR0zV3Hw0EG5PUloqK0n7a1LTIzQHJr
JcaawtVefgHPUK12snb+Un0Ep/L9zryi2ub9ZfjcZoS0742RmM9yqFB1gWgReYfWhZQSjTYZNmql
lDqiHUfr7I5psLauOxlS5+Ib7jRGro8IaClWlqY14NYRWqBkj4yXKlskHzBxndciiW0ksotcjT5G
mIU7mH/KFee1tlhy7FA+m2Sv4MA2hd0Pnq2CfC9ea6KiDXmOQ3H4kDZ1o6dMjFWcTt62TqluvvyQ
kTH2/EOQih7byt/NXY21JfSTVE7pMDGBz0ogYTveL1A6Z3l4gGM2owYgkPhMRQcQLHpfPDgjLzaN
SJ/FDiU2xuCQ+BN+QYPajbSiZUxuHqpJ7SQAKs729CrLLJ5Wle1cuQxVTYY9F/srBJijMv2vMCxu
ygT5y+rERGNgZsu6ntkBSAQMZfi6A+2F6TxuT3u7aygevHn2mnf0z+niL96+j0VmF8AuD1jN3yKc
6yInBD0NkCi9pWBjp3R++owJXEP/fO/USDBh37j4BvSgblwKjCw8sH55VZZUBl9ZDYZG3RJRIOZF
CpOA9RJzeR/IYNJ838j5S9zNa2bxmwf3+QXVjrluYQjlAG2F+Q15N55iD+Ni7ABEPF5I7ZDf8ayQ
7oDWVBdJ8SBjLOl0Q9vUHge/qAaiLwPibU5OflR2pgxd24s0aBAjUIDOcOvbroSSWzqQv++eIacg
Q4PzMPdVvyShc3KBA9bq/5kO4k3WbE/u+yiJbkvGxRBCkYLBaI1aGgfmA+dgiJDlZJG385lhSv7W
bvKUE5Odcff3kdz6qeOiYgEnjHpcRHrrf2rM69y8UAmwOMwOmiDtglytz5F9qqn4pHPb6+yy33hz
8piVNA4zQPixDa0doGF0n1lhkRKMJYIZOVitkE3oxIoXSvqPj9r6OoDJ/s9F/m7wAnYXP1oXP7H7
KQAUr+Wc8IhQOHjQFfoE09eanrF9yoeak4sx6dcqdKo5iC6Crmyu9oTTlUKWFkOCxMeC3JR60ozN
wtyvVDCtAyz2QTD7AIr2V8RBhJmCYuSy6TQzooapeTrB823P7vofv+d+wiU0hXcHYuSQRIpHL/zQ
GuYvKntiveEk7Odim+buOzIkrSlEaS0RfHMQslQBfpDOYjRN+PXGFCOd/npkLPIUYbrCpARQ4ET5
TWtOTjzGKdMGGeI/I6HAACMJ2nDx2IcC96BNkwDePtViOKUDSvTbuR6owO8Iv1SyCDoYIL30pR4i
IK+w5vkFSwjUlWxTZOurAFPaZvK13/s7K+ms3Cwy63ZUz0LvTnXKsjZPkdRjhVt5zd6RADwdelWY
EGcRQLcyYYio4JMqR6YUpqynIev+xC+s396Kj3WnTV2RPaiAp5XogK7QEyokSQD0ncqZxXzfCX4b
rp+k8HEITyxG/UCeT6y4eV3F59aG1OmaAP22S7s0KF0f4ZZQADSFB091hswYielG4mMeoVmblqFK
bzoGpKHeHZqCAFj4+fgHTlVXhAMigFEINlCq62RK3i7QSO+K+cHet6TJjFlGiv8iqRf5JREovF1l
ULS7mMucI0Hac+3U9NBC/FDp54SAXD//a+TCqnLKdFyetPJ9oGCWqu3Y7jLurfPXheYzm7CEovjB
mscBuIotLTMda/tSAPkzsLgzYukr0T/e7ooDO5MSzTxoEdl55tGognxmaGUNPIcrgsH+UYMUy6dj
20GFFXf7EU/ZYx2gmVsONIPiuE+kha2q4CZcstwWvtjGfefCuHxZJCuVEQblQcXAxj9FSamhmfxL
86+B+1aLnvzolwJ1jssBalvYGh/hv/Lh/EN/WPN7FAQeYqu7JMBXac725mIX6U2C/Pc8j+XdeGxN
n8+eIxaIgPQA4C/vReF1knZyvw82VKURQlOiTsmlQ21oVtGHP49y7YSAaUnGB+NEqPtYeRhv8l1i
Wx8bfx/LIBLWMoPvmbvX50hnAZ7ZYGqLNmeJelsxb7/jnP8AodERprCdIBuWkZmTXemqdESrHu7D
Ec+a32NhuAJ+bDF0oKrs/Z5iMPNgBHcssAVSZ9kmrOSLpLYkS8HVPcsIhm22Jkbq9rcNyjpUPciW
PK8RwA6174wTan35E9Z/r3NQvTHJQcTHAXMuGD04TXbkeRWy22LBT9ggYakfbyC0QwTWQJtsfBMD
RYDrbiA/sQxxN+zWr/oiblFfZNG5GdCZB7Cll4k/tinaFjiytwxvdZ8R4r3Isgw3kc8YALbbbXy3
JrfwszDeePJq5CdVQ/6YFrTlnxP+xUIWL2FvRmxU4khpzJQBJD5lQ5OdN2T2WjRQUT9TMDWPD9yk
qft8WNUWpqtxQocCzMwQnaa12RvRUdzDo1f0Ycr1vZvcfNO+rXiGbK3hFcUfWDhbYm5bn/QONIk8
zIxOi9cNcAVasvDGwWv5ZB83KyTW8dBcHjS9QQdxL7WzBDtCJBbW1S9NawZFHmfFU39JxkIkY8oE
82qepdMErJyWm2K2SPRVTTxzgJOdeYnMXFYOY4wY/nVJtlxgVwUmvUdmWW7n+tU8ysLipB+WLQhM
5ihWnfz3KyBJPt74DdbZGzQG5JOJRd3Nj9lWKstyaWynYV6SIe2GNnZoF3qpsHNz8vG9pSaDifYr
X76BdlvRxTp4QWsFeMRJExT60S79Jfj5iBoC5dWj9+5f6AO8V1RUSNwfKjtcXAMSYQvTd/P+800L
WVWfO/v05OcrmMQVVkF9P43KtfkbL+LC6Yhaw6kyqQ9SacO8NB/8BBRKixWnB+qLXSuWv7uRcLSo
beC5A3pt6vFxdBq2lHfXLnmjfnsyiRyNRCmsamBIRtPrs74T97qgqFCKOmHv597mGr4J7rC4vL7/
FxkfdkZhucTluLiqR/o1VepeRCJ0flY/15fkW7fPcGkvqHrV1N9ahBgYYivT3IohDm3ncsqkLesC
FC40DcLQUPSsRGgTtFCf4UyU71AjtrXOKwzNaKf4TYCtuHD5Ysw4BAE8EBwsidljWHVpbEwFIyIQ
h1AqhF9wsjh/oIUDtWdX5PtyOT0c+NRXbZc4dBjAmMbEz2Uc/r7z/kFlTY2TEOXnJDlsieTVeT74
RFLDeYM8JOYrYs55+FRWn9m3dHQaSRkB6+wUvAy0mChCRjaLHkLbRcE3Cav96HJPJMx8iJFsAk9g
+Ic1dhgm6kHTJhOu0DoQhk5HkAZE6FEUpfWGyG89iGGkIydwkt4knYTV7omxbIPxyGiHnBsQWdUy
ydLP1r/h6StA9wGTZPVJukHAUi4xjRXn5g2sECHKlWoqk4H7geV7ZWGKZh1ZCxGwNkUxERW3qAjn
yTurqPu0FRAEipS3CrvZRlzprNHYCyEGzEwUFLYdC+keZY93RVWPc98EaaKWZHKA5zFLEmkNmIYM
jXhLcrOwChphPu+Ywu50o3ZRt1YhzQWttQ87pT4jO/qQoUTium5NYmpWQMjCq4aIs5w1MI0+pyGV
ZXSxmDd1I/OeD3oJd2Y5CVmjU0zDQOUHRP+6wcuOcFHJMUwNf4zFnlPxlssvkL2/FuzDtSPvHClT
bCtdSxruMBp3p1kJhsOhKOnNPxKhVdwj/SKlxdBlZ6w45C+ML/Q5qOQrMQu9OzwWg05dWbksRlQj
yOT/jULfFLXlrNeAlh/Qyn/ry6XAsPikJJSJqfshR0vOZorB9Dy8WEkkShnJk31wQDWbWqzU1zkO
6cbmEFKjpj+D/+4MjLDJLQfnKVZz5/8Sv2hPmcXyO0Pi4f/kjH/34gW8Ve+oZHiooCcbo2K1CYtY
9o8WbbDgndKQgSHKPI6C6bEsAEowJaEYgxSBuSpupLv4pNMhB9WAIGdbKcsiyPxuzyymJ0bAhli5
1St8adfH5f6SxoJi85XniPka3mUVVyL41JYRs/Dcay06itPQgYTnlzJvy2YB+/ZMjSktOG5hzeC9
T49NSyBFwADIkv4EyfTJ6qOU1Lqajlxo1xkOa1pOkRxSRsbs4/xJSwNwVJqL5keorarc0LFS/9HN
mSgCNOsZUCt/Coyw+bJsV7Df0fnrcMpKs5BVVDx4BczL0NdAdyMSvZcHMNs3ZLGpOEcRuOc616Fw
eeUwlfdRHjnALkgkbDBLf++2MxksqlDwh7DDy1OcT+dOc/uqr4fS5Z4KgtqxGoJIO6vJJayXnX1i
+/CWohwgnGfm08ROEYCAYXUf/NFkPk08Rr0lOeUxHubyLBQ4qEX2voGwF5/z9dMcVLwu7Gs+hGRW
U2C/OMergz/bP7C7tZrdZRCSVfFmBuW+KTik962pN9Ruvhb7VdqfCPIOsCdyyzYAb5c1XGdYAOlC
Wi93CtZMDq71f8BgAY9xhMux1AIghVyqjvQh3yxpHOdTO+EJKwuUtRYB0/DThr53muE8pV5VKxnf
3oHZmu3CwH/ERginZ9uJ52qh+tuc5tGheypDGuPzRYPaU5JkmIkMhvAvqRoVq7z8PIV3mdmaHCQD
IPV3NkTHSeaKPdjaWHoTqw4506IjMgzaIPp1VlbSrAJfhh/JJI+u/aNIPxQA/RkyLfTHcH5geU4E
psm6tjIThnjBo56HFtAowKFriJmBfX8oz7nNMg+lGDYLogoMhw7cV4a4amreOAD2RA/jgos7k9Zz
KATKPvuw/A9LCLeA9/jgceO8kHAtdhJq+VeWL+99HfWd666LxCdl2Q1clxEg4GyCQoy8Zipx58mP
nDEHPhAlEksmPliDrziBBT2r5vMcqgqY4VphRuqAKFdJ20Ru4lGW6afG/wQd1HsPvEKCbTgfiglX
mpFEQxp9P/Kqxc7tBbmDDZIV7oPD8ps+A1nbHDQeAP/GUzY4WgVgSdrICsh4njQuMUIRpBDxuvQC
VStylwokuk6ZxdxLIbxeMzzr71cNTyLkiMg/OORUKTJUKr2lAqsGt3rmEjS2a7EA+MLfSv74gn4k
Nfa8sbkwwBYDfBVBBlqTzUGkt2R8ySDkqv5Y0PF63Z5Us03f2d1TuphYQt4cFkXDe/ieM0aKGKx3
6V9JsC0nj0VrCxldj69me8MjtQDGgbXKDY1WcE35HGXLe85Um6BT11VHFkMHsNIjKE4NZGtqGebi
uWarhl2VR4QMpDdXmdj7FzPpO1FIx+nmkQaW9zggbu4XqeHIRC1iu0GTkoE4LDOzj5zOBi6RdQc6
izvQSmvnpEPpwLPc8lVlDO//ZqKuJ9nOgYsNCwkIQxcDNFKAvHP1y33I1rVer69EObTiS+xDLHXW
Gcfun2JtywaHq+NbYlYHZEZa1iOu30EM8Yexfj8Vqo2XLj2Vo6lbcQ0a99+X170JTpv7/20uqXkH
DFWH35JUezOfnQcE6gBb5kVj8KMNKlFCanFsFVNerrW+Ntd5e/E/q0sK8qLQ/F8Zcxm7kCykBjmU
/kI+HhdCMruPIlzLy6MQUTo9D2KJiH2GIxbYKNwyhxD8e9dZ/UfsIqJ6irQCFCdL46EmJ+u4QMr7
wmtztoRY8Gk/K3j5hIKHSXNYzk/45dEAdcnGge8tUGWSggHyAxb4KilTypMrxdn4yOC9BwuqKiVY
mVWByOca2n3RVxZK0Cn8tuvSfDahJ4XG6zyx2nM82UUfCa42lOZsVDclkRUPv/1HCVDiWkd8/E1f
DwQ3n5ug6Dn2QvU2FpNUJ8oACo7Hqr5pPo9JtKCuhVFGX84FhpwIUGkAF1d6GKj1b8LaaMSYqKIL
dSgK4Jn4lu9u0f5i4eMo5n4/0xZT0AlAC1KsmIYK+MaYI2FOCu8E+VPUKNLnvG07t3kOyKlcN1kU
AsPPlTthQON/AydYm98hqcAAd+OufsbUTVeMkau/3qj9NnJM4RDNsYStCvRUIaI3iIiXWAvZECpc
Ec1HmvHKE1YPcYPRBlLNPw1NVMcCMKessqjjVAiIup5TX/2Omou+nTAUqrQIIRNWkFmEL5IZkQyO
cJyUL1cGtX9jzvQH42fwQY21hUxi+TQdjfkVQu9jfeUVQZngb23we9ghIXmMtr0KIrzUC1fZIXX+
ES5pYFefZCSnGnsZ/NmwETdJwquKXN1Nlhadb7kt2VDRXuTWeWZCFMu56j/mADXPxWzor2ERF0ph
XtjvH+Wjh1XnfQ+qfmA4J6UjPd/M+L0FUo7CYxH42UiWCQCmTOsupQ3RoVAeUOfmGoVzlrnOPNDy
m12jhwaxAVDFTScaJ2/5d0MJClWs0zjL6XJAxkBJ50cWpV01DhDvQhKOyXpiTc3aJKBvy9+a6usB
Prz3I6js3rlZCNLs+EjZCkjERMajrmv3LqyOli3JoC3781SisSaqAjKDG5btSPNqJeZlY9fRNFn9
+NBZydIJF6871XVukPmuDHXOJ4OH5dqknURyaDLTBPUn27LvfFNRKxJsg6WIBxiGyx3DHboOgUv7
p4/my6TTnbPz5OD8L8aZJqxS/Rxw0Gi5uXCV4pePiaK4Wtf22iD8Zg9FFroAQkMrRHhratWU8//Z
MFj8ZOIkmrO9gfncs39c6llKgwJu7pntWscws7XuyEhChU/MJt4nt3UoKAIc+0ZBATajRhi6NemA
7wECTqKVGjF+GD53pE1c1p92Kyky25sqoQDzJrGa2ucFudJFI42o7BkIgwVamrzrjBf5hb+GwynH
NBGGOMMX7HonXFV2kEnIp0aypnOvWH6o+JIrA13utSeOCNaFO3F1tcs+On9ysXLJPJDMsEcaJCxd
H3JB2dtQJIHafQQw/nLSzB3ZpoR3cjyjWYea+4hBoE0FP81Iy2AcxSauaTkAliHUvLj/q+lGa0zq
Z7MlnvGpMmc3mHoeVrRNTO0S6PiTDtjFB8MGzxL7AQTRYhWnnToMU9Ta1cOF6fx2GQgawdkSZ9K0
UOppW7yGFwEjSIFXvmfudcsCjEKRobl/FN8aPjrnUilYUv9EJZNXCwS5qZYNwH5XqeCZK44zwa32
Nk+k5LGlYKgh7FTdaD0qMQGJXOrPtX3z22pxHbklYD0QB4x6EzZ4nImrb8YeF300ZK79w5Cus8RP
oAW73kR3ZYZflkwKtX3Kw48VOyV0Vpi1nduwsNKmTWd3PxqSOSGkFYlFYWPKq/8a0p+JagybQ93N
ysj4UY0JgeqJgNCfJI1Jjxgi3QbHDh+EtcaCDkY2FdNaSWnR0CwOSjywJfoMqSJ0E78JHrVHLnr0
Raq1i3GGIpm+IZyTNRYmZpTeU4w3GVEFAygUDtUMkx2cmKCPIWSmNp09d72waQNeYThLDRAN6C5Z
OjUjhkRZwotGg+VIZ+s9xg7EA7hFytC3LOSzJVC+h8QZ53CNxiJZQ3zE5N+7xJSl74Z5ItmJ5mqI
dFW0OtQdjgnk9M4le/J6nAZ+Q2wlNGOgiBCe5dMZ3piL6JiGUF4MNuEzsjFRwQ91JNw4j5GIJrpH
vD3vfnubuchN/iSLKsf+A6kg7kFEntErDkcxjcsbQNRevHI19nis2LYYJP1V8Z7ESH8IrP8dh750
rDL3DY+jgO88owiFEer7eFYdw1YPdSP61NbEwyKKplQ5nirds193jbHNAjTkD9GE4nbXDXbzkUs5
09bUj67b+7Lv8DEduJf0ACLBDY/Yt2BTnoM1Fr1QJM+7y88+L4BXt6Es29wQZgF8N7wd1ZvUwtRq
9oNPkGFBWEPKD+zHNQBbwCmiCPwP2SGpaG1ChbbrTTkP/C+CTHf80EadoXBVgq+xJMfjI83DfqdI
tLnzPgFKSgqRJETVjENa6graoc7iSNm7FsYJxb/EiqUBDQSH0z7AQgqpj82S+db9f+onk7K/HqQ+
JCwox2l8gRIjEQwKxhjzzeYRoyR/ufa2vbU7+JAj3tDRLwK2cijTP0nnGvMof9/ox6NFeXNbLjMY
QHHzvpBlN/9IBx4eUTGd/YThpQ7qXNQjO5bpNq0XAStanqgKq+nE+YLRE3Dnkvq/qDFnv63BCCfv
9xiXnH3m7wNpEAwJXmCoCXhelXb5AdemK8PcErRb6luN8o6XTgk+yDqmuC+wbtckFepWvt+48syZ
U6nAbKv5lai7knjhAzGtgOCs8ypI1Sk4Uji6zq9DHvPQzYyKSGEeDpN7wOb8rFlArdUi3leHzaLL
bAcT0r9/ug+urrzF0CPhoGFhJCRBSID47NlNFEdT0ktgSVQcoVasLxVCGs2poOwDZB45a1y2hbXJ
51Z0RcnqYvFgJ9WtLvmPeG/CEs7S5oGne6z/1MDyGLahmWQLU+OzrJzMal2OGMA6B724oQBsiwPq
RklfJrf5CNlaMRKe2VK4iBDB6enx+mvsodGPVkxhwYD8D0vhOVjSfn27NqAwkjfOE2jp0jwi9MPU
yTUcNAEYa0r4cb0zYsU5VbpaYzFMjlKPdhGtCxe2M9NfTcF5MMJ0276tMzCAJilsKcvaCtxY4vtC
EgUmVMGUPruIMm34QMEnAX9qZwtJPxkt1n7XvtQwNFIvxY9nMornyctlQ9QRr5iNgrTylB7BKtkb
2zHGlM4dnlBfce0IJhK0Z3IKmao4Bn8O/TyLVpurWs7UZGYFY3hGxAtRQoMBmEawrObdPIwcQD4i
ZrwBl47Bft/SC29OLM1TZI6Lwq1vWvzkragdLk6gMf8oYYVNWi7rnSDqvms/knoy43U1IJ1bLNbn
zqAzCIXnTgythRMinAckN67le0kxLS66HPJom+M5I4aAxLCRyWcr+dGXxno3NDL42J9rNHe8AtHD
gEsVDt1aSlN1WRxQZJh/wcfki6qi1unjrExEicdNbO7zO/aYwyFFenaD/GPuU7mSXwM3TzAUojjf
xn2JBVYrk17MmwxND8O9V4XfLMO+MYiXqGTX2N1kJ1Ae6wwdiZIv+dyDJ5g0TPcsRlEo3J4/ZfL6
o72Ks8JnqM+tyE/P3jdDsce/FYHVAEkXkH6tXRbEFMXfI5YWZsu1dsMC1S1AJX2K/TWSDOzXv8do
KTIBv90tuuCk1M8ymPTOTwyEkZYmSpjkU/P852hKhCtzG6hZv15WNCB31rY4Z5dKRqFC0Ziz+PBQ
aSYcBS8tbIIdwZ9a/rGMkg/xoAVsLDkrbZbKWDT58Izvo0g95H+ouBI2ETxAySKkjMP14vBtBagD
AKo2x2zTOKsufyFrvT07eZrbMOOy2xzQVSrK33jQcRPh8pTFhv1+hDF0O3On1Pf8bloMYW/DBpKh
EaSpfaVqBEcYUmLO8emKM07htfIrBv6egDWDB7SmVOvS5Z1skuOQhLarMSunLUmaaU80zldO/wt4
JnCUmYNfhzbKwYDI8/Pw3oGv6NmnGj+P4fCz2duyqyDCPTVLz1WVap8uYBIyWSHsfe+Wjbozdyfl
/BIMX+Uts2MBk5bKDEQPgxFpTPcYRRqGoVQw4NNHC3OfQih8QJlokJn7oOyrRc1VdO1fyJVAimHo
90Ci5hFX4BUXn8VUXGxVOCFmeemRUgvNtKTJe6u6cZcECX7jxBkfnHe1wQ7y7QccyuusgL7RxWmq
2m+OjPWDtV6yRiRwZ2G1skt9DSrKPsm0IxGVzVWvK0NjE0QhD00ahIi31eIYF7lkMDfPH2OnXdZ4
hbc3NNABuNlCJucLBwNXtOJ0eJI0MkkKHKdpQAhUPwIiC9dQJmJOd/e65YhcYMYNppayb5UzB9q1
NzHdOC0CIPR155AjHM13PWQYpYE0zKcR2hM+/5uG+RwyFk3A2bScPZLavdfcHr6ejtvR1Up8FXHz
AuXlUjOk42kEI56Nf4z0AZGLH5CjFZ3Oyz6MWYmJya27oco1DmpQkzr6ILLcqgkpK1PVpZwXciWF
o41dGsXkULHz2cuIt6DekpB9MxjM0BqWExZbZDcUMNNmNewyMS2GCiG9zbSbibXj3MunOedFx6p5
uaQj/W52dAZohqOq2f9BhDsPpvSecm6BzSkbfvrgJ0MA9x4fjmAP6492gh7xbk/qINHLu3tWiLHw
hEwTFo8qbjetCOfrhUZDcK4I0PDJQDm9quSEfELZXWttQtiU2peMQ0Guk4/qOXrRLa92PJiH3rhi
uKgGB5TcY2+elLoKT/RVvP0/wFqDnj3jhKGdMRm19EqRJpUuQSvzVjyRVpc1nGzXxHehxmTPv4VZ
iKz3OvQ4jjd07RHiJZdie6er+IVUADGTNNDpg1aKvmE1pf1oTR2crZpKzjeOPuo0X0Hl5l4rrqBM
7ClgNIQvLRcWM5YSCNmxeY2iheCw92gftkO5rvxz1DDEq7SzUgvknZCEer/riyDdA4cdNekYMb2r
X3z/tpCUw9Uv5YLXzxh+0ogoIcei+V8oOBLV2nV7FyGT7r4Vwk5+k9UQKiZ9/DTo40bgnd59lKG5
6lz/uTwdZQ2lMTm0F3O4ijmALTBkhbmqeegXYXOJX0eJKXIsyXpx1wRQY10O6YkiwG2SQY7MSTIu
zVpvv+OcdOXiD/zoLa39iGlzbIWWoEJpcwyyh/YzWs95zKIdZtfmwtAOE/l//j91l8LKcSLiQ7P6
WVDQX7DCXijkY8ecNEcaWn3mSQ+oV7xnTuuM1bkt1/CoOEqBwr5wbkXLHXgqNRL+Qf+jF4pKyK56
rBpf6nFqP/qi86eFFNCjNcsYzB6jlp7WtMTsTppUX9SmmMH+V2xpDYFAaQCnMHZlvbnVCaEwy+E/
FPCESLRykT5vG66fmb/HzgrhvpsttLbztdKDOyzgbL9D2HdusOn11MIcC4ROf+82fsb+MXia+/59
JIWerThrHDd9FhhwxlBId9O0JCeNeYnW4b/icZf5zuPrbP6uokrQJaTavMMi/+UQYGmfCN71mEin
Li813+vUjZ9LjzMyyVHspSjSx1n0fBzloUg9H8iQ840UJx3b3h/G+YOjFqBX69YEksr8Hw6dr/1l
ACWiVn1vgERlZxjS8i4woa2GsrQGcRG6HHI6PiJDRLlCBQqT+hLlRGa1YJJNrllqslJM08gyETOC
FTcFP1FyWe9zn3eGbD01I586Fs83SBD6s3AMMSw41y6juQrT9f7l6LIRPs7gQ/8XKOR7Fy5OkjS0
R0JskHUckiF5OSNbjWX5U5qMogDkeK9liACd6Nm31lFPQ3Nqo8JzSqAC1On5BOqyne2sXW8bzW6C
hAn2HO3hk6xgBWQJCnTJjJ7fCwvoPju2r2FnlcihvAGwBvEEpI0B3a8Lu2fECteRzgcMn4f8moUH
kch5ziEoj5xrXx3w1OCSPbMLf70NqHUKQVjDI8wU/4V5EvGCSR5CQZlRgsEpsssg73ei2dfIpIXB
gzosjGeLuZnJ7Va0kKM0JDGzsTk6PR5ZTSXmV973QqNpbxjdbPNemImGj6stD0VmedO2sYSxXMmw
ds7jyCf02YFdLQOu3P/h+X9p9JVX1kiRy0B5qD/y6EVwCBupKp6xmYU+bF48qoAV+rbv5fCMIGKE
kFD3sD6hQW147yZuhGZkrCj2lWZZVM7fcmWz0vV0+d5n2TPSuey0Ed+nbv4BvWw2hPeiEbUP5iDS
n1n8gFctM27qmlhJFyEiVmUR18GK7/7zrcg+b4aJWm2x366udC3w1CJAG/e9b5w2iOPW0PsS07DW
goRzvmPESC5JjfIgmaWVRpOtaduMkFFjXBrJrUyMjeyb8fWQOLU6UETxTv822tAb0MYeyDXUyq7d
rtu5JpNBtJ3jWWjcJIg6pBZjFWSPv8yne/HIGaM3ODYnfDR0AfoLTY5xBmqIWjBsTEqrKNJwRhNI
81aMcW8FveeR1GK4ed6ocgR7AaLhN8g7P026+A1g959C57Rsp8zp9kYvqmTU7TwM50Jw7UH9VBXH
/X0JCdw35qcE1tYBfJ34ouIv7wWotpnwGWSQ6oJnaEPZHNvhAYLpRLR5ux1r23gd8vgRTx+SOy6u
N6Pl7gFolglQWSW5Ush9PBI12d8ba5jGteg3jZlJCN3IL5i5YT58CC9npTYd4R0iQPb5ppp9L/eb
cCNp0YCQtaoPf2j31/+D/DgbGbwFZYnyyA7XXjzVTdk1g2LAjSXeuOXMZqrxzB6/KkhdkcD3AqSv
29VoaNjfCC3FRUY/pXuvEPbV/8KIqa4XsDbhqi5HzyOD2OcaIqnKr0w/LHdtgAtWwdR5ynIX5hVO
HVNpc6lfPxO1OYMexcGcPrGnY+T22QrRlDynp+HDZOKhkaY2hmKTq2kyHn8wd5uupliRYySfkxB9
Rbgat3KbQ2kBgRdT4aKUrbyT1um/J3EO8qvoI0Z4Qn80SpkX2LEwiKCvC/jbDtTxf8YK/Q0uxGDa
fqu28mSuTQcT9Uhc7v3DzUwxggz8k+Nz6FF5b9w55OIw19tzIctO/ZHMZALHnqRsvwk+2fRKqjsu
3GOb7sHfu7Kb/SgabLCmIHrhrcui6KbiH+tLdZuSbP5xleklYBbG5PwpE3F1CfskVICkrGwEUgPy
QaJ7A3ibSkCS8nuwbRtSWWiBhdnQl/1qww71H0IHD2GOkLNnm1Lc1k55SmVYoIkeJWZ4skAKrMqb
Mlsx+6rvPnLZhoRwLCGtQJgzbFAPfQ7UFRw0KPkZyKtAdNcNmKT8YZCjCquBz1ii9Y8YooZXKcO5
1H56jlLzD+ehfw1Vhq7f7R4saSNwr5uTXLSnnQ4l3aziqIOKTyOTJ4lUlaAVYFX4AjevF/m1QOAh
uL7zksY5ehMOMgJ5CCoT1x2RezxpmuvTxAYmWiY6Hqn6Kdzy7awMdru2dWKDJgN0S/zFHi1huH+r
7vV864Q4S56sYeEJtgau3fJb80bXHietttUNTkGVmVAfmdUDDk5GSf5/VokxcZh8iBBsiVBIyQFC
1ishjwiJVWRHgfXRUpSDe2QHfLGa1JT3eGmuITQmJsmfZUXal1JlAnzW1/XtjkjKho/fVU9LF0Hu
R21X4Sd92rGZUYQ7wKrte6UGsr0xFZjk2kUpZ+utsiWcKWc2TcFN9+06pMfZ5q8oeJcxtSUSuuof
27775v5yC2Q7hjFa5+BkZ/YLpuaRzMbim6zw4Mr0qVuHedQd3cSkzNFwDS4uRRL8wsI0D7QkWnmB
/uLSF+M8J1JOIKACsxC3Ciu+BL45gkLT2PIhK2NGPqoa8j3UE5vhnBAQ9QfoxET7vDlHCAn4ypJw
EvYNYUATc3/UP+4rbzdjPSkJX1Icb38WeoM0n5KN+zUhr3keQZ9TPNlRhl/CqFGBrna6ALXxSwiu
51hBHd3VfCas/LLdM31Fb1Jjo5p2NBU9H8Rp+kvNEXgXVxH3KmnZNxDho4TlIw1VATtKycNhyhkj
GPZzHgCPd483ddugJVYgwKUNN2uxXTypVqT3WN6jVghTNM+TDtH7pin8RDfCevpEaX4eFg7nBOQ/
O7JSKe0+RSMtpLU+uLhyiYebrLwH+TqnGcY3FIpRrfEjF4/HxXj00dCgFMk4pqt0PeRrO3vwlw4j
W6lpGtuwJBHwsG+FwanaYIhA43cgMrHOJe9T+/H6vYspDxkpQzFIHul72sV6V9VI/NPeBcSxyz6M
LAzphp7nXYcI8OAxmS+eTAYZ/+Qk5rh9bF4HuKqQkDaHR/92KmvGGfLNERmW+fZWYmEw+1Cz0Su3
oADPPCDSO6hjT4+I1QfzeEj3f8QiT58PlKGJsvS+Zn1R2FNYB8YxodmKmWLmSsEcyWIeMAIcb7X/
HoY9jJikg37SCECuZFm4XcHKh8+2QKcGccpNeLAXCQx2YqI+FuUZSuetu8RKIdYVKJoRoNPIRBa5
LY3RKDjPuNx9BzmzWbtfqWC98R//5yvlMV4wpu/wkXkV+frneEqEtdvq81adMsgVMGXx0fLNreCh
1sRP+S6Zo9uKFkNxni20H0J9s227IA//USs//3O5uZGRvoOgyz8SOLRLn9MqV75o0Gk3I+xmp6Av
aPGG9AMppGNdOOWNRBHnxpIoKVt6cBsgyX5Ve6AYxj3JKleMKlQ5NCB/L46y7UDAi2EiqQJ5RXrf
MIOMWMp/sSofJ9EIX8K2e1WJNxEOR2qmCdNsYrnnmKYhbjV+v5idbRlwtOvZAwsNtdkiwz/Knwpw
cYfitjKqtolTAWaa7RBpL5uGlrXjJWAsgJcZjKrayEWs+4rBxzzcWMYcoRByPWCb9Y9P2z8lh6Tn
1UalUoNTAdLsk0CTPDoGKc8dCD4PdLVrqWUZ02es9k2B2C2DBBSKX9Otp1l3xgfGwp4SRE+rNzrd
1sJSMg/7W0wXJfQ1XnTYjfd3+73MNMlhKzU96+1h+hEfEJ3XwmYuygkwl8EakVz0gykZwIom1Cv4
aXZ/p2SAlX/XbjqeIBZnRAvUbpbKb7XH+ehJ46TlCwB3pY/JCVBWCFCRZCp5vxX5xKISAGPNf5g2
h52mcpj4SqWoxdGEU+I/IKq9Nv6VItYi0srW8nj2AyIJL8VhXYnxFsBCTxmf8/xYY4RDFy9rSTI3
znEcMQ+cfC1KNSO275PZFeFCr7AlxUNEjjquT/+BUAfykHe5uA+73vOAiy+Pzp5Rt0IdPRHx28mj
z4SshskLoHQFf8h6jfyBAWZuvqgYGJ8Lot2fz1OKcQ/ZSQJlltSnxA1LhwC4Wb0TJsWLDPPVwthf
NbG4L+PF4xLf9w/ywBf3gwI6cH7T5oLC9o2i+FTJCv0PP5VCB07qQRXXNfVgRjhFA1lbX2E1Bq8E
7Mbs390GByI9iUA+NpJNIrnvXPzJxGEjzm8pBbMC+2Ee3ZkD6zEqz9p5qL429P/pEc+jPcqWs0Bs
5MsSb3eb/tREnNNK8U3k04W1f+4xe4SWNp1m2WnWicRqWqjPZJdZnI1t9t20lAIFq9EwGTwPSfOU
06mdgJVJEGocoNoox70DV3hi/r7aS65ePSQtkj92xPVTn14koggbX0i1y8tPXhPRJgSbzOuf9oum
nc4+T3o/OBSi71WQNEJQY3App9uaAl90bMLHKb6jyPnfU09jlWRO0FZ2d+CLZ9zVW6dCIBsNsYOd
x5dtX+klPVdhVjXh+32JdlBElAejbPhNscTwuI5F7Y46P9FaOxNQCQtU8CER6W0kyoN72CPIZcoZ
RUplmk63Yt/+4rPYTq/uyNomI6ThHO6iahxAyqM1gQlCzAiJCx6AfXSvk1SY7zgfCSDxh4qBT55D
+mR940dut0Kyq3zqM+hYcmlJpvzZnZi6nLDr07Vcb25pHu6Ap2o2Gotp1Ri6EFmPZX18Mjks1Fh3
YU9BENuBRu81+hIisUZvQ3n9aTEOdR/+GF2869yxNijtaBqBZ4ILojYrF+p9mUIsYSPqCLem2IzL
NmokIzqdcXrnV8DO1jSdhZBdpjl911586WKKTD0dZC8W7lLJ7zId5v4FT6rqqp4NylRZtZ0CvdwE
V7VtywjQR5JH7UU9myE9DfTklYryEsiGyYcHQhTmRq1BB3rb9eKipOf4UeBJA10ze9vZ4ZM5eScv
tqFfJ/LxDdjChFiIuUz5T1f5GGL53AKO9NyYQcHQiXbsndvp5siRYE8O25EALpw78lL/JDvSn+Of
LUCWYhpu7aZV3cfc+RVaNgEJw2pUZEaQnHqIct/Arh3x4ZyJ1HKPCBabQsRyBAQCn2isDKtlnpnl
crPFgAXJP8EetPvuhNMCO+QJyoIe4F7cWd0xc6TShk+dHq3DYepCOfs13yBoex7mkHgcF4//FChk
bBxyO4e4j4z6x1jkTobEyyHlQLL+q5y4ysRrzZByCXZlE/386ibpERxaDma84lUpvAmlyYJtdgtT
sMlLmRSdo+WmHmZGqIbr3oOqGkfkfE5ycTLMvdBJE8fCHKu7jAVgpoGI7ZSFNtTUNJi83cI5C94A
35ooddeuXtZ+Tc//rajn9+dWdRVN1h6byxdkFiD9wwi1G/mwjtsMZibJ8RhnjqKSH5I6B381rUJX
fiG2lg5ZSOvIWrclSH2OO5QWQLXlovTQr6cHdKqhcBGK5oMWPK7V1ia1z15JE+6nJJTf42C62nxG
Iypyt/4N6zeSlj/vNqveijDt24qm6fV8/oU1R4X50RmnYdygclFFUrj3ornREQ3Bad6Rde3JL56F
CYD8/Y+D+neKQL/PZKWeyJGU3OVRQrGKoJtyqtUDLk3FNXDULrhZO3Eslb451OjzJ2srRyLDSLvd
tDVMIqwy10tQ4T86Ft3xLZgKbjiQRt5oSjDuPLbGMIG1sa3kZbanv35hx0X1NwyTZKVyk8ngRYD9
6s5jbISqPDNMa/gaqH9dwNoM3StjtSCzH1B9eEpUR1EMA7OsbeWWh/6OkeZc5g9+yYdL5nou0Msy
qdMu6v+jwUQ09ca3SujFM0ARnMjobSGceJBN/p+4XLtoRLl4Cjp9WZ/MrN+8easo5z88iQ2lnxdt
AbAg8Usn7Og+TepExPMVU162DpUu8H+8U5tJedUFHjMrXCNR7UR1j8khhDogfrcpep0Sl6n4Tx+F
oRqQIFYfe1SneEdCueTzZxpfDp6WDl8n1cVmFw9HyNA7ISdCCO0jK0yGR6KEQ1Fyp82Txwm5PN+p
oahlOb2+kMM1Wh8Kyycldq8WKZdekgfhvgjTmSUtWOEqRBhNYR8IrgwRIV+dS5C3lg0Dm55KNqwb
6jbRAO1QPUzE9cbuZhtfIM0/47apN6fe9odTgakT9QVAgv9KamU90NO+SQh6p1091dqAA13Gp14M
GgIIlEimk9VP59eoI42hbjCpYp8KdjuIf+Ynae8eVzNRJpW2mIglKdU1mcTjJV08gXq8TJRh4KLD
IzC1q7x4R55hSgkG1/sAuGSqUI9BBBxOYbQ0VNsl3S4F2LXiL4h/dDwvfGg2/X8M/GDmh+tiXska
cBefUytTLJ7G/ougFH+P3XVHS5n78jYWtCkfWRGTUCl9DVHJL5wpX7/troHRl9QdIBFAvVPGiy7E
VRXFFCwYIiT3Yz8wo7AZFXrM6UCLtowob4rFOouh+aqtTlR2CLiaV5Hu5qeIR6YmSqeZSgzy/XSe
ZXcAc2yD+MmP2Hw6yKaACGVXYo9GsecKGDVDRFp0Ei1JTjgi8sYQh7tSErYENk9T8J92ZuiRE9za
UJdSTRagkeAqitVp0/6pRFxObeavXUS98aANxcP66hAiRxNwL5gcZOEdtlWTrmf4ftfC9iIiAnc0
Dg1eohz53BhYrnUpHf3XHic/ypYwMSOTMVwd8F+YgpNj2fNdkUnf0pOz4CxImgyqLWnnCE+GfMGD
iW330XzbiDvqfb+VguFbOON9i01dNVF/VfQ/b7Vije0+KN26Y3alMSrWP9Dn5VKSf9gV9HbYrl+R
OaDx4sjmvOxyCgssd9WtdEWF65tUs4JfV+DKS0XF8ULP9lUwSnNeyuhUzoZStX7zcqh7z9g+5JlM
euO/Ip8e9yYjAVfnIunYJMvL1vYWyXvA8BkdFIzNY4PBxssYW0hOoRkAKqwyTbjiGq5tA6s0qvcc
iMEIJpey/Ukz7+N/P98lwxw66KpJ47b4LuEOcycQGjThneW3iygEna7ZIuEqXLW8tsKfIAkuFSGe
PlQ+WcvbvuyjYzA1+BhxrqKu7LRaHrgUKEU2NyHKFuOcdeuN/MZ2VRlCkxX2fRCZ/bWD6b0Phk97
M5IMSh6zLof+w4GMVjZeT5o/Tu0l8LGPFrcF5AgvPTB+PVr7LT3Ganml5PQ/UU/5nieiUDpP1m3U
GvvT5uKPmNJiAfEN7YK3irN0fsvAEzg95i69qFZ8H3ORlRZgywi4MbMNRBF5KPzbEDEfTRJxF0Zt
NWrV9s3sT0uU+10ENebhU5paK6bZ4TO2pFU2hMIJ+GJ4p2RsJlNCr17fEsxDgGYUkTworomh/M1/
HfRC1gqC891EtnSHsP1PKDFjp1ga7X5y/AdTTntjXgioNwOwzvTtUQVw6Yu5T2ec/nSqBhlfyi8Z
6Xe6VrPIrzvcERLW3uCmvmGLhpHJBMSspHG1ilD0XHBJM0CT1RF3zIm85VIk8ScMWZKeIn699H0Q
GiMNH+kxzkIaNFOdfQLqyBCvIwDGR3diELXM/UfLnXKN2IcKhnhsOkJxXrCNGNofk8OrTubDhIn3
hnP1ugZBY/Ctukn8oCTq1Cglgz5bugWiJeFAsAkz6XHAD/WTCUtMm5nL4U0YZBIA9fPj9cUyuExU
HjeQAS02wVspXRynPcRf7YWpUzPMreqDFD0BIfa/ZEx9E9kBae/cWDDORJ2wcpUD136fcbUj+7m9
+E+mgZrjt8CftTdbGc76frsLm2ILAy9IpqySPdQ9GD72vqHtHNywEbTPb+Vy1TJSuUggQfF1bwr/
i7EYQpAJTLbk5aTiL3CFscgsoA5exGlDk4kByTC3K1YchTqKrrWEG0xrohXG88sP8HLRVlf2IcYG
UNO1VM0xtp861WIz7yVStENMp7rf7m0XaZm0lEI00br0u2Vu3fyATQYz0AODAeLRHMD3+WPr7NqU
9WFrcftf+PTTsYB2+rtROSc75POWYVXbB+B1zAKCkrrxom9faQ7Ac3Fx4XYzRxeAaSX2HiU5sABV
dCE3EAbXXG1M4HzetR11nfalfrwih1LRZXxY4dWJEY26Ftft/4gWuQxyyGy0YI5NMYxnXnuQaGlX
ZS422qxEpJjTTKMpSwj/FEL+KEOl//r0PQ9ttuwlm0JApDQW4n7LsaM1Q1Le61V0LCKW6FJe1nNm
PRFUX/8id+0qbhkUZv5yAE2vWKPV17TzaXibi7uh/3jdiE4M/s6n9V8mV3hKA8pLO/F1lALvLD4e
sNo6MDxI+fVESPTqtCA5mnyPqXEDLRhG7zw8PWh0nQfANj9Arrrf1jZ4MOiWt6PCujIm3WVkP7Uq
ErW5dMzyalD7JZiU0bcuz+L/5wBQAwmBqnJ8bt2P+cGCSyUVSue+o3LMntgkXRVMjomIu3HtKDpR
lJJQRyECdreya3+yXZqBXEM93aGBRGLhR6cTsjnswBO7lHxAtgnBJ5XGkgM1Wyd5o3hEw8yaAAyA
DVyIxZ1KvGWReHb6dcTYv1FoU1vhAypo7aRMf19goy9wi2VQZ+qRJq02J7cJA/5r2O+RBfu0eCC0
fnQGXZmWIcQ2m9AZT8Dc5T4l8Vu6IqzFAvaiHjQjShsjH5IFvC+FyJ2RtU6NBoZA/ujP5K0x/v7Y
+TdX2D1odQ3HyPs7tCMglCu14EBnpaJapJYxXJBVrnABMEdG99/A1p8HRw+8/qJ7MKv5zCncfro/
s/bRYrXuKiyOrpZQbx9knNtCdva2VTLto9ETFhlXvkQuMM/vLQIMTM2bx8+wtonnlKiSBE5uzj5w
L893/CMJ7HdEfhBrRGscWAtIOsH1Lhu8ekmKspXySJOOHdpYUAL7XbbUjy4x2p55001F7Ku0VGDG
OLYBZWWnpMJq2Vb7/3Dz1a/JzazQOp/iizYqrkkMtZJEE5JyrDCxiVngPljaN6mvsdLPX652T3Tr
nOLlhq2eYaDNpiw6zDysL/A1D52JQnSkD+xK9fJG8UbVrnz+N/H69etPLLtx+CLqHDI0VEf7o5bE
w3Ge6wQ4UQPQYQEt6Mnmh+wYkws0HkpLQd5s5wnSVY3uFF/pmORCKUOyaeJU+2OqDKIG6jSDtwwX
wCSUidDBfWSYgziks1//iJ8iZQri5HI8Ab3xJPL4uLLlFOMNLZOJb97VnYNw9LVIb2VfunIGv6Wu
Im6/w1zKnp3rURZ6SWUHoSlxGsoHWCL/AT66V+uuzNwGiXGBFMMLVNLPA5bR1SUFMpFlhpGUmwzo
Z3b1jHhnSlg6mUb+uop3bim4HN9r6bEYNPoUq+yCkc/YUqbiQdfi25zfjfjtgMgEAB9Pnumh/apL
7l3jPR3dCimmigkwQ/WFQh8xbe3XV5K53f0BrHX9WuLsq74YCzKnJCQRaXvV8xK0sxbJoV04HrVH
RoHgWj0jowShDpnpN5XgfxnNdVILymw2fL3UzNSk1PW9yWB420UeT5zydEc8DP912AiNEovy6vMT
CdQTh6hdNMDaaXey71JO+UCUsM9sMQxEsZs0P2H5cC64ue04rVzBwW0mTlfMDCQ/4ipOj0kuYZ3w
bK1owFHt9fzh7/73VEYfJ07XL2sOYJcamIbzJyb8p/a0cPmzH2UpLUzir8o5nHw2YiPJAnqeKtx3
O+qGDW7r+Dz2MJMg2wd2h8MtawLTUINotZzNymXmwTRyfBfOtKF/HnFGQs+STyKjpcp/pfsP5Mgv
6ZjZQApXAIu+SHCZKY20WY+/PVczibOjNph71Kk5MsnOqgMSSbLP0eJ+epw8DJMLDkr31JfnGFlx
yNK9KTwLsNBFBkHE+VxtSUatDviVlI7nHFc1bAA6n6e29v8cL1N+HeO15nSavpEVBkDHL4UmVhns
Dm2J0G2wZzP01XnyXyJT3mstBLGrcaDF0eJavJqcyzm8y9dPR2UAdyyIclFSJA9NBQg4AZiipKJf
npyoavkAKNw4KbVkaioQ+96xOx3/3ijvloXexVDOMJp9CsBjfCQqrSsAvpQGF0o85ESONGOULDdc
mvPDvptgT8uANUy0nAf6vXnl09p5Oir9/GoUwsTxfe0IoJYJwqCcRZ0s6zlpMf01qUWO+hD5As+O
H+4noqSBMoQLyLXxo52MtexoEJkIqbnNdxOd7vcwMV/PCmg0ZnYdErLpf5JOweiWtxfTuw8sY19h
Ew522I0uFjHKhc1FHGRLqeruQ/JBqHqBB4QutaFQ2k3FQPD6UUbJC+GCEkK3QUB1tLCLTRLTGOz8
fBUjrmU5M3x5TAzz0PfgsbFE+mtnNMCIqYIfIhZfsezOIxWMh+Ahm2K1lFpo6q8mr7IkcnG2UcaV
Cs+4vzgBiEwCtCO7GaYfXoCyju2H5LElqZa91W7Hs5TMErYe8QOeQ4ylUcecTG37ODSp7h6qkjNu
gOsZCsXWGdLhfczJaznwTQInWovMjwZfVzhamw2b1/u9WuMJbmOC+96iluQ4wt/ZEkEbk9H72hhP
w4ns+NkzV6KYJzQ1U56MQbrYqYDv0bSOYSMJDYe9SDENKUokVC1rS4wBJ4mp6bVp3SoTOwn+m2tA
zsrPjjy9zgVZ7IlvFL9c4lFyIiH/DQ+q3zJ0I6OGkrDimspmJrIPxzFWgN4mgNbh3Wd+5HoIJ/Mh
sIj+2xKJuHBp9Oaab2AHR2kdyv7YZsvtuJAMIPwa6bRl0V63RivucPUd69ieRKgfRmc9LagQ7GfR
sEv5J1VmV5lh22eH+6eVJyrRoJAbkoeQxiwjrARItHvhzwL7PGjVZnb9E614Jfr7yjQvtRkC20NW
E3GIiQRxPwfvv2BBefOCtStK6PrfuCtWwv16zB0gr5tlsuKnUGaZZQhzDVhcNYEaxTD/Sqsuh576
VVu+P9zVbTN3SkgAsOTk0JVkcE1KF4KMoj0f6G12carwQtOX5Bnf3rWnrhkGK6A8iOAMEk8jYV61
bECJvTngyj19YbdagZJ7Zdtf2WnWyx8c0VqZe8CDcozc+sFcEbsmEqtIH9iRwNJ5MrJEwHVwEVEk
CabCMQ0JIHQ2HkbgxkswAoGf1k6c24YDxbmf9QAGqLpMZ0R6uWXNneHWtOAfCwzcM5JV43+WI1OG
3uZ50xH9Pj9hlH2tWc2l49Bsuc5xb638u9yfRBbWovV8d5E4a/4FBf/RfuWAN14w2vzeHR9fY9Ty
8Qn8D+vJdz2UqFXktxgka4Ka73PNI5tP7Yi8AGRDH6+T/MHp/xDLbCBKAbaewoMpyhvCwel0naLI
R6YJQx+mxopYnHDMYc1g3ZtO0aC1WgNSyCPVtO65lVhpKTz34GxUAcP7PrLRczmKZcknw2uWpcya
K+MYBGtBVuY88Zf37vnEXIuVDF1JSo5HmWLtXbXLk1hqI7UADjqjIrmY8cJHQENUPWlnSLSYop77
6I+kXzoZfUBeajj/K+PHDD2BObkaG2N4QPmjFRA3D9dz1HUtQtjUhmlwGt8GXwkqrYF2OXyh3VpI
PF44bMe1esW7NIAWZfQXo1RwD2xkx8h0seJSZ/D92F8mWhtO8BZvh1/yTGOA0fLQGmvZAQbaI0x8
K7oRa/4ThMm4pwQ0CsZn/daNVjpEmNjdOcxXmVao5wCEsoO7GEYrQ0olnmD616S3bVEGlpQBzEdB
tt0fbD0rPAqdUUnWPqMPjCRk6309VM8tzf5A4kMxKOUF+m+fxvqsmO125JlYb6Pwq0jT4lusiO28
WSmaFNxARVsajXtSyhy8S7zvfpicxcoy7z5uEG9YpHse6G/gbFoHXwD3wQnkjKFb+PM/ViTBBIwj
zFQVhPO9IwI8gHEi7FWNusi0TFIOYaw+UwvMN2pSTvp4fbisJtIDpduh1SnoDVfU9WOEkgjfw1Q6
bjqvsSKzGxUb+mplAfpS8z2aCq760LHo2B2v+9HRRVLoULuzZqD4upEKsRJbG8k1Kl9pBmtbkX6f
+P/s0nMoxIPsdphNeUgNY+EHRB1zn673NUJP5bkVSNUgO1/lSI3TW3I4FnJZRlE18aMS98ej8UNy
rUNIvwr98yg15kxk+CpVSFZu5K06fOjap5T/espDN7pGCy762u6T1u08pl8Imb/Ta8QBmpPXdRRw
0HBElK6dUtEk5Sdmzp1R21NEccax+IGcTEq9e1EmuEmosiZ1McUtlfbvlwp0Ui0q6HPAPyauXeeI
s5juTFmRz2Dx+6h7lJSJBrJfCSGMwChR2Tgn/xF7FdXFDA4C5HG1W1aRBzFdBV3jMbN04oxHSkXg
VSnBptI1VpO5cniNj5/3lkK2g5s6gYvVq3w80/nz7iKnSt/msstlYlA7fmcU4ZXV/tILw7EbsHAR
wFJa6aRh0eSgin33GpegwYCN6beSHDnSao2snGNUGPGm38/S4bOlw3fdfJtfaCwSaD4LvVuz2V4J
RvlZNhuuZPMY7gt797PRC+tKvNvsbYpIxOpPWtn0lC3IW1yz9red8Pw29Vm2p4LDaeIPG82PtnCd
vBcy9YGviWQp81ontueUQ/mHWyFShvogX4TPFwA64kA2g6MDI2iDb9Ytr1ABPlPljRqv/W0mO82I
WsEJGadEZn6R41thbZ+f6CnWpGaD/joQSoSTSx/s8VzfWcY5hs2Ueg0Ic0Di39WCpgV+/9pFfBAx
jChzEi0lgXF3X2z2JSG1kybTbSuOncO3riqTKmHWJBMb/DxGWTuBXBlfBzZL2BbopncsMybJcJzx
VGmDGaTjrRYxsfZG4/XrsNL+vP3QMtCy7p+uVcJfbwioHD0G0xJqdljWV5E8nzh6pfoLyHUGESKU
HjFXdvAThvWEjaXBhgRxDNnRQFJvf+FQWcQFut9Fa3C5R2yKepaog4bLDeb85k5DgHxBYc2xBpHs
y0TPcc9Yxg0jtofL5bU5kCoE9eIhFIbQNZ7P4rQztrWCi6pRwhk1ycfjY0VU0CezAMaouFSR8J6Z
kbTTE5Bw6/RXMW/DYmK0l2ctIU88IN5+DSqvl3Pcg3HIuXeb5fGSV51QKatlbW+F/kZUoxIWdygB
9RKPKX/ibk7TjhPUN4Ts21y0y7u1jPEerHa7W5CNE5dc6W5yUl5DCG3J8zIapQWhvanNEcA8Xiqi
3ZJ/pi4D1EL0YCwCdRlWJKjvFgY9obywZpZHkZg2cnIRXW9XLJFbjQ8HaUyVs3IZgI2rY+sxjjXD
GeLg2/KYzZIiLiClawrZz6+KTQT5GWrRxKMGZX1GtE2Axydo2NbJBfPl/Mbp9pFJdGZ4JBVKWSQZ
wnPrpU4aJCFFyc/z/rvpdm1OKB9+j5AJsK7w9cj8HzyXkFQlrIIybWHkJvBSlv+IvjujlCQ/ysic
Xa4yw8Q7KcvfAyMX11QVaeNvpJ+Ac/G5IZ7liOi+5sjdxgl4D1C6kjb7miBhXPAiq+/rdLkmUBT6
mxaXswEEeYPTPNlTvSBpTDCm9BNOOs29aDKBiiCeOBMtNNN1WBa2/H0llqTzwH/MmDqBhDGhqUQk
qKj7tq0HLdROYkH1BZUdDdArfFoGN27jl5Wx2gjNf9ESn/E4EAzQge+2UXaIjIl4HkzRfbsnUH5Q
jS2VxKgt5DtNE9FSrhHEXl9WzOfOezdTnlxcmpRp+FgdxT5yORxPwy8N/tBcH/DmUdUito11SHvK
h26TyBwo5jZT/eFlXlVSt5NEKO4OQOeUFTmdeSyG65DOZLD2TRc0gaIA1uMvKd+N+YiYx6ixRCNa
Oss7z0y3pXZCY5UhXMkrWHxHfafjKoh4YelJs2dYN5fGL4G4oqRJyL/s4lGVBJV99x2RbSRxfXmQ
78uhK6hiRUnVDKCOUK8eRNR/ORAyRSkD7tHDSpOk/xZm0ucBbPb+dcRjhAJK3BJtuZ8Mnf3cvzIQ
DWeitaTqBHajx8wr60hHNHsp36lJt9XP2qoY4Uk9OsAz+dHVZ7WAYA+2YRBbYHTSwSbzXhdrz2E7
exKvNCq5MH3lGrhRv5fTKzDbgcDjfT2I2BAv2mZoMNPcG+nzA8rxr42O+JvB3uE7WJPcVeUBrsZc
9WRKgW0vVaKBiLtUW4+FJQzSEX1i+oE0j9uGbcOPGUEWHOxxIpKuFapsBlI5IrspuBId5ovcioVj
VAvUCuVMeUviM3WEjGo9+z6pMVPdjELkn5zHg2ia3CzrXxx/raLVqQcczwalXDV/QCyvo+K+ObQB
ESwR2uwO6kbrDaPET0CqD7bmYybfFImpF+Zd8PfpC7uXjp1Dgb/pjfPCY2GtFbPI58zdTSyxfmxE
lnbbBiZmasyg/iY059u9PVpZ6OUwT6Z/1/xs46wAgb4wA/ZEoHtVMwsELfAJ4qAKBEs4RUI6DW+9
SOn909Crcjsi/TblIFw3U0T7Akv+bMe8Fy1JWWMAo726JCtlGQhYBVA7UFnE7VbygZfMig3uyWR7
+U4xtOQp1ekTbadtmibMcWEXeFv1iwsRMtuRfuyTYQj1kMzuBB8Al96Tnpvx1CndSeGnuHvKX7gI
Q+Nwl5FDH6KQE5qET//61L793UJ1+nhxGq7TNMfSIeHLp5Sfe0FtfQb2EYtdw2Rrmz/L49Hdll9k
nd3s0yT7s/AoaAYNczC4eEuZ4A+FRSEiR6w4RrG0/HLL2gMlsLabYx+RocPYoHDoOm/1gC47+7FB
rSYL1dS81NCgzsu58tm8twqLhhjtOjBpQe9dzloJBkcmRUs1+h4nzYDTtBkVMZpl79yIQwpxMVGZ
4WnaQUM53cQTXnVVll8xJR6o40RPazCSUyoCk/OeMrvSFvlgQBdS+C9kE4k0PWrWi5MbXg87hNkG
eNL1y7v+YF+L+kK/I68EYgmqgjPMYgnWx2Xy6xf9LspbUJcmcbZYIiJCj0Gac4F309i7A+NpAyZw
OZp/BYp6S9v/aPmic5kNWccDw492AJhrm7dp2Ya7Aoa6FTR3SCB2CMIpwvUB8hBYCO6BEXNpiKgh
O1v2MSlFuO4LgaWdN815Q400m9In9A0GdM7+n2eiERm4HVZ8PvkO7Eh1BIbqjL0W/cmvdcWy5QW3
d3AnesWtPdWAC+yksYsXCEMC2t7yQwl76KAusweDbgMajXBLPi9KQahRtiD6xd2E47fnO2wJMRhJ
zzqI7C5zdsCSTMqCe9GWmbxJBiNGYjUJ6YpOFcQacAGOc1blIj8F7zsmHqIumcYfQ1HvmzCNq/MR
Ul9Yyq7zK6agZmtBTj2+9C1tWwILVamOAmXPih8XSpLo8//RG31Mnz6u4N+YdMW7j0WPRsACYKTi
EyqmCHGh9YvpKGBzrhx/mLkMecJfJP1tyLS75b6jwYmkv0bLkYP5vu4wwqRf495gSa8wg/qcxf1o
DxQ4AlGdbGt0CYCMF8bwyswQcBYwprl6XM8q7OyJaMXv//YOLFcvaEp2teC4Y2ZI336TCTEAFQHX
A3vvQA+eik+IPIbVkYzJ+cjkNGuQBSTiWeGArPjjq+IA1DEac23Kwhpeljr/D4e2Kealov9IY8lr
/SxY4LhPecIlmD2mZLlEaTK1J7sXxJK9fLp7WYnXQ5Pv8UHOahRRJntXcD06nwp3kYmn6AyeeVQs
Uf/sgF9HHkWVCvXDjjyJG2BeVXpe+F2PyhJjtD5jHYSyFb2Tw3+CKBfEx4yK5EXzFj4rigok9sbD
Bia0B0nJ23EnC3P9oYbBnSmBWzci483VjJRj3qJsLsP35C0o8sZtqfNoCzkfszMrZSn+92ThsqD9
16MENcP5FNvM0HQ3aX6XfGj2TmAw8qbpWh0dc4UQNo3pdFUmeCxcUfmu2Hts5dlvx8pX1Gv4Z2i0
0agxZ7sFvk3LmItvlIL0skipqaa7EYlnsTHBEHk1/7RHl31tTLzY3VeAwQj+AiBFJW9ECxGWaGJq
aEIDqig7W2ZWdITl0bMW8CxcNC0HH2ThS4fuJxGMRCr9ru9NEfImNPAeWc1MM+7dDWVNbBcRBLSl
dwzB+v2jen4yTFx/y4eLzveM8jreTEHDXoNlIuhZbw3Hoo11/r5vNHYjbuRn4k3lNHGpcAEqSZx6
M3kGkZaGnUajkCON0vMUgf0V6orKm5LicLgsRC3DCeVaYNJkfG4g/323bkCxWk4qgTucT/aYyk9v
R+8dPtB5M809xUsWHP9Ok5r56+w99dR4s8pJggrGIFhlG4p2I8qpmKB7nPzNf5fDoWn2yMNcL4vc
EKXmTdFA7Ldr3tKPyIr8zTm19uHbzvRYGv2LYp1GtaENKqp3e5O5K4o2LbjaMr8nmb8tCxU6k/YC
gGSJePzK1K0Du8EiC6yEPGcMKlTP41Q67+QI32/vlVBeWiVaD6eaG5A6lx04nK8No4qJQ/TMDHEg
bIOP4wO75mvr+l2wLRcwq/MQCV0jOI2OtgN3YdeUequnaV/zeH/y7B2wiS6ECBGun4aP/X17R2TI
sUIqNUBdmH9Llbn4Fe9XGdt8ug6SqktOlNfYUsU799uEAgVhURSF3m3Gyu9ea2cHlAJzpTz1GTKz
8hzrO8Wl61MvuKrDfNzSlxSVuH255j+Wk2Gezaqp1fy5Fj3WrX2fM73am36IRzEl7rtFnQBLp+/f
+Yg5QWbo7Vtz0B3bqKptbEOcUOEwHiRRI4Gx5D58Dx2KOUApR2jC+U42LHrihT/PYv+CNoVs4ZCL
WvcWhk2v+zz9Ouf9MkgRRmNTcA6hdIXqBEOGlIqUzggbLC7wZfz1yJwpQ/4PIRJNc6z/4oALEe/X
ra2tTjQZnasnosnRsyHRYL9FcpylwtN6Wo+5wHMm80VyOgjP+lBT442BCGdhQUdeBt78Mr32D1jM
9wsReh4pooHEI0SVTSdVpqFmsgcD8Wh8IYpem7jRjr+4eHFFmCoZTnnRSS3CCRFuHPDanORPPXCN
LsEbWlBpojILoIpm3h3neWt5SoxDEywf6tycDqtOPyGL8tNlL6BN7fgQ0gqlQNsdHW+oiiS+rL3b
ao9jsVuC8VIXOgmzsj/gUq50Rzq/LEboW527fIo1f/dWwJwT+BDMknthiWAVKUkMfzitkqx/pd2b
Kqe+SeqoXKrTQ8DUTLtLOkAnJI9TDvwv1bJtEFKFYvM8D7f6yC6qDj0JAyrXSlB9PW2RbYKyYXKm
lF559YITS1LUwMVH4ZJZOvlZ9IVIm9Il1T2EzkZw450oG1DXoHL8C+CUr1XK1LeXCvtUOeh9kjUL
se8XJxtp8JU1NXqAJYDZqpQcNKXtvabeRVR6uC1TFVammMHN/zIwOQtcLZI6I+VbNJeXDm6MLWqp
/mVXdVfNBdTEvGrhNaki0IpH/E/Siap8wIJywcECMV9wp7Be9lWAd9pfBAfQaI9JIi3oXwdNh4kv
+l3ndDML5TAL0K8lliqI1rVJhxR9SOu5AgbMqQzqS2rcjr9zTSu8Dnw0puhBEKtGmhklJHYd83jw
teDQt1OABi6muT4zXPr2HV+2QPffHbezmLA6jX7OWO19pF3/IxocGHuVMbMJjqkqOyWOUunA55kn
0OKv/LffnG3tqBeYhVH8U9jLUV4BTZbTLtiyxJEd3mJ4YHY9XeCu6kAs/STClJzhLqH7GI4ufw+Z
d8bJOY10gSedFPVzyX36+8vOaheWhYGOtX3ueiMqcq+Cb0QnK0Pf0RVsWbUpLhxh43WSek7Vr5Np
7x89RcwFjFpw0fSxvuAixZlFvjLOTK0hS2PwDRPRXPOhAc+IxDjQnw6WYltWNLiaP9DRGV5HMg1a
5fRdw9JhIT6tmHhbENj04FhqM7vtFIPTcSmVQHVVh+Oh/3+fjSNTfCcCt8caUcbj3BLawCthzwzc
JxT26RUrcgJMUVsQE3T5NY6TJrc9SO42tSS6Gk4YGdfPmMVDXPYAW8aTTpoCBU3sOk4/BqHqGOVY
mqsKjbOeb7AepadNiqMqhW074zFOdTPrS+icyxIBoH+BnIWjpSYXf6OlCE+iyLdzqC0bPHH1YXgL
7b1CTYHPpDVbdmrC9yzrOwkVq3/RP5yd/odCOtHm2lDpQUEgD45bJjkPxLWdIIy1GUvBif3NCsjM
3xIm4A91A28YpWmVZ9cXH4nvlHv7JROykcTC/g94x3xOo/xM4KmYv0fP1ijD8r/DYRwuPL+ur4Co
iWuiemtE0I5g1ZlSfoMmNDNTHGKokXiNBl4BQxwJSdCJwLuRNZ+7LBlPdlmT9nh/JCfzkSXJgVJw
OQO4rHFl1tFI7rJYP/C9JswmZRbQ4jpr7Oav62hRJXpBODHs840a6jdqhgXhegJRXmE0xmE7Yy8/
xlPHNOFXqxoHWO/AlN5hAky7T5bkIaMNqhsBqbxArNRT0vmIpv8WMxUBxe+tEIGba6hh3Klze6x9
PT0Tefhb4rQzaBRTxKlcjF2G4y9vDYLoWubWPf1+zhL0HdsBOsOOdWVHIM8NmnsLcsKChHP/BZQ6
f9e17f50T6c9mhRGex2tfdfOBMZET9/k5rVW8qnROpSTa9PpjnBwlEZGhot2O/aXS/DntIM4RapV
DcstpkGsh6YM4nrUXujf5x2AzJ6LVGTcVv5x4pUF3foRCx7GDXnAvB9XTWlmv03QfiUxBBBspAWK
p+u+N3PFRGVUd01L/4VsFZAL1WOwhPkUjEYc/mnxY/8icROiWagyBk0Le2y6j9k484wLja+j1j9Q
uIuBlcEuwjOGmxhhlYwmqBedIRNBNnR6AgWN7EJk4cee3D1r4nMW9jXCSz9gttBoTBNKoCLhL0KH
eq6PZUl2pyhREXi1bLUP9YnOyX1mXfwE/+wNBcl2gcMjualAI0v0CKf9o/nY2rDWtJaTZb0NwIrp
5E8UuYqHjGtp2piHn5y+vTWw9tF/uti7/UoX5vK9vfWEGYISbG/NVCPZhjDTOxvT+VI7eX55wPYG
ql7U6nwBp4TNgrI/iCcXdVW1v6fJeiyHgEDfSncWlv5JxgKWHRa3BdzUn6JvCK0mQKrFszPLGWrb
gTqARuw1HB/kRngqIptPfppY4gy5uRkWX/rIhI8CNij50U9lglgZth/WSS26sr2icIDAIAHU5AIT
R53ER4lRuctAiXLiX5C3FApboh5cFQFkRe4bkfWHKM4/Aw3ybtxhW/U4OahGo15rq5bewcIZxkEE
rNoFKNiyYN7e5A1n6Amkp9gw+eUwoUI6k1CHpfqEVgrKhDeuTDnkGxMCuMKK649YwdJ4t2IdiV7o
D3oGlJpD4Oe0IOl1/t+3uSOxTzhrrS9HIFHKyKKSdtjvB98473sPOx6TmlUpU4ys6F615SgPF1u4
jfb1nTxF1iDsxkGntFDJviAohtn9A2N1ITWkqwUK/IbxEs0c2vqHFwq3eJrL+cfRmIiH/wwA4STg
ocLPtL/joJ4yP4NiCMQVqqrAi8WXaYeVtTgsnibzUlCut2Grq9yLW5AxyEuRSHZXjM3U0kLB9nqS
Riw3f7oEEQUc4kHGmOAypIZvbOZLUR5F+ccZOPpn8iHaXAr5UsQ5h2DfpY/biT2l29JKCq4RiajX
K7dL3MhB2Rg7EwJxVJn5hYbSbxQsHArvexsLWFHy8yUGD7sPVr7rSh9B4gbcAAwZSowqCcpMgBNG
7JCWo9oG65TovBbJtzpXz+Qj9po5OQprUUKHJLjq5Dh84v7/UZJYNWEkZ8X7GRTfZ/PNP7GLsTAn
iBHeU4fR522HNMe+JyhWP+REpwODrARt5z8/m35KDGpnpGBDsv2/7Lz/IH7w7YSWuBKJ7KIyTSTD
bx33UQEJVsnIqYKO63aPv+1gsejT6gL9GdocBPPJLZlMFLKzhjNGY45OrGSEZd6eXj7y7dS12Gbj
+7orvMMzo8lZj+x+3/WEqBngkEFM0Co7hykxZxPb1UWKPcfQoDYXw9/BLFNDK/pXKoT4Nvoc1Lc6
KJ5TVt46y0P2scqnkVck5v7L63C3UPDu/DP2Qy6HDWLpo63RECYNsKTBMbhTdf5nuK06e3xN0rl3
+goB547Ydf+FKQbST15Ybkyk6Wbxg7jfKQ/X9O5ZzTcw9tRFYGTqUq/uoFyzYRkgBDwuaZ52Mz6H
9Q7DF+UoSH6OBKPh+XacNeDnbWp0gvCxTzNaLPc836etLJnnio5AqS5P6Wb9klGNH29kF4CgJbJp
BXl9MaBliQM+fZe+iOw24rNrQHcYER6L/WyUCuSuWTrloI9A21KmZYtyKdQxTRO79ZfhGHy8wMeR
GFXzN18Get6fT0FEayiI5Zn6Sqa6KolMj2ENeH5YZi1h5ezm21ZXzPr4ze1CjTwGaMmzuk5OJx5o
wXwmMx6JBVYMpozfq+Hqchka8RrVTQQsXl2MGTOIi7aJEvOuHRgcAZjbL+KnujvLeHwwSU/nDB2P
FGssrRmbS+sztYx6Hx36EWuiZe0wsEmK9PU7jU0AZl8JDUuEj/M2kXunbwaO6kVkalD0H9xBh4Z3
RjxviRXvXYEPS/H0G+rbeifxyxOMCiznj8ko8J2WG74kYseEQ/VJuqE9TE886qOvlQwkI+fMbgDg
xp8djvoGnFua8hDoFwWDu6mEqUsgH4MBbM4Knwl0B1aAqZ7M9ypqBggtH5+yLH60FhWrstJdEptH
qlTLwmXiaEP/WQVKfz64vf3e9ddLSGtWf7Rr2XBtUUvByGwhBzHVPdWIhv5qUttwIMQS40Vq9puC
7g0HSpVDk/OVYq0nql/pJTUy62fnXJyeWAvnf1aBL4M9BCE9T0Y9QG3z+cKA2dObuEHPR0n78seV
9oveaXan/Q9BC0aK5CrSJr5vlBfjvazNjXcWRjvoxDRfp08jYrUcGdVOH5zX2REgD3UO+nwDfcgN
Vzg2s1na1sH6r/N0iCPhyrpKwwH69BZGH5q1yd3r/L3nznRx/8MaRWRcYcf6ZtCBta3thGtr1nhA
wX0HdPmIaDpEpUllMGrLdIzZKYiFj0ZISUGv+THlchWSPbqm5Q7UZnh5wPiNReGM1hi74/WmZYsa
rdErjNAlzZK5tzSnsXlOIey6593zwzJ5Xk8WYKtHVh2lgUKXaz6hFwKVNtLowHAfJHnNy2lVD1IT
/oyILzoS8iJdNEDOA+01z/S5xJASqXN4OmFhy88HQEsbYHy7CSZ0FSrMXHvE8Xpo/UhW5IzvaO5t
cSrPe35ZBIL1gcvzj6Paei2oPzHhybs3m/o79KL5mF7o68vxq2m/ZRrFpSUv846h5NRESXDkyO1z
3RktC5lv3D1rM9vbwODI4F+Goy7o+2DIpqE700ActFxO6NiyYGmic7tm0N2gSKMwMETC4y6+K+G9
FFcWyWR8TsuG/0EliDW0HCkLG7/yPBWCOyyZ0fXHqUl2N8+emJ+IQauXLzGXxKIJHzUVu0kmi9w/
wry5wRoMzTeGjJzkLLmaBJmo/mKiCJY4fWhf2sb3KIySTZ1dn1KDcvkRp/6AnDYc+TCs+VW1/6/i
NnyNJCnRn7+0w1dqxddzt0VhL27+IY4QULg3dAwtcAvAym7/WaeWsbwgGBQF0COwUmowma9ZQnbH
fIKD38qL3GEAO1RT3VWTv0fq/Vdj1gpV4gRXCw+F5Xs//EMpDO5GCvl9AdYdQVe03ZjQyLx8eskw
3AqSbYBdHQurax9s9sw8loCHdbNmSINoy03+P1f14gvm0g3itXfoJP8vXlYq53ydOSS5Ow1HhGZq
HhLV/1vNXbaS13KvAyhy7g//rtrzbylxDeIvkh1xQYz1ID4KgDyLAINyyGntcLDLtmwzrAWNg6+O
pysGjQLM8Gk5M+5ec62KJOqyXXewEcdNU53eYYG1r7PjJtgyBaefAfJjOY4ok/FMBAcomn2xgOws
a2pu3GpY/y1gOtSo14eGaS8WGQ3Ncka9bdhT/mvmvn7ES6Q1otGFoHFiK/IbYWPxaSbiCoH3J9mz
zb5zzAzcPOdmGEz7ECkVfVKAhLlzh0g7ILjyyjrVCJbamGNmTqPqqut2z/e3gwZJowvJ8GGPOZVo
1kYKu54a7/kQsFOHelef7aCjxXVBPfHkIHQQWTR5nA+nJPpXpKvmVZ+CUXw3W2s/rCgcS9Cz0/af
1CnoamOdYafu9Ej5aVSkaplRhGY1YT1RigNRx6a2VIUbMMXUJbaZ+eV7cWShpky07+136nR62Ugf
wssMRRX+67NyTG2ryUUL+K+n6oj018WmURwzO8mzUph33dsKlh0e2XCdxkmhPtIoStMdQPMeAWX3
GBY67RA4f2DdrEVheS3AskFFwAXYLP6MQ9Ko0N9ZeehEAQbOLJAs2IBGfDEwDsbyP9nDVyj5fqFw
7zT7xYqwZRUrnQxSDyYDWYGKnl92vZUwusm6XSOeudmFaoCXvO9l7i+75I00YSuD/fuxmngmpya6
GwNulUoCcr4u15Dlo7W0W6MUJMyJ4igBQFAzYR3FbNOr5IckUmmmSkUCFa6MEDWSavyr27attArB
rppYWwjtokJ1gy/1RtEfMLshhww4FsGNu3XrObjBBqoKK5HB8yJfMObsr4oPAWCyJeOIQeYL8pB5
F91NNFxoKybfZY1KUCJeobCkuMg9HjKmCTgyqFVzO1dPwZUe5Zg2o3m+NN3U20RkStPpv3yjre57
suO1C4IwOtfDo7ot0yxowvrEWOAn9QACbVnJweJUnu8wWuUt2SP+QGGp0Xvw7L6wGA5kawoP9RNs
BIb0ZR5WcEe3jDi9hGMctYIfKXhfzreMSQ8QCr7JFRZBHgTeEQCNQOcBQp+qKKEDDpkgCx1UajcF
NxSh5xvyvTVQQlYoNhjFApJzHA3FuUKFrp81LP/q0aM4Cnw6S0WW7oh1hSGka5HDgF66E0YTfRj5
6jNj6K0SAOuyBNnh1RK1wyODflgkyPXwHXeMP+9jL4sG2QIFyhPCn6BsnMJ89itpXQ9w7iZIkAdr
eLTiE0ePjTBS+TmI/GKncZiMqTq4eknunEHqZAlzunhsNp8EWKiI3wCefG1R37If4/o20FrMw5GI
FJzRPBJAY0DOVcGjWIvdAzfg4o+46l7KGdZye3qQroDIBlZj97rSIWZEaxK1eYzy5+wEfcru2J8E
wDcRbKxRR7mqlYLEhNEMvuwtzsXyOGYZWQUQPGtt6omHfph5P5PGy8n9MgvvRZrSKtfH8HV0Sbl3
Pi8R/aFEz9vId4vLCYsNrEJj3aF58ugraVhraFRW3mKY96pIUIC8aarvQwbyu1DfQqs9FVhO1zj+
ylz+yGyoiGrpK5Lox28eJg0xVrj1bBRg6XoTA42ppLhzgOGSv7xPX9rB+JttwuF1bFpptVI8DhKk
PBTQ4n82gl7rDw8vx2GZg6GO1WZJWA97gPzGavfNxEx20XDCHFgY61Xl65zDc+KmHRtm5jRtG5xU
dKfSYw6cf9o9+stdHDLxsc5sJpRKf5hmu8hvHM5MGYXhMg6Oei1Cz0i0L+L0YZIV9XDIwubu8xBn
ycKZTyDfO6k58hihpHLirIM8s/znFlf69fqJmBf+0ooFum6BjX5O0yTVfwxtK8g0auQdUK6k4sfm
2VrVs8UfSSn26iRm+T7XeWX6Ha1VSY/tiN9TkVOKvZwaFJcPXNaLRQcf2Dbz3BS7trqWYDs7SOBv
dWm7MaBZdhLkI/dqp9PPMS4KfIMHIFG5O7zMM4i9Ycv+lJfinWK7PLlCeRQ+uHPUE0TrI0uk+4Zu
+2ROPWstzSW/MAr3e26M76tgmk93EZ8JLq0SAXKBkrX+vgwwlXct0KtplSoZfF0lQo7WLPcGa7Jp
HpPH+4svjmqCVicPVQNouoAmjmYcjXj3ziUClVuVr7d3oGuQZdtbDu1nvi09T9aQPaysLuSCsPlU
49hq7Asm8CLL4bjx4Oy3CKLVkqku90IUmRW8q4QhHaFtc9QRa8SKZpyZiojx7iJAn69BFXlpvFbm
Tba86VNJL4yWZhDqfHQIF62UINZsml+uVwG8W7motx3C7yMuLQ63EjRAV/LV2jsmwKL5Lez28IHf
YBzInFU6C6OowVQpT38brHLfHXzlPr9t5xRR1s2HDiCM/wSfnZvODnmfG7XLpGh+8n7DI15ViaDy
ccfG1wXW3W1magQjqJ7VvMaRVEjKam99XmIZhiBw/Ae/eaWtptJg4lucXHp5TzhO/Eicwn6/Y8bk
i4rLcSRVYhGvirL+fIWvs/jpWlCdgsIr+DiP/r/+008tHodcQ76a71t2RMaP+1u6I4D9K9RFOZ1q
r+FXlCPp2db9V2aeHzXbRJ84CXt0LEPEKRRVkFlZhQDVKuVKGR8wmjT3lEq3DCH9V3wHWxVEmJA2
VryOZQQvyGGwudIiXwLyP2+kZbvESQ0Ti4dAYwqDtsyMo80ZDh1MR9IkVmVipcqpmwoi+iWLbvU5
5xYlaAwcosOsVkU6QpveckX1iFESf0gsmJOgbDKbjd4xGrfJvjt8UXRElITdCFE4+1FARv9GnOcv
WYhX986O+i4JTbXy3XONB8ctALMV4CLcnRXAdKUQ8q3AloHI0SZY1jBWXMG4SWXQZnXYaM7HKwyp
h+WASVtRXNjIfjQ472pvMhqa3vyVlta2W81YY0ZaeuylURiJFVb/+trDv+d9PssnR5hz8xiNPzzP
0fzLwbyTT/ktlzVMDSh7ILdcYFpN2cPVlmkibCJWSafR95OzkjEQsJ4/hcItpnEk/HMFG8cDcWg9
SLwQ5y/p3DdS1UmRfEHnyxO6sDeG3nQSDxQwMF4CCnbnB04DSzKf38diWWNvo3ctGcvr/5u04Ij0
MK0TyVK5zBzid+L8IiLB1K7zZdi9LoIA8C0R3fOwhiyFnB+KK5/SP57GGJbYrmGc5AecK/VHvWXq
3DFBHxGjZo98eO+Hs9W8rfhDCeMAzrYL2FQknz3VVwYb6oqALsy0qUT5Vob1xZQh4b0yEaxyFvwn
JCJBfwbuvetGTVQ2nsLS6xbijks3UhQQQ40vZAx4qtJ4WtKyCNPkqpE4hlqxH001stee/6b1sKUk
ryYhrfLnU8D+HlENHTOGTWNxFT5QtA2y3MIOJxpEZbNHnHYZutEaLSXgM1IGrRy+O5DeTyztq0wX
0jCH0w1rJ20fzzGT1UuQwgXn+M/Mse6yPmIkZKdPnnf17oKPFIS2W12JBYlXJpGAcgTaILQszG3A
DThPsZOQREsBMDVPoO0YmP2opfqZbzdoaS66SXwT15DFrGZfI+sCeFUoNV3OVoZQeOaYUzGPvjsB
3SX9DbiwbjVY1aGErkgTIcDC99XRnzt6I023OcAUIO/uE+0jmQflWQk4X1sUQCE4XnWYHyuDXuBz
FNXab+ndCxGQOVP4oISdA2UeVxCc29uKP1QA+ksdwrF3O8aZlHEuJKxNwvz8DF1xJUDb0SinbdDu
za945h6gCswIdZ9XhjfLkrhHWSOfo+EQApc+oRFVVnlSIMA+9p+gbQCLGxSHTiEvJsbEZjuxoyUT
sj6WxCMnjXU7Vg8TS1crfpmxtyi16CAD3u8wDCdQeY7BWdlIvcU00akW/o5xY2QP1adt7e6hmwpC
W2mNS6s5xFygm7WhWxDGWQ45fFhdNWYhpQSQ4+G/DeIgR9Vq3cRFykMmA+AO3T6GxyRb48TzoOgw
1s78SQB+6nQimhVA8xyCQcniPyuAeKTnooRbATdrKpN1Mr5DwXTQGUJbuhk1Y00ChyDmwwsyhpUc
29G/o9Y5cTcvsg7E3vj1MUoiORXPAZRL8k16tRBGMfuEq501FGp7ZBU0Oxg2iZyt3TBL1yeBjxp+
EVToG3IgVd1c643JOKtUzeDhyqHsqRMTCSLp+OeCHskuzt3z8/TCiqtn9puW8L4SR+SAb4rqCNTW
cCpvZlOVrHChf2pdvqc3b9WoeTpPu6++1egJWKr2ROmoNv3+h5UHrn9djCK11E9vM+325BjnkSuK
P+wISd86Rj3VflryU/59MFmDleHus46jXIBNWEsuNZO4CoFR/i23NIOsQujV0t8l0wAIIx3wz9/v
sCutQnTAmJwU5EfYVeCGfrhRsgOrc+BuN34BEqqVfy33jXE06E2na6UDkN/ID8jXDoN4p8kueB3T
XMuQmZmOZHiT/vDSfSQLfSncv45C4XjFFGIgD0SxPL8T5FbHhOMawhAG6hNpPFqC63uriYXVrSG8
X/oBFInIARLkU5UrbZT7BaZrmvG2KjIVHBj34ib4/pD/5m/yxCxZlCbiYkFBUESQG+nx0ev8vzyQ
PbfuPthXquotdeHX58a8g1MJ+07+WfC8T8cJhDjTujwyLGkXnZi0j99GE1//Pekm8q6R1f50p74T
rF9YaKRp8JKUT0xXyx2h0QyBpqKf0pqm3tsIGQ7qRqDReIA1x+Ix/1QjvOon9Ic/jZY+Exvmr7mW
S7GHhAz30E+oBfRau7moQjuVyhrUW/wO8Ust1rCf8hAme1rVtmMdXb9YAqrmn6X5sGOYQUbbuTb4
NBsvB6IfKrrXYiCuaqnhrKMQFMGu3o2xr9ZxJZGQasIg2Tw6kiI3Zv97K5Vo2vkmze3gdai2DE5z
sAsVSo/nPqOapBudDYEOIUVergE8UX8Ow/0u/pQT2OWU1iFCGEk4EiQdDptqY/0kT0GyKE/XSQUE
I4MNSSAWl3vOe1njxxpFE6BabzTu354jStK3+kRtazkomFcQnT0VqARLPlc5yxuF4QAUIKMSM9/R
QJt1FadZGHWI90z8gDrnr6uHTiRLrkHD+Z4Ovc8lBtWy8d2bzyk6QTRgsp3/uaLZkzJm5IGRK9Sf
Ov3dBIP2ShVgpim99hKodfJShEcY5PpkjEUv9+p1I4nVDP2T3KWR2NTPaxinwfO/TbwcV8UEThRc
qUU64bE9r77CAiWz9dvnAAnW2FWXVMK2Su5H9bayr120OReS6dQLyCLM3afufCcRh0178WUZMBFi
67nZOCwVWzGceY6YTSoF3bQwu7kx8xOO8ovBWLtHzgaZWhywtUdybD/81RnGfZwQqYFXtq9NFxdR
vw3MCBbiRBbs8d4wf0BqwHqkJxN8X9sCEWCtWYDmSpvcf7J6rJQ3ev/k8bEbU81cRjpyb8SrFsJ+
rgZDfgPJT6mEMsq2jKeIU0avBfpRog01LYPCh6qM6MHORM+Pfhi1nHPzEhY6RoNQyBVw5cKvP/QQ
KAzRCwPs6ffr5SBbyJgMd85ZArpH4TfA1Mg8VBoMPvOp0qRHgK7PXlJ+3X+px996Wbbo+jS7+J0+
fiNA+AIqxfIOXRtcZIsDA2QdvkXGbYdtUb7aMAq1460pHJEKOyQGd7kFyw+sEy6c7ClwUltpGxg/
AoczfpMc9vEtHSOJfPuBNMHFlu+DYG+Xzm26NfkgA2enYr164KZcjk5tLm4FgSKoeKbn0zBHu+Np
AcCiiAhB0MCULA470oh6Wz2Xujapsms57cDMmNGWuhQGbhrqGqAC/5IGzA5DHlJst6U0EtiJo7Ew
xrImGKeb0eD6APr/tRb8qxLBIUMMVSKeFq2wJ3wt44XElUeqzQ9nEZxaLzY6IxfEPgi9oq8AcA/A
0ydtF/7/E0HmbXTf4skdXPybebKkYMukhQCHXQ75x2Q9rFTdnlcD8TtmdHjjKsVi9QI2b5prHLP4
BIA9R+uv9YwisUSYqKNhbFLMOimE7l6tcmu87gFno7QftoAq8KQKASn4jzqN6V5RrBQL/bZErwEQ
F9P6XGAFp/nl3RT8vn3yCs7R9STSMMkQNElC/temlrOUu2YZAZ4RjB8rXvxJyfYVw+49ab4R98/R
9+QP5Zn8paNa04/AYCdubeDclnFt7dENnUPl4kC5E1bKA7vJgRrM6rt597hq/dbbUIV+jX/rRx9V
1zY8Y+AiVT7d+rm6hu+ce5QSNCmYuR9TnGfs+NUWB4Z5wlq3V+1r1COlkfzyVxhqg6kWoBt2vNwG
79lHrN8qMKfnd00FGgVAJwi0sELp0bkqA1m29BvxvRe7HEECg8UmWMkyZCqBIdUYWQz4c0YWzFwu
q9+JH23pZeeejcZP1ABrW35vR0TtQXt6TblaagDXHsS/23AQloFcU7GoKQrHxQALLc0XYPUygAoc
7abuzwXVJ3ZMEqXRnc9hNWGkb1476mstEDp0z6xxXQvYqlhjSxsaGC8fp2Qfs90xeoQScABRYia4
1vAZO+uB0aYNHAPbZX7NvHc8cSp/BpF2Ig5W4Sr53onHhp5brb22jik6TewyM43XmfN7L3m8sghn
s2P+QQhNQF9hEp2YODWfOFwKhzatPfQ5+ssgFPX+caAMwVCd0PT4wJ2MP2u2yG112v7bjDG/AdOd
Ptazshe8xnRl1NdDofbLLsOxSDX4ZZHmrBUs97jg0dTZFIagHEE6DoGCtPgc6T0lC+zhUVxo3V9f
jPTlt4o9b9JTh+ydCkskucR8/G2xYab+V3BPiL9hN8ypL9UANnq8e3g3fy2kFwtb7lc7sPz6WXt5
OZCZmnr3+OoAPNLz2sNvbPEBQntf+WOGuu0vDJ6btuP6pkG9OmkgDkFVqHYjxxX2WWoFLprEv5Q2
cRsr5g6V8iqUbodhvMT9nOZtWGfNb5hnOT0WOlOGDYGLXTISV+T1vYaahq/0pXP68whxVwkPUqrg
hDmtEKdcFDDoXJ6aIs+fUc5OFTMHb32kcvdIfrpxAazhbfUDRHWW+If6twK0txVd8P7IRV1GhCN4
eRgKcy2eF0tuustmRp61nuh4rFQ2jqui3OCeJ4k7xkdZbJ+hkEb/yIfiSH26mzOkq+VllGodR1sA
Wr1xbLZEVQRPvXnW8Oq/CWlA4vm8pgam269rMpjCZIM5D3H0ieWrH91ruAqpZNAvp5YZaxeAZ7MO
2BLxtuRHjSzme7/HqRFqwtRV0kisDzJncoVVtEDGtiw08PdsxQW53C7PWwQuQd81KwLy8KBcFZvq
w8lhA7Tf9LTv4ZBxEfgTtOKPbAZ6VMHjBUZylF9TtXG5OqrTHSVuMnip+5Vy1M6P9dOx3YMsEuhi
MGxiF4iZ8E+T5VN0zwu1dOiln/l0h9cPlCMXpvGkjMjprWwtXOG/7dViNpEXpu/V5bKoqM/zw86+
euyxRscDcF0oPGrnEoKYQv+xCitmCoIJmWMCkDxtY0pthwCCpm7hwouvEOKMgPOssYr9tT1fujVM
Z6hlsWn+afqixtCY/xTIO3Ttqqbxe1M1VP2sYur1wXzSqUKvFY0n0xt3UTRzMSI+VL+molGzRtAF
8aeDnbhzcFCTPcFQf/xrtamN5SbaZjegic2cQQzPDdLknOLKcHCsh6mJPPj+O8JKaM+3JWA/ic+4
/yx2t1fAU1hUIHv/thgEy2r8pVeqOfM0bau8tIAxpzEeg7vJbBmzOS7QYNdXN/s4EQhRRRS9F1em
uDnryT/5FV9pJr3SKPtdkBvrjnp3sp0SQW8HrWIdVlFDZItvwpt7gG6mlqtZLmVR91DPLisFqhQJ
fLNCgaTZY9n5ZVkEQNErZxkkV2ENqrbNQyDfSWhOLJw5GmaJMd8bhIjfH1Vy24Qt7yNS+UoBC0nP
ObhokBolz/D/3oDMgsnGApgCS0qDljeAJ1JFpsZqkAeJ2fhNXdZkkGcJHUwI/QJmbUDppb/yPELe
DGtKsKCcMXMYwWDfKmpPllJFiWIsYkmHuEMB/w2jXjRt88JpFLBKRNEbuE8auVlyTYOUMn0XeYlv
ahhKMxuqk/28TFCqrKI+9QeCGXrhc/obMQZr9DlIy37cHcq7yPQJd2iWQE0T94AVDjxLUe0LlowK
H4BiQcAhLEYhLQQg56OfjeKpBzzd6QKdxFp0al4+zmLlNUrS0gmftsJ89wjCDsvGonhjAE6snC8K
+4P1W5cTe5KFgEJrdc86Aej/M0MTVZpgnI6NiBtABlYMd2laqjEfg2pvshWypAwbhWpU0B5HIcz/
+Tw7e8T81VJ1PDR8xnK1qvcNzz/hQ3+T1TJnpl1sh1vuqbKKRkHVAo5+W4gBuSXAn8y+bMUnmM+c
5Dtm2DFmPvDT+NM+gxoNmrHQAAr/mZLgCDEIHdBmuT8PyVih0FJXaTSLhnTQ/ZXM4YneHDU1YGkD
5It0XQYATtNmALSWmPbjyLUu8xHIAG9iLvdSTMCJX2irw8HQ1KEl+8cb2J1Jl3m2/WfYC5A2Ji8M
xgmfJ2fZGpd8YlfWwtCOyEsiRVkV5kcpj3Jxztf2fpNOMOcBSh6haFmDj8/uLDdceJoI2MQel5Xt
ceZT+v8PuXOKQc2vIXo7Q+4Ke7uHcm30eQCd5Z9yllhi5Pw5phkPrxoYR3b/TUiBwmJ7nPBMfHpJ
vayODB5Er8gaKx9wEqDr9R+ps9DZbkYGhzCIE94yMM4XoOwbibgTp39Jd29EzMR5QcSDbOh2knm0
lH+qWVQeDlolnBTL7F5JWhVLvbJZd7OnTNG+Ksh7YdRcPuP1ehMSA+bqh5mQyZ7sbxyaZIjiQa4j
TTrHE/LI/6t5u4aJYAzf+Pg14rwAE92G4kEnsjCaIPYzGXORTsvJkgj/qqSedduTzF6p6QVF9Yz7
Kp6abjlaMvLlcE83NviwCTpzZ53TLqnfEfMDrYL1ccXIv35ak4cI4KKKxIBI+9/+eZq5EUzVv0ro
E/SW7FDjRJHkqVkKiiLpJAlEq9WUnKVMoFDhWeba9fQZzNZHBrbuqsASgascyPXoehfVzvRHox8u
nQE/U9IdJC/xIVekiKjwDZdqCVKenDNNyoGGsXmG5YpwDHZy1l29TRJTPnuLo5aP/IdW6RecdKIZ
TeIAjtODkhVCP5t27Z+ADXS1bF03vmj7yCFmadIAkz6Mg6MsVdRMDIVYxdDMtnY0QDOFXbFztBYd
zJe9fI4ngQ21X8hVW3PCyb749yuIe0E0dX1x5nkVmNfN+l1YxoH0QIgQNFaUKK2gzGnxvMwUnGm5
wRIHfpnb5BmyjPLOCpxbZ7zlb241L9LUwi/3j8d4hXGZild4/5uuRbO2rMrmBq8rITED+O50xAyw
YTYTRZ9KVx6QpO+K2Q0H4yGC0xLkR4UepDIbPzb4WhDumL5D3/CwS9/CmzD3XfOVzwyElzE+8cN0
N2rqfKPBfCdtptbWzeRKzJ2AfiOYUuHiHYWfznN8X4/gtyDK8fNp9DYrFVPsggdZc+4FrgNQLdV5
mbfSmNz6fEyVOCc/O/zZkZ6uyQHi+VmaudXO+0c630QcMCT4petvdG8FLLMEcFlXTvwiRJTJII7T
ZPckrv00rI2Xw5pdBYNxQw1RG1mUhyp2u7nPUtKGMLuA82eVzW7B7tQ13OBmGla6Wa1y9lGqFeHD
kJgKSpwpAu6obwj1e2bp7EMozbGd90Is3iqzyOw+PbM+ri0djXdEuT0ZBBGsAXHWhy08XvXVG3hm
yFZPPgDUN1HnASXIWMxx7U3ISjriwfIXGeUnh+U0a0FZYbRuL6erQxjGnVM1DD0soYeS/xmeHXui
JSzVUHhMRNkNkrcxi2JSg0AquegXvfWqkCWPN2IPeDN4jO02YfE7OcojhV88scgtLWF86g9PJSbt
G8Tex9wBat74qAdGtHNlTn4iJpB99XH1QueCHqfGwOC2PDycuajIhMqnIoLg6uJYT8nHgS1XnN09
LkftOLzi2JusyV3EW1DzgmQZfCNnadQLuVgv0iX5jtowmXrM68sTfrVHxVONIT1xX4EZJkhhBMK5
eQkvrSIBsojdrBq9xudoBA32bph2/Zn0B3E1PKgV875YNo87p6MbXRk9pe6aMU/mwjJDsr/fc+V8
GJmv8bdTqcaW1THebOu0JictNC9rL80hxKmhxlu0KQgi3gn90gQEE+VMs5V2VaaOXMH4GJ0BNKG+
hiMaoqA+6rNNRg3BbQSkVWvfAvbzs++iia2psXi3zTMsXqr+u67TXAIF0D53ecaV+R7hRv3jHVS2
JCZfPIwjKXsq9KdEeRP/672eH/fJzcd0qcnsjauWz2ttKwtgJNNgZ5jeooqBMHHnj9lcT+uxW4zo
Y2ROcYcSrPOAljjBgXT7G+ecSBO3oCzPCIWUTyGaY/RfM5J5iqwXx+DdbIfSuzz3H8nTPazPU0IC
csq+MpGToO/5m73Ys8/eK6cvqnCIH0j0Hb1Q2ZJ1fwkDW0lwXcGgKobY+45L0pZDIlYdEHNv9F5c
yaTXGshXHIvhxr98FO8jGd1ZD/xBmvb3DorgXah3o5f81SryCnXDSQDMG4emaY+brNUiy3CtfyQJ
mXTeKSX9fYNiOIoLFd1p5Kxf1/52CrbP3GMt3+CQt4LtF4feLLXWwKwbjA7LYD8m4mbYCVeGM7/F
lgY7G7G4YqeASJr7rEuAUiv+HRBLt22uqkGcM81uQX4vQLP4RmImgWkD9EmuzvhLNeRO4onzee9E
9I0u2hhY8sFfaLeBOKAh2TyMbZmQIm5awQtBzbgltTrILH+A0rhPJ7M1O+/9B31tDLkHz4bdVbis
0btUCgp7tpAjLQ2ai7bAjeDZuGVqOBH14C2Vu8326FtQnuV1KA/AKmdH0f1lXpzWk52mJBnlP+96
1i+PI+MFyG1SR5+huLGaDTU2mai43/QOrv3B4c39WcBNHFgdbcDO/d1QHxV83A0M6kxEnkZFwe0D
4Gp/A5bqe978n0zjs89d0GYoMwmFBlXTKc5TKNwT2H6x4aXhTLD+69yfMcmMEByvu/6TyY7SAPPn
Tt5zOQyP+KzayWKnuyBGB8KMET9SLbn7n5Qh9dP/XFzvNoHULAYEzaUNyudRMO1ouyqfOL5eRFiD
hDpVFqrqtbk9KY61ikpbgbH9Bl/TC2YHHhRTlQyVIi4D/rzTh6/X2R0C3iJHGya6GjH2rYV6j7+d
G7CP+IjZKb0GmFJcB1HKyBKYV9AfJIk91V0DZxz4VJDVrz7AmOyXGpCRLCln4Xzsr7w8PdyMcras
O8IIuW7fa7vplIym+jfD/SQDX6N6E98WiRoGGikFAAKd/T13U3ON13LrGTKzuN8NPJDLDqDDcAML
F7imlH3YUHhE2z7GtaO9V7wOPIlc4ZJRYri1D30IVfyWjxHKpFW2XbkDAyTxc28BAVsLUtsUeVpQ
c45C5Lvnq93JqHxXE/Dmefeni+AJrqorAVLFMuSbpybYM6naON5uxgqm23CWDwMaeTTIme4XJF1k
Vioad1/bkZd/N0CHMpnK2v6wZjJJOwl3aA9mSVNbys0uBAcZ4B/+x46WsbKbYH4iRYK3U4pMSN3O
EEr0dDDEJlEqRWXmuqCZmv2/Kyyyy7d3Df5AsBzCOy/I6q7qJVMupmaHTw9gtud7Ed3BNmQQ51Dm
H2p705zY6F/MxhiGfxK3+wImk4HUgrnSyqXR64NzHydJAj6sNPzVVrPkWrVphdt2PiZdG1QShpE0
/SYJIHALFnC+Cv+/Qm+cEK3W2U/NQs/7ZR/UcsGsHAtIVRznix0kThCaCCZl/oBKL8Nkvb2AJ6WH
VV8TQq2s7530sYpgnLOtTBUwcrin7cxLxVdkv/whCByJOnvDE23ispSmzTsny1c6tFczsUcFaCeS
JY6veY5tB23x9ME4mKEtV5PfcqNyxa4JGQZgDpZ1j3mutVG4wms5vrKOrNkzIzPQ7y7Q+G5kuo0K
weN+A17gE31a258d+zN+pzzANoLR1RwB0G2pvZ86/jn6BrhmOKn/JSHaJiZwsPM9Clw5+JDRg0TK
aeEqIKjogeuxmfAZVICCcJA8scvdbIfG5UsKpM1W2Ax7II4MHZ0LEaCQesGVbocYE3oxLROtQfKc
Dpfpg39HzPVWyC6CsZ/nB2sJW+62JzyH87aZTMqlWsuBzRcRMYJ3egPc2+K84PBLp87s2VtzvvPH
h0RkB9jA8PYzq+fb33iCfhqSoqexh4LKOJCIpl1oVdjyHOHdATUE4tm69ATOdskhNz9ociBfO3oD
Qp8WJ54uwREcKW36De+ESoCfg2QzPMYT3dxGkOMwULHktQjPsoBCVkXrcjdRYg+ujJK06468sooP
uatw+gnuMKe2Lgbw5b/CNG6PND34Z8OoxQvyScXlHvSQmbREbNZ/E3DrFsVCXTHpIk32wZi0n3Ap
mAwXUzXNX/R4mvxVTRJ6NgfrbMHQ+KJlQxaIGSrDMmbR5J2tkZw3Jn3qlw4hDnLocdG5VHCJ0ba2
veIgRP+vOco7/9hpipDOVrW2z2IFictD8DUEe8PkPoT4i4H17fOQS7jNbJtloGnd60tcfBrzC1Vi
dMfO6mBmxjqR+Yn72pQ50gFm40epbRmzUCKY3BNLqWxKAbFZYSmmhAxbAIatZdMzdeIjvvK8HrOt
/8uLeLDr9x8VlIqwbojlxgamCOJNmS33KvOTelA7WTY0mhQmcY34QiS5aEzxdeB7FlKs9y3hgO8i
Bv28Okf3+pkHcSwJr2yzM0FDqiJgkBrnjEAtGNHfZwBFnbnVK+CIcFxdrcV4FpJ8VmKUlMcFqkDG
SltJMZLrpr9gVnWy+NUwYaImVDuHT4XOdKgc2iIZy6sgnbBGUx6DneUC4yo1aQxRrkxdFEw24Nd5
inmyuw2QrhwjhdVFNj2mitwr5bQghhCuGpsddrDnEmq6Une4iUHLNFGhmhEksPw0Aydlm39859d5
OTUsKkxLAcy1tnQmPah4uzmo/8wii3OivGMXUAabgVUrH3CffRS2S4tpvwBkTmOPhnZ6z1y2BM0T
XzXsRjQ9zRRfPIjwrS986I0oxVhYzHsQym0NSQfVS0XwHea21pF3cY8SG3XX9JdHxmoMwKjJd6Vq
dhDV28LU2/iZKQ+GZ9FSt+Ojokd/Gx57O5o0MDC9itDfsK7iAEK69Qpqbl6GuXvS2A9O2HaSzhrU
j8J6rnYqQ85l0dN+0NzvWjGvMAhNCFTJQj914tDE10anvW92fXJv//Gbhyxr62KayCBIeCF+9QA6
wWDzwuGHjQguGWBChsK3GZCKg/5U4DY/w2OIKIanQ2VbTPm6SRyGKmkuzrQDi5RIwsKNrkd8UD68
yzLv2tQVuwXqKiRYVX47g7fFr+DN7oP6s/PtJlFS+OwunTrHynExk5Efme/6jxh5bFf6wdQAcaCV
+hcV2OtXPbdbPWXbEmT2Tm6yz+t5Ic+altFVLgq23I9j1Bd2jefl32PXj/pNoJiWG2AYCsyYlKnh
CN9mJAaXR42xUV7WVIRoGdLkxnxcJpxapmRUXfl+y9oB/qRqxySHSQ5DDOtoZNK24svlq73kGeV3
b36SLamskeUsSNMqNa7+sMg5nulKs5AUoC3k4xhowJnqMY1RKiBVh2iq0vq4Hj+KKpFFPDaems4I
jEEqOXuRlUnENrLNqmkhMX93MgGGw6FIvfayqnPKBXebrHAM4EVlNZ69p57nvWyWE6Qd9QFjz6hq
YXB0bjNrRrOOIcVIcz4Sbfs3mldghta72ozuGNr9h97c4J+UEYHcTRmHoMp4KXM9YrWoyMQElVP3
8v21k26sCdbLXn+XX8tLbl+TCBemcbJpygNo1Rkf2gY5Dv7nLWaUzxVqOKGifV58BdTwLahHgoSG
8bY1XfWQW7VeAGYzxXxPoNKyT+8ApJr3kj7/AfI+fzOBFOT7glzxbh80Yx416M6EIJ8E1fEB2pmw
EXq5vCZABhqmkp24LhE4WzcpyrDoUSOwv6Qw6N4WZWri8ICTn2hge0zjdQlRIqyH0isiYcy2uHMq
420CvRYE59HkO3EMminJh4ll7QsFoFLHKNLtfl9MixtE2DWQWyN4lrVR+BA0gZJPuYqIi8vBZ7yQ
T9oryLfxhHmZjSIkyLgyBf5TFkD1mvCkP4oB0QQXcIOK+dNWY2B8xwXPU7DeX0UW9B/0utzAokUF
C3A6QQJed8q1MWGdF6iPFzG9oxOR3TlNRUXb5qDyYlcMBcLAKepn3Nyu78qQo+yGzU2vYkG/alE/
z0mq5GZxlMSUbLaCqHEYVysE0K+fyNrXZ4v19tql+KdYkDRfwVMvT1/Zx/17Qf7UwuUYjfPKIVU6
r5RmqyR6U5umuWc+jyGteErlr5vwT8znCnaft9yTaoiCYia1apntEMOxhHmxm9OGGVwQlT6zM669
x/vUFQH2B3hPK5NembNL0ZFsaFxnih4ZyoFwNjRnvqP7lTI3o2+GU/7lRA7EFx40klOJ6Zklj+a/
JZaLJwsvwuInE8qph5O+4uc5TyZFHjtmOOqraAtdNCP8sOPrO1VJtrlZEHHxlxuQE/ibs8iZeHmJ
nt9VMpyGAWUtVi7eJbL+Xx7/ScloXY2EUmPKrwCUgWu8sOLJrPGYXT5Zs/upfEThx3gQgxEiQ85d
vDR0ygW+3a2Mg3aPFixtUrDTrg5XhcLoqJp/J6GS8NCDhOAKFLQCHcxP4b+Pm3nl2jlV9ApCU22f
CtAi7NGuDb/DCLe2Cv4pNs/INKGVxGOZB1tt5Sp92GIUZzQG+Gbg3DEZYuVE9IQHXu8n/QovTFAE
3fjrl29OHXLT7JDHBiBnT3c2/YQ7zokw2xBqzip3jQSSplLekK0kvyt5mU39IQuJw3hmPSyJavdu
GGss2O4oUu3doLxRUnL1L8+GcNVm3SYnE9J5/TC7x/xsbIlyYex7yUqnlBVigcrJsAebqq221XEp
vklSH32tFuIHus61mHi7plVnXBUb/AGWrTuNoIMfZLlEHBbFAW0dBktJ4v+T0nhs8SumfZ1TlWty
uD50bqOFB5hte1VLFJXm7YBfKvfe0FPPKXsuo33oeEcYFXWQUOfCka6sCMbYY1I0Hx69CAdVPey+
N+lk/bfvzOqfAK4x3FiERERX/ZJh5q7EzdYD1VQfGdZickidvTq1fZTLCze/WCBN+XdwnO7s76qG
a4rtteCuJAOybqEgZPIpACFNvPSwlerC344G3bUxFiAwtqihLy3aSlZ9JTgjEEKf2EmL43WcIGl6
akw7fmPB8sl6LC9z1ecrzvnNQ8Pwz4dcWHmq5Zn64ft6Pxq5NsL+jnet5ZsMx+dCfjUkiGwcmsFY
GsKX7tP5MMzKb1o9JEGdeOgQS1/nexgbPPSLIUySLwimL6SC7ynW2QJEcQLqhUjtATfGpx9QwFr0
zOCQGWlcyik8uhvHeiSBG682VYqD5/njnlcBbCYvd596R/uowBgWyMlKzB2kXzr9lXJN0Ap4F64U
tLbhDkeY5f+qxxylAajn3N8dkEB6ET6mG375n5OsjizJV8dP/kZmYbK/+rCNYTXPaf4aw9R/dssN
GEJkwiQ24OCF0fXN4M+nyqk7Gg/RwGe0NZnUIkrWA+QxG0pSx3dmG1t9Gl2pqSVNFkqu9FrJzfNN
aEObN6RBsNyuwflmiuH8VWnGE4iUQcjLXSC+/pXd68WTFqw7VkXqbOgJPJXIIP2j4kjvqedKK5tQ
dSE8wztLfwSbrjfk3EZBngICFFtY+MwdS8nR2F278W4oL/0QUYZwhSOCy2z4SXDIseRS3v3+Y9TW
afPJFVEc6UMkNykPDZKjJyoYU77hJ7GCDrsAye78SdBvTc0Ch9Etj1liPjYygXecPdtKHF8B3kEb
xjwMF1ZNQtnJLtryrhVBcBSh1oo/4V0+qe5bMAkoVCegENbbwNFYn9lVH2EMbS3crl4r5ogsB11J
F4MaadC3xGCU2v1cofNwgrmq+CatHxJcUWHbDUnlCZwPgVtYN74iuchwR9UeW7gm4M8YSxnJKaqM
6Q/Hsffi5JdSq1ao83fix9TI5VnfY7zy+YZm/IVQmQttU8xZNhtPPfcBqfoH5bR/O0tAKsFfOw5F
SG2REcqFRSzj0oLbo3O6zffsN5hanwm6ysCDjFdPZdEjkP0inNGjKARRjleYE4QdUK8+LcWUwDeE
9Czx9HTfLf2XxuGSzzBZlqJHgECrZ4Riwrkje7rKlycdGkQYrssxvBKFVJKhedwHXJlr+GUwdo3h
TKViV5Fb5FFvJufIA1O/cbERive9gBAF9tWEnYjQDhqLz7cir2z1tzoKjV1sXgUnu9d0oo6SpaGn
o79etPZPHK3koavl35FRYDjUic2sijPjKSapHnqzwofBNXjALVdsDuTJtWFW1eBLhVLNG/TywX8P
2kE5Qbmx966aaF30hCphNiUcfmLfmzIQVpJSCWc048ZT9yKr4U8A5tBtL0lHPx33TH1G30pcswsO
CuOrKDoiYW2Je//i01iEuKTQ6QaIAhIqSa/fPTIGBpAecvmf/PnVFpVIHidUN7fPrc7GCxHv6Upd
VB3upPmIwxIWZRw+VhGMHlQYcRASJuxEhj4Z6J+mFyhbKhIFj0Zh7DltrXVEWuRXbeafI/M/TGLT
+335x/pHw+E4bk2VOIk+2y+TPAj2jeQvMVVszDD8X25hMmIjeWLnjuPNofy2BRk1NbDXKW7JMeXz
HEYC2YSr67vu1sJr4kJsMj/uFTSbRv31GOzPSFum+mxPPahVHd5F8xTtHwdf+MJtaZgOQEDf+pvo
/mKv4iNgzS2h3EjBiHXsxCiWDvGcVxKmPGDRuPfiIW/LlZe+zHJrFDKWKhrhnrUGQSuU1y9z4cwd
cMPSap3SoOLHZpmrnR4aP0W2zvutZ9RutMuLjaGJq48oSft0zYgLO+R3Rt0kOWaWLRk60ZuMuuku
qGgjsJn2Iz4uq8i2i52iooJHNh7JDTMhlSuN6n0aCCTdwD8HGk0a1g4vITZSXwBMVboEmp4uFBXm
RGJx0jIX5R5vIA6OoTp5O+eTc0a1qJCbGXXNN/LZHWWyIoA0/SLc6byaykvq/orwSZnHggKhS76t
yrL6763R0+tyyfSrpehyd/LfOW8l/h/chDlvHLg84aYQwXOnTVpVFVAFPEuxrdBxJ+IGMfXiOTp9
n4LaFtqWBYReoDqrOLYXDOZ5y6hGuqDtnl5ofzHvlujIrVxQ4RwruEB9cZ0HuhFkyt9fwWWqvJfr
VDp63esXXjPVNHgnVm/nmz/FjOwJQT8ooH+NrgpidImV+0V4YdKEYQjM22G+X6WiWaqBq2sTD4xq
VDsI/Td2aTrwvrqV2f/0+54i+/7HabeYe51de3n3/0rP0e20DtFPu3w8DlqGT4B8OUvnzb5kuWyb
Ub5b81nVKTbYJqPv5B95mcTFndzNctRfJeb7TRM/CUiEWQM0g2yQ6BxdLd9UhRCe/z5qhP6ggU0e
sXw5+g4rHuR7B3NYBIJKzrxEfrjBfHgbirgfu0FPuUaQYOVI2qv2QiExS1HkMctTBPdwneErcRC4
bej6/P5qgQEaJ5MJVadBrSP3L6lTPiD9o/VIBeM3hGpWm5HIWOduymg7s7E+Y1PQeQhewna7hI7d
ZR9dRmbUtFkUyf+wGfmAzFSiyp8GqGA26tLCgsAAvzisdrYQEMU54tmZ+KS4jwdVkncKB3iTsuN2
Ch6PDpTk8agziX1aVZ+w7dwEbvSyMMPk/PW66CN9OSYjAh3Zx6Y6CqKiLaxWrdVBk73UZS43EE8J
kLRuaV4aPtXCdCokTa/8kzagBZ5HQ/lIgbxz2OADLncmkAs5571bwCBEK80MwK/GBoMlLTZRvRwO
Nx5xpbqZS/9hiZyiR0M1byF8jmEIrx4Eq9mg/xcvDqS3esHiWa2pjaVfG8wv1idMm5qNLvljzWo8
UbB631BtQ/XPCxqk9PsQYJkl6M5ziKItj6fc/3DFk2RGaHqhnLkJlvzict5tmY1ZeQG1oTVwIAxg
hyZlTb7CQubWSqO7phQgiZX4DNNavWwgy4FED6pM4mPQKSEgbxBjrImxiSRWgeddZYkGwkqOOvWx
m012YDqH9JXyWJL8pKEoO5QoflVzbaT+Njv0NI/RNv1xLk8LIIiDYBPluRBxElwH6WF2Zol6kTi8
OYi4rx+C37IS0/1sCpb6b2LVKjeIZzZK3bKooNJ6/whFuaKudqXsXdt3hbRrUd2MjhLYAUUuBvI7
lT+HRypsZFt9SurBDeuhkVno7emctJu1fXI+TMa3DsxVB7eJ3IZYMeIy0uJOLzV0Tr4CWVGzJWxe
C8GMuEWCn6wbavpA+JjV7ohb4UqdZIYIl6KRpcDWOWkO9mHcGjeoUzLf6JxODdKXCrNG7DVXLRfq
ihn2LxMSLdh3IOdpY7m6BWN3vj0K6AV18mIZ+7ZzO3deiYHaYRYjPfZEJ9iIPQ9lo46DVUSTbTuf
SZ5VWPQ/+vY+rkhD2ZD7fxaBOYyrWc0zfdl5IQQ1JIO2JNcvXHA9f7Pst6RPNE78dJ+3225dqzYy
6Y/Ajv1QBx6mwQ6QogkMnSmXNiMFom3jZt80jM93s5lI91288hCSQVWtvjud+bF07oNbWKi+GmPC
V5UKK6E4JibdjetZa0ixap1nfgPB5olaRoc8ZR1ZjrWlmROlt532Y9XV/EobvVzZjv9mol91q/Ee
ezm9gvI142qUc9VuiDAMXgcuYsSNz8s1qY59Biu7hTgUN8fTkiejCklFQTxO5hi0P4T/d+h6zTlV
fzWWpGAWNoebs/Ii79gEM99246T9uRN4VRbSggNZaSDHQTBXBlBRwoQ1jbc+69QStyBb1ILibnR9
4IPKMvKTq2GezyuDYJ/Kxb5g9UxK4F1wE+Y85AIjzvIEtW8g6YOG8Nk/CB2KF7oRM3DvTCVO0SVi
Ua2hCqcAar9WgchefSnbKP7XCtsEUoJ23HjEOm2aKA/C02yhLTOw1Edcfe4cn9Wt++PE94UNu1GD
41yK83qFsE0pO/w4Ei824MB9F1OF8QPe6rj4EEraG1QazdmncR4WIee/YcXPhrbg5X35VKz7HoWy
nOCz0F5aQRpcpY927WIXledHMngt5DYV3B3TQQ7qkm+mNrL9S477P5GQG20xaRuuO3awfvo0B1qf
GH8tlYCtgWx3oP0bULCXXVzuafUm0W3LohGn8mdh8R938ouiY+UdiZTjpqvkotJteGGsmOZZEcM9
wVtw9SOJZoATiomp0Gkb3i7/M2g/EsDixQ0+L8L2HXlVCjZgmknTSWhehuELZxtfh27ZoxhcyW8b
Mksp6TYuySsfL/9wmK7dmG1aVUK7WKJgpt8PIZLEH9A8aa9dKgaQlYmbxkym6WboNLaSzMdGr+yx
25INYKXNFDP1x72pOnyCTH7gs2qv9NovBjQ+RwKg5GshdoXEl8lbFqEq7XidCwf3zh0waQEm63f4
LJGOfXMZSyHTp5ZYnLXfOauBwocn+ujUTv0KgRHROsaNDHHf4TTb2L2PBI8iX56OFR4zCKc9/BJ6
Pj8OyjcrgQh1z86vbVAojmpEPvczslZHbuXHGJhlRwiKq5dwEP0SSaJ/SJ6bpwpwTsPtXC+AhCfx
yIG6f3cdML7tuOlmb75URQ5iFBoYOUtU5MfBq+Kz1kY++egq9TqdUYAeK2VRy3r3JNfluPfVLosG
QLk9SbzDHdWtdxpu5xN+5iDKRa29qe8wkG9ixVaKcWpjznr7ZBuwy2eHqZCxrhEbShwjBNuFxjUI
XujyS4xVp2l24JXRX3CvHWZY1TF/l0r3GW7K11KKh43/leVXkv1Yx2QdJyUCyunk+OYLnvydU5IN
HtEgdwJc5GuHTQcciZLCLW/NZiy6Ky+07Tlvfr3V3ZElR/KMOylWusdL7vlw+UhhP4FisNYEPKf2
gbCDsHBQ3qCc0G+39ZYspU8eYHHsxxUARC1SrOkdS1aXiuZhXkVoob8boVVNUe01BN6h9MYHNoe6
Gxy+tD9yHaZ12lHTGQeNNI68yCAtCYNfxTgVW12hZMBJ5jxqq9gSy4Jq5pAK2ijsbkM2BBPqab4Y
G6pWZt5Fc/vTUvcrCCB+AcD9hTcoDx5P/GXtBoEHqNPh1BKVY+J/sE1zFbj38wEFeEva7C3RIKKG
Go51Y0zqEkhc5XUfbHXA12IOdQ4WfcU7F7Vi6ckyZE7XEJ3NbOIaaUHY7Mhc888f/rDjjzWC3Njo
FblK5mL+2SeMGJY17heiCx7yBO/vVnMbvwtb8rr5yiEMoUkOosWzmpRrGQhPCormp5DHXOv18rpJ
R5dEzABuYgYSIh6rdpqPUVWCr/0angx5/Siqugrv6+xuVSL0xgIWcbg3LMzDvWhiwa3hhQUGKWBi
Qmb3HahqG0QiUT0mW4HAvQB67SRbujzZfgCeiI05i7x8s1pqGwHxL2wpR7x44GjBD9JIsrSu0rsK
7pVjaSPiC0kk3h5m1VKGvx7/QoTvyIaiAIoEjFQXlmBWGBGNo+deMae8fE+l1Hfd9HdNIiNoLxZC
vka6brDXVXGAbu5nydU1jGXzBHEV/kIN/whyRWAKAatCGMQgq68nR7AM7heY5x7+r/3JX3Al+0Mx
ebMrtVUSefOQlyJ+RUphhlDZqBNy3nc2mxFy/BhLwbOjvpsiwaAxnRicbia1saqWkx14nxrHwmD+
mhxPdOG49NEiS+BGaP2NqPEwFoFOVqQBeKuu7s7ac5aa+Z53rekLNsjpYefk4dyChjay8rsSdWQM
oSrdQ2qynJweo1+sO8IZPOFVcc0kxol1BVXOYN9EbphjQdecCC3ijmrrCpKIo5wV9KIp08tHZfvv
yKGiI3Ab+RLF7mGQ75oI+IdeG3bP3xP1g7rhGBxvrnDk4H3YcA1eNQwBaxyJrLE0j/TY1LtPM3IS
/DlHtC7ywp+OFxtRBlrdriaX7CCmZM1LvZ42TvgHao1qDA96ZIzb2m7nnUCq+BHt91fYIE5bvdQO
yrQ9pEHHEo188VMenruqKGz6ayiqq4yNbKGh8BaGou/1CUDCHL4tXCd7BFeFdxX6Ub5mOkBtRAhx
uWe4iNJUlvZ4yDlqg7/qin8ZGXDXziJOvZ5u4JtbTc2LbDdtSEoL9GU+AmISnSZoziMuD9D0G7RQ
ynLLV1ASs/ve8Nl+01WkmtLsBOmxomWd11CKFHh5i9nydzyNwwC6yJsyyodu0id3hDKwJkCpC13R
vs7/QZkRqT4f/GdJfSnMfLWWaipyOFX6KD4vFwRVfID/+DSGx7BMgWSXLLNoj+mzu2myRlj61wTH
fUk4NxsBfCZ4ZOgriyt/mh5JhWPfe/0ktVCfxlVNMEPyuby7wypA26adzvYIEKY0ZMp3XqByCr4e
MOsH+xnqClrjkiKiIZes3wLcuE26SPzdUuBSeCu44tOoYMS+p/fxLaJZKCdhFhmSH9t6e2nRan3O
p4+hRSNSO7Qd7aliAKaOgekRDA9oCjrZDdSyzha7lzYOkJQLYvFbXxKXdVvyhmCkDYngdtMAMp5o
EbE6koEzJGR4oHxpseJ98rarw5cahxbgV2/GeT7YKN+0MvmvC8pOO1lJYDYY+uOca1CRmSJrCJkM
0UKSzsz1V49IFRfckV2zTUJUWQcQ6KVWT85e7bRRzNDpjRkkrzZMcvCSrwQWl7SPeselXfTk9HXd
J1snkd4qGtu/O9nUesPWGF8qwcAAnZjX0aPsCLFSLeguf8K26fq6dmwpXFzxf+055WyGvHWFn39b
zjw9v7wU+Xec8oL2b5z4HILfO1hcyrRXUuFtA7QIlJZ28IIp/BdoBmyaXymsRqkSe6PGBs86KOrO
EQQXGDvMGmeNxXrRZnmqQV1UGk1HZijnN/y6PAHEUZV+GW3ARrRWpbvv4QUmwRSvlH3VWZ0pURwl
ZFtSCtn5tD9XDRXCClXbqx/xzzV+BW/vhWeZSAci1aEYLCbirtu5QkC1yMk1NeSJdRhOVMAxNqhn
o/F8yfEcmMyjkGAy9qVixjiPqExqHcH3xryL7nQ8S4KLBqhg4plf1rorG1fY9DqwzMI1/0byJGlc
4i8UcP9wonNTTlIG5SAiidlc1ORTQKno4wTX9Bmn1ALMrRoRP196BW9+gdo5hKUHbIKS9XuZORba
m8Vhyzd1V2Ykt3Gpvr1O1rICZXuIkrHUITGn9OWKLlBON08DgGnYb0ptmEvTNSd62CYn21UaXSxU
dNESrQOHlsnSOTbzDjlGVEUw0D5qDqKnZzKoXXSfwqRi8NN5PkXbCsldmD5NHC8tDjsAOHBq0Ds5
eFWz3anQERdcK4biclSBlER35ect/BdOnfmEgO1HOZY0f0Fdayjod5pyZFHrUeeJ2HjilcVgBzf+
7dCSNphXWgxIb1rLw6K54Ch2ZYgg3rAbeRP5N+rx10s+f1tSd+6hcJyqwdQVKAg6xGXf5cuGwnfZ
wEWbs9vjBGw6b6lFAiwJEAQWkngpzJTSFozxBPVRKBnp7/Jvr4ohDOdYVeDzBYNiRfPF1S8NLQDB
FKz8pZZIyODI9VCDssS883jbqmpZ+rjYjSKnp+1KvlyFwogZzPj9+5OzbG1mQEbRIxKaew7K50Vb
H0DjFlqHnY0V2zXQvH5bYlvRZYv2oBu1o9O+fyROf7Llp6+EdvJSkeg9iH8oMJenF6lKua0XngFv
3yfkTHzUxmgtrddb2XpRdhLyMMAJrrrwl8C9je/RKbYrNEqGz6r53K0I40wga8/V3PTGGfmpokjn
+45cPkPB+uGsT7GU0QqAiJfE3yu95ON4K/NpuwrYkjThGKe8UboQ3riagg+i2Mud/JwvHkbZVpCS
sAX9kUDmMzl4l2Lq0zkVMHu/LJVyWXg8a0WS0LLgyVhYYU+bRD1OiNp8tG1zKBtII8tfhHZxAyO3
0zEf+ryqWL9PjOdQgY33LVXsYe1NBRj92ypAnaSXeNtW2kU6hda4CaZoWlc8Q+M9Gb153dB8srnG
2cpipevgFTG2ERHEo7jgmF05nsuoY4NbKk+8/eDqb8VReEAjo/Du3KFaEp98V5D+eZK9hnYo6wsA
0KHjg6MXX1JN0cJzU5F3EzkdLtszGrR3/N/fNK4kep7a4BxqTTJDnqQldG+WfIsqGBNnc76HyxjI
kuoYCpr5Gi8W0EKhvB0lFw7tRCenFjDplcMFtUqDPaZQBZIBzyoBxLQzHLz7ROCWcObKSwU/hr5E
GFNMshZuQQXXp6Gvr5M4ofM7cC7OI+gF3VkfRitB4wiPSvmjqENidfkNuYf5DYDnEg0TISi920W9
cTT3XqwYeQms2GO13gGBLSGPIgBhrxvNHD1tkigh50d7lC+YIZtCrJY/2irJVpDS1UwK+GfwNq3h
UroxI9WMZ/qEaWxod8kTBKD5MzulR67x70ZZonDNpafXEjgwZPBYEHTZk3MfKMZhpiF7hb4jyAUI
s7Lct1nNALjUtBOUyLQxYVUTtW4H2PnLsJp0Uq7XpxemztoP5UlEEaFLorZhQnF6IFKxTTwvX7Lu
GOqNGpM1rqguSq+hZUVaMWOLmCD6JOgZFHUYdtkwDL5Rl+j9jQoUcPSqrKxhjML2cyS87ocSH2Zm
NEkE6pMJyTyExfdJ5RdT+rbnyQ9ueLNeU3LZ3/Smd6Zd7ZpuiD76DCH+XwNNgQPkrGtbpZkiBpsr
ay1e03yc8Tb5x1yEqF4ibKCLp+WIMdsAlHoPJGU4iKod6qBFOo6+ZiDVireHut1i9q7lSrsUg/wN
3emm4SaM3D6agzH+hXNxG4hj55zIc6bBOcShgWmvldxEODO+hIbloKRgBGPt5PITMOCg1ijAfKla
ziEZwzxJc472lq7aQNW5WW3H41nZXaFW/16h7K13CpgXDlOBkNGPWuA6ZiXFNmSigzX2fPFP0x03
oLzCOrTbkkVk3ag/sCPACbmZWpoyswsyqLvg28M0NSA5501VhX5UaU6DX61wYs/AGB1606hpvS+J
2Bd4LNPBkEXerfuaVWqRMGmkP6J7UfNZw8Jh/n4IotxiHSDtvy6CMHw89ctb0KD4zaEtGlT1p76M
lID0Fe6ORI5a/vBJNVhRQGUZ8QwYEQtTlRpaQHzWG4m3ft6wEU30L8hJkiRCsesslQ9zf8GrJGq7
Da3HtvNo0ZDkN5aONspkMLNUbtLFW8Somg6aXeUEVj6i8cn67R6fVgGL+KzSPuXbqHZCbow5PV1g
R2unHa7xGQ/ThdIl/pTfOLxislL2ygJX3PShZAD+uF4i5rAG+bvfGni80BUovf7BJzJwTNlagEuU
PParZQ6dxcvae+2W2zuAoyaI8braC7ZSTKgXhzinRiMaac3YzFALDlkKoAaM6tS5UzzU2wadiOM+
XhvsX45AXuc+sMOnI6kgUUH3IlzcB0oWylVrqmS2yMS/RH7dk/xNtY1NsrhkMgbUgEdC2Fswmi8t
vVgLCrauLj78w9A6m0FCJZ2wZ+bRX30V5AEJX13wenl/nAkc9jsL7xwy0h6dqAlHRwMkliHdnejU
Qdge9HBek0aWmCML0Pu6F22Ir8fU3oY3GYswjk8zsFX0WBPY+JtL3FYILr1ivLVuDg1gPaFwMv/g
n5jiqnQneMxXuz5LmKvJnmfyAuG9sL7PVbhz/a+wliNb9pwMhmF4E+3n2O3IA11LhYwXOfT5MGqz
qHlysUAxVWCEPx448N+pr8ScjBQyZMst0KdgGk3X7mIIG75ycVroS+V4dFPt4TpfMnt2tjLIz800
mKviqN2WwPFt2wyjic+nYTw87HaXJDUwnDu169elaZOzhIT8bIOuZMPoCwpCTl0wltn4Y5IQ1UtJ
pCqfz5eLVzXAfrlPvGmjcBALWBMDUy/CIc/OkS7OXs9tfwS4mgMZQpS0gTrheDTAM9USuW49f2aP
wAYf2VmPSgKXaj2AEwTURVhy4JYdzJzFFfS+4gARjgLiPtZWsga1j1hX18km8Qccj6YvU6Q8mOEE
VRKhVNJrGBuM1c0iV5F3yq1eHmN9iC5eHIpEy4YiyZTUOprnNFti3WxYxuO5Z+XxpUWeCc6xmokU
vWRNXC5t+V0Rb0Ojo33HyzDvittJcQ5dpy/6tw/w0fDdzhHb2TL33Mt9o7lRm9+DekcpvMBhiqfn
yBZHWaW3kAOwAe4hf3wTWm+ezaG9blv8pBzuvq4QO92uqhX10UBeC/QDfDVucM8RPGPcGIcR3y+K
Q+wKC72U9dEzpiq201OXfeVqX3XiVBh/lGTS80HGKYbzsfhPWFBQ6WdafooDTtt8I33p4ZsJmEyu
TVPw+Afckms6+LTTo8FgUQXvBFs+B6AMtjj2N2L3Bu0F0R9X7nvgac9bdQIo666pjv/8ab85Zulg
xEHyFmybPWKIf3MXpeD9TPdi8b4OEKiz3aJDWur4lvN0MI9Kr0GFrwsh6MN7fkP1gjYDAEz8rQMf
g/EQrgYV6BQMVh/Ste7YCCvpZrm1tUpwNrk9RWu78QxFwoXMRl2Xwh5C6w6WduI3zmmIK63xvVHF
IwakvKcgfTz2jajk11Jo8PuswNq3/OPsE+xrbp+JMBrzlhwM2HA4okM0linQMxb/FCFV0xaFlg81
rfATMl1S8ksFZUdo5ONNKxGM1rfJReCEWX0tCWbh09dRSQbtq6Eyv/xUoh4Bn6TVYhQqB2vQcKph
LgM6hFKtJEyEiGyYwkBMU1M15vtJkN5t+chIwdgPCQpHfv2Dc9DdW36T9+UaWTlRxjIff4Ke4ap+
+O/rGRexNOg3h8rSJ3JrFmGZT0CUjvx6Hb/gnrVxEF9fuV/hWvhqA0OmIz9D28tcM+2/ABFQgRFQ
VUzFsbqGJiwPPlqdlAq0eya//hEsqTALNmCwRbGqrwapvNET5YErH6rKUkd3XYR0VcLLHNppE13I
WBXhdVqlNEe3HYrA59RpFaJ2hLkUlIQjkDhMH2SPIaDvXNa/G1DJYlGyE6LZi0iFZmYDSRoIjFHX
/bfpAXG05Iubb1oXS5oDxRPHjqV/gq3T8vOblWXuEBKIAWomvzJCNxZVxLZAAkdjGe4Byc2QcKZ1
/hVFdQLbx1OQ3OsuUS8ecqTn+xi/Gl5v5XFQE85Kgto+O15nIJqBKzLGFf0PwRmgaMp/9WA75TX7
MzcZhoXiO23QDwSHLIzy2EdkzsACH+1uJiKYUiw0M9xkK5hTB3p0zPSNPCmFegrStQZ/hfjpNO67
RNekTHT+mQhVzyOL5juUNxth4sKP8+Q8wQ9EAx+g62kLsAErpSn9LjJTQ6e7MiMoZBQHv1d+leFb
bjtmR1zHjp58bNqWHQeb8Zv1rK/zONk5/FF1VNAMyaZOwX2mg2NTI8Ue5WiPtIE8chZQY7KmPVVM
0PnHKCxH++cZ5BLA4fet1eayomDblALEPjW8cqZOpfqpibSY0/2JnAxn7RMlUrwh0bt3gFNvgvoT
hFITTfkYgwxLa8XzO5fXTEeDpFZEEWgCTXpoJqkRiGR2k0gkkQEoJcJ0B8U4CcfcLMegKUkALRO8
4hzYA0sUYn+oZ09wjnVopsUs7HPfDCr1wAaRCOR3ip//pATWB9VsAyHpebgDUEflRb3VIKMbBtdv
nc0aBWJjdEtWdNTy2EGw5d6qE6Xc6TgM1Md5uUe71Uolv5Ts+1UNpd89SRbSghglrz2r/bjSnvAT
yp4vbr5XSmi6FKw/1ZELcOVZEOa3fqDvsZozwECggihJhSzipy0DKrjrUWTdvnbKWMvdGcwBGtF7
TxPLVnnQg3Ej3RPbOnBos03CLZ+AsoPDa/AEy4zsDHVe1BmSbQhrZ7WQGtyPIO5i6FccTD5Ks1jY
mLrAGHA4xepExHPCaBZ/B2YoGMGvUgGt4QiLmxKArrVOBvYG1SeTkZZ2plQH7wmmnmLSmYbwrxFn
7lK8j2ircq+Z5ETGEePUL6yWqpn8DJDieow30MVj50nHhCEHwF41gD3kjrHHpYZTHpq9BdUu687N
s4w7uQfQLz9Kll+IuZiQ0qxw3wPljMJFCpGm+GjZSdB7SZOXph48YLen/Nf6lR8g4aozWFliu/sw
Yu3df4pP++FGWnxX87eGXkXMkzWv1ZE/lQc9SjdwCpJl1ajdePFveo30uRDUn8Fj0Ytdj3h/fkRW
+f1I9IVTFr9QvwEX35Wr9ouNGn1HIbLGc/2fkGuX8fh8tCf9rL5jq+BTekLJ7Jc2ap++10nV/zcd
yEwnVGjz0HMN67srQ9tyvANpfMqodv2zfQ4FWoCOMJThqyqm3jPkkWwMLK8GQPRENfFZYo3xFVD+
Z96zKdBmd+xpkbbabWIqif+J/t2KgCJCjgJ3dDvPGjoUOKQ7nTPpELTiMbVS//3RfYgibS4TDWiW
DG3ZWgtMY06yZbEO5OzAhBVySCdX1tb1zll2lt2fVMSYJVxzDByoPBL6yQwtT09Fr7hN4bwe//a+
PPmFfm/Twy9+BP2yjUvkSD21gQqb3lWzvQ/bqb79iEIqSy+RatbwbW3o21IdCyOgAI5NC/y94lFv
j3DPd/q5Yo9N5bmEagyW/jdQMLi5qbmkBTjXoDNe1bvpH5Vqxm3/7b00hTwW/J9ztUbo2Bu7yLFH
YpDPp40/3AE7t/6MnBY9R1o6aBhnzQF9iFefgepsKkW0nYXUVuZ8KXY7l8FvzwqjKm0F+U2g7Anv
RLOQm9zCoicrF3Is3Vdkr1R1o+ASgik5/J36N98XOQnLLjafeS32zDKC4pvkOTn2Wg3gLpwiMF3K
PzFFHWqpjUUkzcVX1mXfgVaK0vkn1MA9ubNSYsLZmOwRcYW5PmmR/LlvRZpeqIom+wcrXlrm44KJ
WVYef1Ew/xeP+au6zAp2vqx/013ELOZ5Gss0Ma7P+jA4RiwFV6L4FMlCHfJqTlhlCsbey1NyBGNa
Hgw5MfCF1TT116UqipbX8XrocRbujnA0LEr3YSXARSGolzz0/MHDWgc7/9Wswr9JRnxHpRSxnRFz
a4x8MfBhuxJ19gVShjWT2B9BMMEXw1P0RXeZxNnkUa3UjUdPuvV4SZux4TRWKOkUtOQbz0nykjvW
wnYvg2LO3a9smsM17LCY2iwiV52idWkONn85lojyq4G+cw/5x5MJAz3o7/H3+Pt++ocDiOgsl6py
1IaYSiAuKJb2pcBe6N4wn6mUMbzdpElSz/kqPJBIHS2kYqLXLf/OlTg3kc0vV8BQV+h+FvmOWzfj
Oz1GCUjaY+ldGEjPHiQN4biVuVm4kKhoFVgsaPjkX3D21LU2k8Ae/NXwfOssRq5jL+KFG5FRI1Q8
soOGDk0oBO19K+gU2bR9G3tvB56ilpYd8x9hM8nLDuCEmGxapLfssoKrQWp+eyDBrogX1uBlXkCu
2gCBs05Kvtm8xs2M6VQJWd0F5ADTK1lcPOHMlIa2heRoLPtBNRHF/yn076jY2Mc9Gz/aYNjoZ+cu
0Njw+PpdTix5Oha8PtQ5bZLyhpfPv6dF4CiMKW8sT0tSPALI2NsRQssi1H4UQVVA7fqynLbL5PKh
kSlaIpmHRZRCxfuRuu/i04aPRhUbTzR0HXuuFFP8IdLUi0NiCy2Ci0g3E+cJsDJRxRmzPNPnATxP
G46FjxCzCrR3KFWEn74YzZu7bwkv6VG6Dn8k9XnvXiRXKNJeO3tMsZgyIznB8qL2smjzxyD6FoSA
gsaOOZo03auSnDVH0ghWLtX+gz91uPRc+LoBC3yy3qK2l7IB7ssKxvgQxtYtLZhS0nL+PL8/a5Z0
yCx3/1SKOLqA9UkBoLcKHzfJ8JMf3TVyobiTnw+IW6DxhJDfCvqOIIK494YtxkezN3VVLBOtjA/8
97vVVJZpdZPMtGLjCPi8QIoVGrd13T1PEqvjkVsQF265A1IbddsEH84vn6rqeI0hPl/e9pZHAeFr
ij92KjOQn+DIZJqqTJtUZ+I+z8MDsQv/3pdOrH53hR7Trn5dU2cbmj4b1h+vRmowCpSMyzK50wb7
0aCEO4aSpgJiDyv2eP5scWhFAV+nkTNttIEjxri7hAviwOghmrdla9y2vLEphNq1J7q5gPyPIbJp
dFQVncrYZnOD2/CKyIDCKbITgja2XINof6OpXWFk9vHLMD54/0XlULEXT0EkT+pI5qvFya3zoDbR
DjeNo922Fmz87KOQYVoEHa3YZFQiSW3e8M2ICOtIEZs2OwKM9u+cUPcHd3xWiUL6ciLxW5HpSiTc
PeLxt3qutWRXJdnycsyiADwmlH+4/NgGs/XWXKn0Ceol+u5q6PDRJHmneo3EIrvny6IcnK+2jLZM
6qKl7iB2e2lhS6XwmQruPda5CFG3NCzWKxyV0VtRG2Ffh/vGzg0ZH9lhopOZr4ceU+S62Yo+3mmz
EOF4lSt2CNuVvJGbzhe2SvdnP16qqih4XAP4rEsqwKxXWp+PetB8NKt7YRLNh+OqbpX/Altodgco
Jy52dFJ5Jjbgga4ri3TB6Le6NK3SSfYg2v/zZUlm1luHhRl/PfmOHNY4kGeQQcrcuCNm4uwE10WB
Y/DKdg0PRWE3TCHokNJQxTTK1wuhOCHyPb0ptcCtXFtrstZwGQ4eHW2xJMG/O4omYNe0+VblAgrP
BjQKXYlMDBK6PJgPKaXuKhWxnrj3aTu3iSyGWeSek3lhsBrZXSSiYlcJWKZqByS87nClRnvDRYpH
h5lfMW8sp6ZeFXl/V2YaS+cNNLxwyy6B7PtPx2hGRXr4MIM3V/8yjbcwhKpMGt8QhhBHxPZr4E3I
7k/JT8NyOQWd7gteJMxSyw8euN4ZxKjfuJM5KhofiT4AVDzawUK6ZdfUbPmLK5pTw1gOjiHaIoIc
g2bD+pe+LIt0Ky+Sli4JRwnXvr5FdEoIzS+e2IufP7dkJ+4B9lcYV5pFKdqabUK48wCdGvMwmtnB
g74zBAnLPJ98Zc9fVMFp2hsFB1ExXIDSqAcYZXzUGVdSSFE4pN2RoGULbi657KRYRLymt6fLMsQD
ogIElwRNbP+zW77+gmgMMCplEjGIU+9Yt8tVGj9TvINVhjn5NhZUHMA/UAK48P1A6ntgrecGOIHI
amRNLJ6dq55kCNhx3WZuSWLHIL74qBzqxJzTibaNG6qTO7V4Guk+1uc4dSWa7zckKk/n5Pii9QFE
jHh9XIa2kJAVnLYNC/FTNdduDH5g1N2Rz34zI5V3q/nKYpmQ5zBk9PpF+mFmoSzD+jWKSDG1QZHx
x5eimyHL9tLdgJmYQxflbLfqXTYcQF/qbXnS4m1vO7cwlp0NKpB0yqX4W3D3j3mdft6remv7vt7Q
QRDb8ka58hAMZQmG3H/AHJclrK/JuMj5BmHLvjpjstqPpxvKTBpDWaHHL+OZka+pAjMWB7Zy+uNg
Nnh8Q/q//4vm5MURmKBHpDHaoXEcsSHyRTrMb+rOpRd4LOaNp9EVBZYd/nhZQH5W0hArddDj2U51
ILiuFfxZtScbDRcbNGzXHt9DqF8eBAqi7gyV29Z17+8hsxD6o/g7MDME5X7s1cbjf4Q0Z9cuNvzf
6P/jbYQ7397be5SQPaR9ATSHcfQTW8DeK3a0Mk5P5lT48HPSx9+waZUAByRSY1BQtl82JzfSSZ22
LjIUKsMssk9I55PNHX/4cK3HWOWFbwS7/H7RKQQd17ejvSB2ln+f6wtuLlOAKAZZSQBWpaVL39cK
GkqT+NqznrHJrNYJpDGjx9E0LrQM2TaWcX+bkLUgVFH4Il3oZ9VXdlDQXIKlmF6k0bLgdur26QdX
pUKGQwxEJM8NOw9gPsA9msuM529UC9suiR9SXd8y24njcIse1gjaxyo6pWuf7MGDer4wnAOzgVX+
AcahUfAsOcl74uhw0PP81b0y0yDjZbSRK0wOtJAYxxgF0736uzUiovmAGW8PrG1IRbNScviwcKB+
LIFATOiux2rKT8S+2JJ/HFJq5tG2DAA8gj+nZXgI3JbEIAa94+Bl/Ca2FTeY7l8/7uuBCuEyoNEj
+qHU+bvCyd1xFlcqs9IoJoSloyXlGaI0puU/r/U2DX6J1WOgP3E/yiUCUFwjAxRlBCsmd6iAYiLQ
G9zpJKbrX4WUhIHKKFDzo2JWx8zPJatTaXoHaTZhvnIKpHz7V/ST6/NeYD//+UenpJk45Dj8Q/ot
534vSiXabLO4isgh0Wtk3/71AmCHD+sHZWC2o6atUm66d7ms5eluMG8Tbq9a40mB5rx5gvWb3TKf
INgWmvN8vVUvl8nEsu/OcoupY4M+cfwYVuIp/TsbJVXeP6syTQEEYPFzwbmDt37GO0RMG8ndvB+q
XkyiuQWHiagEwTdgF7WSKokgjnS1p7bafmYnXfJtbctBy+b2pphVUYv2vxb72D3OouVxy8MV9Bs8
Cv2LD89r6fYZMPs7do7uDQnpvh1fZNaM1Zzm1HJw9q4X8WXAkhyMtbirULp1/tYYbyQts4OkmgK8
g9UDS0fz8p4oZwRxcBPilWx3wF5QuTmWxtdw2nv4NNFhWm7YZQNdl5CRn209EbRXH0oVQ3FQ2UMt
h133+pnh590//dQTOMzlFipbBrmd2rhn22cgZAJwuMAT/XdYyZ2kRd9Bm80G7WDA1xCwQmRbNknh
7/nH4UaCSV3GQejunzxnEDPJrTj04V8tyO9VPegqNvwbxcAkCUfc7V/DcWAXCVMmJH495y7nfoyH
T6MAFY1/NmJ7PZWn/o2A491g+yXJnWjoMJmsN8JeJx21kAieEsxcXEDI9jNKkeqsF9pZFSycxRZ6
u/8lV5QrhptMjafZjQc0YD/leNof3zF5bNFXdlM4lhJ+yt7P46mzactVEMYfNNv37MsRMiyqmv7h
txlCFmoSz+R/9gnvMRaPGN6r07A2jhTP0cKAbcR4MAafkiGA1E5vufZqXxrsEPJPlm6M1o6FcFLl
qRktiS2MUeb9ZpnpIc7zFVU3Yjms15yjlQ6dmv6sxHPlXBFUtDZxCvu88XZZV5Z9fzGqS5v/usJD
GkSLWpSyd49LomV6FwNulKwo2NHHZMWmeENlPz8ZSmZerAJBscAiF1tV7Bi1xpI7rweVwMGCqGeA
UTlNAqmf8u/ZmJ2IIDtpjwK/plu197/Kogq1XpmZUvLjgYnyWKdNwWAS9BDUhVCzHOHv6wfKHGxx
DwdR0W/4wIedGRWhgc9Lqv3cw3IvYnBMJmezhzNHuHUb2SqeC7OYMc+Tx2aUtDhmdZhw4WBBQ2lk
EbkjBHQvzdtetVFV5BPAaNgIAUnTyzL4tAwTd7rPjw0T5MMa3Q9pMyegjhh4SMepfqgzBOzpvIiS
xjnd7N+KpBnzFGTfmxPD6Qck7monU1LLx8+bk8xZ7Ba+G+lI0wzpS1MTnf+hPbRAuSSuvXingjyj
eKbvDK8fnQIowbs+P9xbqWAzJmRUt4M66uSek3E8hp28vM5U2gaCAs4/Yjaq+4uVK1uXNDLojVCq
epLO47Uw3DeeSgfU+JsG7k/LOwgMmV0pfG+5Lrl4E90UMaHlVC6/5djN7zcyKA9VwWJ09TTfhlWG
dX6bNKIVPVR2xu/kQXElbjkpYt1gdcgT3Ly26zCTH9guq/A3Q9arB8ECOO4hRfNsVPHhJzu2qcAW
6j1c4bX5eltm21ITBJfcX0Mi3GvsdMRVwx9pb3a095FSZgLOjhQ7q6AOguYe22F9aWgdI/4+0+c1
QwRzh6g5D9bsOuvgrVsmQ2Y/eZ2Z77gWEfUQHDAFZT1/7a3UlUnNeeXS4bBTaQcZIyp6qEGm7cqV
dAkoh16X89zrfwV/Dp+s4hf0vO/bTzmb27wwPt/jRq3e8/yIqJcNO5j8VEFNDSdTK7qzvdLZYL2L
rEDJYtaZkM13tp0eLtB6JyNFcHE2jIZriW5/L+Gl8cHQjp7Cwe3KWdOo82O8apbbf9ri5QjJL7fY
LcQGrnoG9zv+6soX4viN+GGrgyjw1QIdBWwj4wZhyPoO2/h+7oB9sfVvdqaqQ1kLIBKGlhfN1HbT
l2p1Hx7wcs4g4fofuhi8bNOEVRRUDO+X4/2I0B0pTveFSnDb31yrmKli1p3dr77CocaJC6K7f2mf
TGsYV2Nk4ZEoHrLX4hdrkIHwpT1V6Yv7tCKURGQ2jf+c078uESTgk7sY6nIXBmFFf7P32gcISNoZ
GlM7jNKqY5ubYO/iiAgGD5JtXn7UxEMyJtRs8R3X4b0mnloRfOfuDFnGQpsd2I99NR1PZxSSkGDx
dz4bXVnZa3jdfcZVGNKKiU1pFk/dYTmc4WosmmPtRs8hSRzC4go6NbjvmMCYF5/lfu1KDZN00ePT
Wfxn5mWthTB9pHtlxK8j+ECas97mELYKFNf8tI/P2/C1f0bP7PVJNuEyzxPy7yAu28mKZ5PunM9p
O/6/aCg7MeJl5PkHZb7mK10SdOYBrG5/m4VMJgYbx3yMYbWhsdVjafZZ7TzOtVG1I3VBJSIgajYb
imx9O+OMPVSScE61Ms11gd6yF9v8nb92LXBuVlfEBbzFrH9G92KLDs3qyba7m7U0Caz8XS9cF9Ei
8QY+c1a8GX+HXMb+vmPh6KWs6Q0JyNltXxl0iRwWqPNDhcrctKLaNK4SGHOhtb/3jwpzLH52iI6B
tCg4s9XBu80By6OI86PHJg0tRKSQ0v54lMs/hVz3XbBPTWanuScfDSHNsw8R3GEU3qLBITLSn/ja
Z3/tUvqhoCpxcTWcF4aVc3TQS20hdAamHoil2UVKOmHlX8qW9WqYg6UOdtA3tqVYflXW18m5pwql
k2iuRdqEITfaU4RVQfIz5Xo44Xcx1qHGU5MIyf/V6VfZXO1C08jQEdPgmt1Dng3FVSU9YmzMbjqV
Grisuil9IcqcPEE5al20bhPaPf1g6IhXepFT4C2CMyxdPdvcWNhvJQHvuXGTrHv2Xfm7JfRt+RbD
AFYuLs/kvpVuKWRQmMDgvnoYjjQtOaV53kGeiObXeyv1mA82SZ1KDFPKAGqs/CY1lhL7RzrPTOb5
HZHQYn+BnLYcdiQ1mOP/sE6Z8mebtDGP51DR47SRRutlTGZFd8lbbsCAWAoLJ/ANg0hkXHCyFsfv
CJLQVQrl/RFNoFBxT+SmOFjCYDBEVHp9oSKd4Nw6TJt9qj0V0Q3SqBYtwSyPxGDrQA0pF3J8n9aN
7dWxKnzEJ++vTrAI2sXpY7GStChHPRBz9fVKoa1AAe7JeRBsn5+eydJQe58h9jwD0Lmnw1RN0RNA
Q47de9qOEP5v8hahvCxwhR4tRpkEn23Kc5gUEV8iuWPWmYnkRk4ZgrFpwIUyf/nj8RhWvSfuRlWm
LtwkmkXb6lAAt719Ot39ppYVHrsD5gjzoP9r4sOrwF1YTJyLG8Ll4i9qUohDcpe/O50xQzxWx75j
UeqEoaQuJb7mM20L5Ganee8//LDHX+KhFO56DpH9AbLgJAz0lDicRTmBYXiblQ6IVvgPzoKHVTBN
AzkbrdCphtZXTDbijDr6EHXjgDZCh5/ULdGUtoULBdKrosPjNNSRfUwArWmawiJGwEKOBLvWRXTk
yR2mIJBiEOcuVorgUTbjdm5KU2cdgdBoWqnh+0vscxi7s8Wdeb7BSYseezxUSlH/KcdD87srTyUF
nBc3jDrcyCDvI9ILRbeRpPCNdjkCLtfQayNOlzpw8STxZjOuNYWk2QTIxixXGDHQJMAzpGK/v/XX
0XrmIvV0lnP4lVAH+RJO9O8yLF0zy6vMgvPuG8DAZw4bxQytvogytGO/n9k2XxTgkHNPCmZyCmxY
vlMIgh5Qv6IHq5VFlEvWCYyFbhLIhj2DXRvnukCWS15nAhLtI9OXQHdndblRkSDKWN3rmWRHYHDv
qmBHMRmy7Dm3n9f0VrVWIdNmSCZexT7Zk6e8eE1oCvWQHPRQ1jfMCxpwkz71cmNjnUAUtaL19jiH
NoY/Et6wCxGnJyVjWFfvYh7tWkh5XvCkkg++GmaoeEHk2QdDR6OSUmh7Qsuc2JdZfSY6ODCdez10
ilEQ24BlvaO2m0ynqmRcLLvNs9RowTyYdKZgpcEt4g6L9AzfFByWSh+FK9lCH9Ph1AWUc2ID7ZVH
nUax2suGYAZZTPY1oaRMuMsvCgW1uSYnZW5yTRRWWXbxrR0pAlxfuRMMHhY06Z9qBn2OoFOJg9aV
NjU9HHMf7yqZ8oEalYvFrXca6dbDc4DkyYR0chebnq14Cq1VUlUB4ZbzKU8P2Eh9AhRzkk+hCaYK
8/rksnOBjZys71//d+AeW+Nz+i9++xx4W5xbRpiczIb3+30DO2ymUoYpt2DsgfWw8+J/ebOW42r9
7SfHoG6yO6TDypqhAibUtyMPvlJ6fa/BkgI77ISvTM/4fJTjyd4+OvLxjWBSYJJbJto6TnPGmH/I
uJHPbRmctbyOOrqWuDByFTYa/eJHjGcJwNZuD62bAiOw2IHCUYQsiLPa2yR9Lxvf5wz8i/PlpAN3
yEM+CFErWj/yP5VTkhyKGGUE6Keu0KLVc4lPNkZkd0vHW9hiVCmq2uUrojPIcZVixeZ1GXczvIrL
wSrJa/p82xFEpm7ElNGESdcgpFjusWyi9eCNL5eOVsodsD025l7TV7FCI/CmAGaecvFeV4MVXsyn
DVAiEWhUMHQdStDNpLN+i10JMknt5GGvKXNKCJpqxucjcE211hzagS5rzW+TKlQPjiPEqujP1PN3
+YO2mx/1STRtceaL1GgtGIA5tLJxWedEIZO0fRnOC3tSddr964IRr1mupDfENACK+v0jcd50zfnJ
EKYCxUN5E3ebSOB6oQBJ9q06BjPGd7f91Nv2whoqdoWz0JUEMxxu7CqOtzh1DsSovJWRlk+cMfm3
37KrTEDWGrBrxb9oIRiIJDD6OQgjjnvl6cDKHMlHT6b/b/a7PEenKFxcsOsn+dFKkOJX83LacuKe
IwYf4tAZn7bigO3KdSG63yL6rOQsmRuMXa/Kj77vPZ0lnL9GN/mtzQffmpmgnkdl36LP1IQgFALq
R72vHJIBPGpaLIZkDc6Xb5mwJXZ0s/x5XVzKzRmJYbSuPGxULm6TEJ4XeManIVnHZUpRLUe8EGmT
z4+8xWtPHP8pwUhkWsAJKVdEYlv0E7g8/LZRssuwdP7HbcXwLiUXvRGWU7GJzRVmDF3v8EkLdAJj
gAebW+6TY/FfSnBeK8J/9bVAp+8KR1cebfWpjs2HHUco9Bx5dd59DsOeatQRV1jK7UJZITOQJjb2
p1qC3V7OLC0D8FXnA012mudM+39tS3LuwHiWOfWs+0J7yv5YcgSDQvdDBxnBA/GR2jZYqzL7rypR
vtRsYr5dVTMup29ZDmS1pTJ5Ljmwfx3R3F8R0JS9PthlkHkadqlrW37nr3KSOLVuV1wU/jD9uRdc
l8SnKj6fgXaAMwG/X7PwHhB1aMcSvNa+QGpYCjYEe54XaBdDYXAMkXtGKG135uCO6UlSAqA20gL9
+I6VMehTBmuXBKeJ9Aptqy8TfBe7YnxDAi0PvDwJ6uq1WtqeP5sxwJw/lQ+DF/eMmFZ/OjcmfRqm
3bMdohCdO2JR5AGil3eRxvsOXGB4IHcc5VnLOQnQVbr6xP3EUHqApPZ4Fzt0aiB7rdzswRTipnBk
gbnI9EHdrReXI5aN3HkxjmNj7M52pK+cf0oY03wV0KPgEUxpzNg123YYlFJTVNVp/8RJVmOt/+RE
BLOA1B3nkrh246xx6F+eV3C3GtJb0LadO45BUbqd9H8sebXl3W696keRvbMVtj+y6fBMB7olxWEZ
Gh4oeklh/mZTEE0sWxVv3PtKgdHZhx8fS26D2JiZLExejOIeA9rZkLeKWo13+z4c5CsvDzRO0VPM
Z5cmrPd++v+mc4/DKCXYRJkOPWd4IfePSKZJXIglmTf4l8PHFko8qcqhEgMXDA6tt/7e78xiXYnr
/vnZaK4OVjGY1BIDtKeJLPhQt7BEw/IylQJZcOUInBFeOy+yyQSqjCi/QJVQmChpJy5dcKX5AiaI
/SE1tGn6eCRJqEFZ3jg0hUHY319P9Eoco9/6Au1xrEbj/6S9eGtXtpoKlfzAP3iZwC1FrMptrB2Z
f9w3h6to+/e+igM89tzvKiSUjw/pCsR8MRKl8AVaXf4XdTz5qnE/Bu0664mQhBid5sF2Iyl92sQ6
gfG82+dNKyKsVomrRBLELQbUdedq7DBozjefBrOasP7eyZ8SRiFan1htnTpdjplsm/yJSfhD/qmJ
/76LExnp4pMDjW82NbvQB1uy4dUpwS8GcuporGC2Yh6AriotosApsVMZu3V65FyeYoxwYLNGcSlk
vBpTwW4iYsDnHoLq6GCwgsTs2Cw2BNyZkq8veu90dKjAqz5E/KrmHMmgotW38Ll/fxsYbf9XXN5Y
Nya/wSZrbtM9hn998ZwyW/IBuZUZgDReFkbuG/iqoWh6s3o4Zl9eO5VRVJo+foiC3e+Mpks42+16
n17HwtppOVcpJ2mPQgdFITdQ618mVUwmevF8S9h0lxEX97D6vCwudFZ3sCCUUTSDLxSuKQSU1Yjb
KaoKBDrZLJtQwcxp3/iGhBjLSx80giYgbEaS+aTVwqEyBIMdB6WYnyvlkQbFQfmQQ18rgMS34oUF
Muh6Wajp+/b91oUTZeKw3qTj76+C/Zj1PqhCKxVjvW81Tg7ixloYaqqwtwXvgVZ/OD6MmJPnyao2
8CbTtqPhWrq9p5Ro6iODZ4lTjghZ3iU6l8aUWgBZxv4DpSnLI6HKg3odrI+s30j+4T8xA++vkzQH
FE7yWX4iNFeTgckLg0fhkeC//lFZs+cT1Hyz8djIaUxnCM/BM+RgBUR6VDP29MfrrNiJB5ZUebmh
eoP4vR4gUbEhRLlFASMfcDKtDxbTm9WQ2unb5p+HKZs0ppD5boKKLBGswMWWZwAWfIgfBfOPu90F
fGuP4eMu9ZgJBcJM7b8+orKMttfuhwJ/3UyDk4JJ92YKHbuhZKYrLlsCMMKHcnlYpNhff2Qw5EI2
1ljp1rO5nAngDcqyHQsWDy0aDdnDQuJqOJcGpvoogHgmaUR1V/PbAWg2enfahvtmxcgPE5AHMWsG
BJ5Ho6mPvvAid1NgIYpbwEl4P0uNimgWqn3GcYEHSby5xmZVXfPdQgZZHHA7W3B8t7aVD2EYzwt+
C/ulAVyHLljvjibpw5sO9zuIdmx5jt+GPURsevjAcobY32k54xDfIc4p2adSD1aAHgWjtnOUNi+X
KZBK49vi8KFGg+qbKVfPwvPpj4k7FU+8OX92B0k38yzdoCQoiVOJa/HF+Tcd0WpU/K0qtZ0Sn4MX
V3If53Dt5n54/WzmcuF/oi8qZNN6xPov5zuJnJvcBTJtNnCD3uq53oMSDKUDmIf7UCpD2nSnBcBa
Mbsz0m5gd+laD2ABLa+yA+6/gwL4jmCBmE/mOngNWqvtBj5qIvoXvNIWkntMg8wUkp+TSldIgxPC
fJe7D36MO6kYbPxHYFpAWzWwjYlS+g+sgjyVp4ozN3olCiz+jZ0+TyP/6WEiBblJGy1KqtfNudEH
5zYrn+C6XxGSv2YA7yhNkJ1gjV47v8Dp6XQs5OTOQnxKU6UqNP1R4DMM4wY1VHAYgOgUYIyjNVtW
xNxVZNd4oKY8Qz8tpRDlPpgl0H9r4cV+QtWfiuEPion95z6Wu4KNXhVaJr5otlflBXNgj8h9qGfh
ojUnwrEAXKX+XoxULQJOUej3MITgV00J170kyEecoBmW95g767qbmfMJHncJJX3I2/8/Ob5qDDl9
8TyicdJw/5Z79vCrW8NOl7M3Rw0uXYyX0HkBgKtwROCqlwhcwp5zi7spbZfLsYF71gm8p2hHJcKs
p8q61JQ7TGNTxAecW8cUDMClwipQez+0EY8as26mT3KqGSQuO0qAsQ5yVDXzvI0K3NYkZpMxPtbw
/UsQVmn50KfcHyDGBU9GbR2nG+AB0A6cfCLaFzjQ94bK9FBzcURCnMQYQ8fac1Apx77c378XG/h5
Icxm0jfK68uHSWWe5iIxss3wg7vwNAOyyVMMJE+Q9uT5PHQcxN9lN6LFHCFnvBezslzgQKvoTvDY
BIYTfR4oY2/Zwfilo/4aDDJJolmD/epz+yk0QHtSyctoRF1dQ6UYhh81P1Jtjrzp2k8c5EsbxbO3
u2TukGwKNnlVJSSYy31RdRU2gQj7xfa4qDCXruMvKb6wTlIRx/jb2y6M6tiSjTmXj6/QqvEIj2aP
WSYvV0bqMO+wi2p48XY+A3CkNtvBpo0b8Fa0fM9jTQsPCjw0kjlQbb8VMcocfxtNSuEOKEYXCgZz
RLZxvAGw2lHBdthgM1+vLPHonPGMAEkOqiiwOg2AfwYHS9hZLu93p5jimySzUw1wrosL3DGVCIMv
Mh7YLWeJtWlPbkE9/6JA11xU1jKgKZMjGqyugV+5Xka0zyaFOs8YwRPXHlh4bGWioYQUE6xAnR8m
2h110YC20KLb54GlrJ/JTaUfl4+wwduF6AT7Fz8m5RVqRzYUHBZ+4mUNVz5LR/yYArKSialejouX
HJSrK9YiazEZqgnP8AKQlMN3hpCMVDryGrl0jCGUeE+vRTlumJLf0ZntsFKp7VeDXl9zXjaF4Kob
VlmJ1DZNDSgDFq8fwSBUWKDD964GL4th0dYaa/ApPtZVjYLFY1p1ywAawhiryhmnmGR61jf4C9C6
4mJrxHJEYJ+jY2rMU/2DyoN4JCaYTFaJeffmGPoOWEAMv8KFPwstFAef/e1I8ZCSW9pOB1j4wJx1
6XV5hKhoE/hqKDcxVL8SX0zBsD8jJcjxXQPvXt3w4/f14D7WvAJqCggxWAEzmNAi2oKKDcPnFqMn
sysOBkaqhIpHVtMfQc9kpqh+JdQb47oKz1ScNM3lDx7RoIjUCh5msPExu5B2njnkTnvhxIb+M5Ol
VJnTY2A57ll2+N9G/pRHG0FBYmkgU1dZU1ws02e7+spWD7i+KChbpwJi2nLoHmdE4mKu2qS++1CX
UGsyw5O4lccKaIogmxpsNrrOwGdU/GGNWHDxQYwjw6/+9ioXomh1qv2uJOt9CXnTGPaxAZ4F+a7w
w432MX1chwFg/3nLScffIqcshz5AQeKy7cRba8eh9aHG+tY4rtt6x74ds6pQPM/MkB/GiShdn93g
pNbRQGN5yK31SkLWVH13U269z9iTc2dyen+eBZoQ176sxavODeHu+c7uciBLxn8vXFAirEGirfEV
7vQ4P99C2S4ZEVYuitgTtRKGFuJK8BS+7y0+1V0sodZXKhpeVzCa9BjPUeK8oKYjihPDwmvifKyc
3l3iLoRmZBsG/olHwWjupnxZ6wfatFoiBCAMCidYPKornEY7OYqmBSc4EikOWmzHrSp7897R3Vmc
kPeW6JyUt43BCun8s9gnputIxnekTAI7u21KaqR0qMk2t7MjNfa17A7pxBWEhcd99imAfj50vxfM
s+85x6q3vC4wBeiGEyMTwxUpWcvL8EHciJhp36IQSQzN5OthVBYT32h7DsZPxxF4hQKsr8X+POrY
+iWC0WFFl4czce5jVs3QftEhZLM2qGAQUslVnvH887egKcGg7pXP5t/6rxSHAEiu/sa04KnZ5XHl
aNKHugvmX2aDJAVicBy5f+hTR77wcfBOZPEuoII6PhAWSX2WiW2SXmWGxVFNXTA1nYVnyPHL3hy5
GNKq2Yx/4nhFqOGtGceAfjei/hyZePlmNfgY7B0gV5YJ7L8z8mp7Q9OlM6dyv2s7c4PZGJ+a7Z5H
ICmzkK82KYcDNqygJtuvFFo5gP5a3p8S3txYx6dqZp1KDWTiB8TBhUzftcXMsR2WkRrzzUlvTYlF
BTvz3SfevJqJO/E7TvH9ZI/aaCxzx2fywd3+6KxnjgBPQGBuRfYF7LXePxOaaJLIrRN8SQgO6xvB
INYuy8HHHT3yGomR+zF5xFde5LTfmsepVSQPhXddIkzYYiwyebMQSy6JuXCvkhsLNUP0WExBYKmP
6oM9ZQLoX0iz47woE//zBHwoLFbZrXbYPX3pcXplpxPDSxhcnAPxOM2NqvU3v8UrLp9/jFstmsYq
nE15Zru4ZUzWAS09QKubaDpuIhDumZjWk0IMhSyzvXB+MRkLZVrNkKhtJ8t9LOyCR9PkPlSGTw/n
T5j/ep09B8EW9l5DP7MtOUrtOX+9OgyvqQm+wKMSe0NMaUilYvOQOfyZYktVkWFqIH0wSbL4Oi8t
mt8j9MRSMiZPIsiFF/RCTq5/e5i0mrK3ezUL28RBCG4ENiYJ/QaxbNGjFSn+DekXcmM+UusMEDYY
mSonViROyYKZetpjHieIoiO5eepgWceXNJvDG8vxPqGDU9CTMzcDkm5b2yhq4xjSfTqdmK+PwLvE
k3DIQ9CBw5/kOhccu1S3rZAes2Unh22nl+QnVUvVy8CgvPaip6XtF5rzDYg2TzppMPqUoDUPriU5
LgN8lQZP0Itzp0RPHbMN7V/IDHOBDpiF0WPal78ayYfFUFB/egTQEs/8J6wyxA/fnOC6opdJIB6n
yJX/IWDRZuXAwLWdKOW9ZikXURnBb2IBs/ExHd1PZgPGk/2kZ57Y6zmj8lLZkKohayc1XVh6fzc5
C9RHM2idp8fA8I+O+Va7YlqLm/WnE9ilwVM117PRdfE1Ru2WAuhQ9kRNDC3HcwR6zU4D3LnJ47Xp
aQEDMPSNpr3y7iRYLF3m9LtNVq1sETYYhucwsyA4GVJ32X0tdbg2b9dlZbTjp2OAHRTHuNwa/ioY
E0pfDvJcsQ+CDiQD17i7UGAncNvyREk64h4cD9jnbKu7hAISyp5mFh3ojKr7Ji9OleOQuCLI6NqO
sdfJigXEHxevrm02Fs2AgPZJ/j4B6qzynhNALmUXbuIwkHuI+opgFPmsHfkv1kYj8AxP37onyxNS
IECP40317l8Bj1oV6P7WJixgQfDDO2S7rOfo0vCmGeZXkMBpBpuhWf4hWeRu7ZSMp/lgY9ZNSteZ
V22rEYG95iPkeyoET17oz2Y2P1XTKnujhtenjHmN51XzmfmKV9frn9DwXtDktlNdyn8X+0+gaM7/
xsGD4d+kpC3R7XilrIcMXmoL4wvCLSQot8brtRc7+UejO2JAPcXU4c/8mqmqPhfx9Kxta3OKvUSi
LJWyJV2AdpGKItG7Pc/NSySM3s5do7F3isAwSwXZnmlRXHodcQsYlL4m5lG+7baOUN15o+jqJ1aN
9LkV7/mOH42hYJzLetwVbp8q4tOiRjlyOvyrU4gtPh/UPyD1/fLWYZ9IczUxHKdhS4Nyun4sJFKP
Xk20dRwYjrowsAd/5/ZRoLsFLq6YYgAErDRk8zxjITzn/c9gAkfm+EX0h5URdyV+gvVLcZTiHYKi
WQigzKImpzcXBZglY1ezmUnncV9XFvqdB5V4/ubuC9l1XSDK5LURo1Pcukx7Wng0lSBpAr058lER
mkgJN7eBr86c4ZFv2G8tR1e7wCduYsuQ6ClK3BZ+b8Er8jFxq0hwqWVkaW6SZ7jCe5qddt+48sQz
92gVui16mDxfaId17kfwwkPqQWCbdCpJpxkKAc6TkmLndwfUJ93ILfjWPS6jACnxXpv4Eyb0Pvhk
loUmnFneZidUSesnoGUGFPDuOPyfPmVEXZ70wUEbCLeRj2R+MK79cqjOYzsIRkU15EyWclBE1M7/
BqXJdGU/sI4fuEZaLlgQTk2QzzA10yqTOI2V0B1DzAIvzowtBOyKe8s9LIFy42U7EGfLNzijO6FJ
xs18cDMtg0k8cioKICh1yTrfc97rlUUc+UuyA40TWi3YdpLxSNo8DNQn0Jqvi8bNtdLhlt9AN6z/
rDneLlTpIlh/lovshkt51Th5A6a4BrXLYfUc4hja4MWDTletxhPzCFSFKzAj+Kh5wBk5Gs1FWNPk
macIzeFTCs3XdlvgKn5zVFDD53jM+qkDBqoiVXsO+f0ZRO+S4uHMd9RazGPfZLcnUbFtfDVoKuAD
UKnpx/dbNg4CJzUb+0sdbPmiZQKvc17QxO6HzzZ5ACAgbBb5YXlCqsanJbvd2RLzUTKS8tCsxDHw
U993M7MXg0OfZYlsIBMAMW+wkuOsflen2sgPgvyo00CYhBwcrfd7yRsKma2ON7ff/CKbKleV56/S
8jIZ2+67qDQJk+dqaKrfehsF/Q4iPiwYN8Wyr/Uh4WfN4jSzlDoxNN+qnYhY2w/20mqAFKR/euPa
xjjg1orfhfLFHtpirFIiXI1DXuGqKyIzSypAR/rWN/2hmEpTD7QH5DT8lrEpXlv74aOcXO1XsUeJ
NPKmSkPzPW24owfbGz0euw/kNFL0kqFcEIYt52hgCOj74iFK88XZOdySCVCPjpho6TofyPRiQG5R
/m6Mhyl0wE/vgaZD3ahJA7Ta+AfpTmXJX701BZN4fBQUxpMl3lXBIE2qEtdEh7VhYaU0m8ZwzD3/
7DQ8KsiqEYdQK0BXz+AcSquTBJUhXXdZuZgmGaOS1IfdNOTJItTrEc78r1Xz3tbzt/k/aYSAlRSH
r7tH7e8kQTb/XHs2IalaIa0qZvqzkZfIn4JV+wGDJM+DYHY2l/Y70DBfjzjdKPUaeDo5NMGrV55B
vXMeDSHzEDZuXdIAaG498uTKkBLsq1DWpEgh1hqpPbSovvwYXZQPBYxcKJsTkI3eEP2xrbbElO1k
4W/4RTHz9vXksu6dqF+jELdgSfIo2NosCVwpDtKK8ULYRWcjsdBYY4NTbNpGjWm5wpNKIDUDBUpY
k39bcCEfyzJJk0LYDEB+ls32BaywZLd8cq/PLa5lcedd7LiTkE4LoM4x5aj9c3gGhwYcgCfEkVf1
casa/KEiDhlUTcfIZ7ucYtYMHyrwgxd1CIP38At2M2o/ecHhvFvM1dQgV8gCs3YQOUB/haOB88sn
AX7WiT4E7T5Kg7WUn0iL9Ue13J6EZOL3SvveKkezOrIktgpcnhtTY18GSNLaN3Ltdjt7/Vx3AxAg
k7EB6B5KFNwisfmFWVyT4mvr8E1ewmCphPdHSZz7USjWi/4zslRuzXKCMW5zfKKy80cKvTk6QYPS
1BokRFfqFfJd5tyBWpSeNbWUhQtTSClHKsYPuhKzIpldf7mXIaEi7OTcfzYwnRX/TTmOScgG9Wnb
EUISvMsYmF4Vc2sZFNYEvVoNEppw6yMLtwhVWMVsTiXM+H09NyscMSyIMCX+XBRpbplnsZL2QlVC
eE2VQFggfI9IhmuOrY6E+sxTmoY+0vao0MTgWAi9f8FqpYU7TeZoVUJ+jHzxdgtNivRK1h0U63UB
qlDNmZrhLw4NxZeLlBNq3qfx26b2NpVgHvJCjEs1Xi4xMU+cVAHhkcVuZI4Hw5QxA9DUIU/Eimds
J7v5dIDQ5ihGMRLmfzkyALZ1/Lrh256pU9L6SO3gyVQlTEGnoZ8qA6Q15Y90hwmkBx6BrcHM5CTk
vSzqAKVpw9khll1Gg/aMlG6MOedePg2FqR6euGYp6Oj0/IWhXmyv9MemumpGhd+L+tGsQGe/M15n
pxJwLQeHHteic2IZ8D4lTrUcOcWWHXXmsD39c30/VDItRPcKh2n/sqyhPymQ6LgUqOycCa/fAiCS
pBy7B4IWGm0QpYMTp99MZPr6grEOFTyLTS3NNgV17oKnyAmG60O2g7pCXDVq+OTuILblFmUqtfE3
ZRJs8cFmBSMqM7812BeW9k1kBIRZ++pan8PlA58j1byegVVkJFLwL0eXU56jgRGS9izTjHQ+Rhvf
ZwhOjjB0RW/8FVvNXiArStSnKfZd498mv7VqtInG3tUcVUAMhtFNy14s73HtdteX4EDIcsNdVI1v
f1Mnfv0dGo0SYBqKWqAekqqdrdbDIfcqp526UZJ3255buSIBO2MqLrb+NdWR8WxVGmxF1bdEWlKK
vF4XKeoN0uTUwueMWsU+LEOJngTdXneKx9687GnyF2RgWOtm78KGzI21JzMdAHDx9Q9DMWDtQF/l
nro9tO1bvMvWajX6dsHT7V/z0zmUwb+GoG3+iqkR+6inF4XVMRvtBbQOyO8Y7qBZffz7cPTpXO8o
Oirvhx2om3V2LQIwBsLLIWODsTPJPy8+Hl630Y49qQumjck9ChJC4k7hZbF5OSOV6M8QdcCWb89h
SOQEXfBOLxmDBz5VnlYiKCT/n9F35RrgjZ2NjH4kSI/0yujsY2IwmZhKax83SLNKWtJFd2e1/Rj1
m168qOrj8EsHRUN+AZB52ut9QsMpH1mH25tEfHfPSXRCMOhDp6PEIMldUNgL/6dkUC+dCGeEbohf
XAtIjfh7Ehd02XxxD71gVEbs897sI1Hd5CZBXvCUdlLh/IX5Oe6l6H+7CNleuacdz60jDbRY+dMD
/oD6dpLqficRoBmuqSYXSpxecHOIZkttNrBzDwbdNN5dpos9NfRlCL9csl5iRMueRiFo/8+8zxcv
Nbq8/r+BTKq2ZnAmAOLM89k8BHXUDKUKTpJcQinF2F7r4YqqRj2PRtgGIx+4NWx7IsphYJtpsfpk
YTLBMRao+Z+n/vmMgN6BL7+5KxuR93fxdCWS8PhI5uLhpfDFFjqPl+XQlpBPGK/jH1/pD+uyE7wF
7YhL9T5aFZ4G7bmE/qmOOJUT4dWA+nilHgytZMdPMJzWNu+drAs1fLVJO5zgbN3OV1sfFKTCsSPl
IAxUIUS6Sazd6OQbsKuGlt+d4563sW51YMHdV1j1TPjAUxol9DAzglC/JG307aewGlJARgU99v1E
XSSlagEdUuFaPjpHM0lYQ+WfhO4iUjCgDjLLqXkszeMzus4f2ZeJ+HkTBpIHIoFutIgMBiY7hEaG
4OtYSm2usvEWGbbm4+KVdg1Q1/OJDeExjjIpVsLC08SrbF6e+gWPnnTCuoZqdyxt6L9wOKi9fMg+
xyEBemDtqzGurj4gPYdBfW8tbf8BMDS26kbVDe+7Kfg/j1txfQeUHoro0bqOi63qe1ep7CNfU6QH
D3QE876IA8ByzT6eMV2zb283DmbdbsjXq3hfiKYKsSC+KyBUkH2PyzZHjaZi3ec3SHgNQMo8MACr
3GgC0hGPs9Zp/c57k0ZmoFxG1Nz2JBcZ2GBiUM86hOmZmlCTbg0mx2gsTMDSxl9oO4QltcIEPz7c
jFxVuWvH9O+FwJcH6KwH8FSTb+zsSC+R+ptJGXgIfpBr0Y+tyVr2FbQ5H6GNI7jKvAdwoM7/3c78
KtvWNZigyRpiEJYAM8r5eaKFNDg2lBdJ7FmpT1esF/iknHWz7AHG1xt1nQJKJFG3bGyo3v+ACISJ
uR8VLM5EsMp+KZubGXTvm3dilEunteP1wBSjXQIYArTOWA0wt2fRZgU5DPZxpQcD0P/dbVXWDnlO
1upAYst4xXWBboq61VQyiMni8yUd8oOuqd0CSCA+opdqtJoH91TglZ9J4rZt5giSSLNljCblkzD8
eoorolM6xZL7cxv2lplAzowh0zssLiPv9imTsrx4VoG1k3il5O2DpG+4kVrNeN/OUBxnbN+gr+/I
8uXEXCPDmvvHd8Nia4LQ7Q7sVXzOrk/2UUJbB5QRBthb+PZtNirhLXQSw1zNwajiY0w+3tsHeaEW
CyMwmEnB+Fc/HKc8SLKt3EA4BZlIEzLT6ObOrzhsaNJiVgTfveE0GkG8lGAFJkml1twldcKPA96o
MU2Pofsa53inMpMZ8Rty8KSpeFFtxP4AMh3cCu/hlZJ++L1jffWZd07gV8tNe9bpFzbBPWnBRE+O
N6OZ06/N53Dpe7rMfCQ1geQVB+BHtRftJb8q8qTvNkxQG4eHUcBBw0fAikqgAH4Zg4CpMuIEB/AL
vWsbMx+CrE40vi/2U+Ijr8oApfEPPJTvbjaldutIaOTpYTjqkUxc05KBb/Gm19Zd7fI/Q3ZV/DSS
KSC/aS89d0iW2bRBX0WQLgWztTpila0Vye6T1K/DfzVkGsermhiAjkzXFanvgOXxpXGy7E+IF8eS
J8QywEHVjrV3/wwLv27Pi6yBpbVsP5T35I+JSStMj8cntNcc3rZ/2koIamn4Lq6/Z6gtHYjwrEaq
6RBFJv2mVVwFyjsBt+dcIt6ws1eRCFAATjdowcnkuD3+bP1ZdQ7O66oysNEObp5exbcPTQysGBYX
zClL0ZCCGhdul71YhpNZtZShozqaBkRggolvfSjqAicLjWvijHOzakcTVpdfgVfGx7R9HnZJr2hc
cZFk1MWE4gdvN58HRmd/5cm9+TRTZZ6vswBMrr/Y5rVmyBO37ZhqUL/2ZbEZQmiYNOa+EQop0BIH
3ucMvOn+3wpnKzswCd/7Q0AbsPgitLNJkrgWAFeMOLyXQnthsmKTyso73alvz+CT5Ke3rRmA1nI7
WCmHLqgZcr4qUG9Qi+xq8YDouvjtn72Hb37GbDOwUyH3uaRfSDR0R9KFS2UqHZvIJ9PJnHs59fLC
7CX9XkyXJCc000SIRuXQ/HR0gqnV/jUULcF4m+OCnydxcSzM13jm88PqYPMXdsqNeKuuP/xorN0G
cuOOzYjZpuJoXV+On4RiUkE9rTjzUodpCM9fUUcdfoT++TUVTFs6vYap6amsewMMVzqqmSsnMUvb
d9JcPoWz3FCjctY4z327Z2zSGY/3+XBKjwTDEADKvOC477+5rXlU3EIfyeIWtRdm0hhsPAescjQq
b2pLuWbo4+BdsVeshrr8exmW/WSLxswG3bP9M6LQb6Nn+UJAiUaTAWweplR3yZ/uMkogHQdL9nwD
HjdsMCltTsvkq3krFRnlMMVULMSRsqopHKFJ6IUXKmgmnjKH878frCnusy91aanFGOYaQEcXM6Hp
FpKb/8TM9YYMsgW2LyYeamJDFrtJjco43jMDOyTgh+Sd+6+xG8Q9olmTK+47PvJ+qgKHEHazEXGs
i1lvLy9F6fJH2+WxmaVGM53EulYO5vLF0laK0BvJPv/jCh5kXFL00Mka9+mzRbP1nxEgp+L5M3bI
tFVRp8DnuMxDQmDf19EEf9nwLWtoLhbmTsGofysAYxJ6iJxxlXcljwl7dRRdC7v1aB5ZTCSeKn6Y
aTXmTNj8gnrKQRVxzuhfI3oH8/cNWgEUugLoqFqjz9XI7R+JX7M3JLl7Q45RXKeOQY4+1wYV5+ne
zVlbYPzHrjrikeisOML44ncj501Y49kVHrOOeXQiWQTciypKtS7DKWHhStmrUUSETdXV58Z7u3PS
O94WVlRK8TUljduk8nivqO0bpd/dkTEtf4yWARVxKNYOzMLo7cN9ZPgRQ0QCY1RNpRnpgrhMKuI4
R++rTxGV0zt3v2POrqhy/gtIKlhEdZl3/50zWbKHEUiwqeAht8FzZk4lS72ShYzoUNE8tJI3M1br
5HlEp+zqB9SurToQSCDort69+ifSBHnz5D8X06j6E6TzvxWTfMIUhjZbw/jxDLacqWNdWnuChSC3
lDTR4dOhkbrKkI0fcpPA2YEAqOIoRzcP7YlXhDKvctI8tg5nuRlOSdMS5mAZ3HNw64sqveyiEg/N
MUEMotjDzVRTT2N1ijPVXMl0y6GuuL17TLSA0toDKAyqj0T0ohbMeOGmEnpWSKPyLTgJJTo7PuYE
dwmG+OAGMbHT4+hrn2rmwKbRsyTqfGYuM9+McP6yPxhkKGtJ5k4kSPVTUZcB+Ee5y5NlOoVOaLPr
pn9P1pB55IL3HwH6JKASnS2Lp4hKPIcUEPrz8knnb4kG+YY0hKQS7MRiox/Dz87typJ2m5bL8ISZ
K1sUo/4NxfPe+/ZIC7VnbhtqfXcrw+xnltU6lKcTeTFNsRY/6Iz4AMX3E2K96DQvJt1ZrCjaovXk
K9PxFSIKLcBM+D+5Mvgt6xEqG441lRw7ULfZyEd3gngVUG32L9Puzxu7fWEraC5WEDPwF0ilkl1C
tVnCu5prPdGojeleQ+s59KYd38fephpViXZqvxzxHsawaIHEmetUbDP4pcPbXY6NJRyL9i3DEZeA
xpvP3Eb+8yuF7dsIEw9ETn9McMsAuUvdexM2fWyjTx31XEV50xH7UFesgfCt2qteH3y3n4ZFpMzi
9l9Um6fWEwCVbhCdHswBK3r6tGsEYDutOOmrkI20+FtBERi5BAnH++HT0IGKtRR+vUaG5JS+bIRG
VJphHjVl+aDHN4t9GTjhxaAtSBnqnv9qa+cAyxUIG+fgeKLzA2wikIpVsD84eivdQIdBA0NbG41d
3Ppoi8wqyKLnyySLE/DvtObIm1XC8nxr/hgVZXSytYrJ6AHxoHF7REOAoU3WIekoS6TKjvKuZmlO
32ns45UOHYGFn7fhgDiPTIt1sjprJWWXUfNUA7PcZyl8ippqOegFs1hbRCwFyGgndq6yveVen4Xj
44SSViz1kkIO76JSRInvVasat2jG//flaYfnwmtWkUnGHVwBtPwxy+tmwzf87qnGaYUAEuK+ranE
qGhP3wV5f42eP/6AWIaTIO2PUXJdpsoEgPMRpye3gy3bJo8wOtUJwZIIxd8zcBfkGEzZU4TCJDgI
3vrcwC5SWH3BJ3IJALusdV0ESAzxQ5qg2dToE2xZsIiOjXZuR+R/lBuWU+JIHm2cArUp4Bgoz2L+
C8S5LnY5fK8nJzvPPss8dXst3XA9XMY+viGyMndC40Ld7srgOGSeKDunAnaY+PnewoTPr2xYnVyQ
yrViDPodPsFtrm4xVvvMt2CBNQnoOmxGDQuS21gEaV9DMi9N9jjjKYtPs6oXoC8shplyI7IhGzEx
QJwVdr1HEpUgDrYBjgWJ+O1FMENpNrWNBlbN0M/bOWSnpSVoeNQ7zj4kJb7OWH4j6hoaC582o9jf
GGvWePevEi635OFxH75HV2R+Czk3o9sp5xZEbiisdvzEcUXGUMBbEpccs1/OTfzVpXepGes8wZHo
HLo88nzJ617i1shWOQAjYoX/l0C7J/+LievYaluMMybBnJk3n9enm8CyBBPLL0jjGmzAWdYgxkFD
W/r1PlmhAOf2R84G3RMRekXvWp7xtvR2bZplT1V8Skq51JzVQAL290/rqUu/GWKglPYokgCZAGL4
xrIKuRMFu1mxNPqLeC0VVZyO4XEvIOyaEAZGyVlfKj5cKEI2b6I1vtaabutnsG5EbyM+9PHNnkIU
piQAGaA4fz4ODT4S0EU+oZaIm2Tr3qchFvNAJ8fLvGIcccRvlttwAme5pgmz3SC9aju4XHnZpEWQ
iOAIsA9Yfx1dIrxqAJ4hejOyktdpz5jaVSQkripRujG7JB4YxsJI4L/HyoSDWiphZzb2qqf12XtC
Z598M+66OhBQwjVmj2d7aTT8xoomxckrnvShWKpowr6sHau3aRH4Hu2bUY3k70jOruDBH8rPbiRp
kjaAKHhzy7u6/XC8UX3lSdCUaAHn0Aim7H468xvyovzc2Mk+kDE8oMcKP6G1dFKLDUacQ/mUovyE
lWUTjf7RQf8p0FG38VPkrTexT66TsVKkc4OCfldJF0IoSp8zi8q8S0vWM4qNTBhmjLcOSF5NQl1Z
jlmO455pHysj2Jp1q7YFHZtAiJaW3y0SCUyou8kaEqrGhLE6cih0ZeTVMH2HdlON5SfEnl6M/tXx
omwF7iHSwM4Ucjmx1/N20j0ZxqbLlY79nFjrhwa/HbC0a1sofNzK0uMtWNOW8zUDEsGwKiH/5Lx3
Jjoiqk/aQXI/+pNHUvO1fgn9mnomLUQrTE0VmfU6g/+VEG8L3HW73BoCv6RgsGKWzQ/547nNHvuX
5mu3gfxperCJSM6MoMCnHuy/2kVJAYf7S6kCt2zYAa+nDlfTRUPDgbAIXhqFfn91JS2Ni8XMw2sh
eYymaN0tzbI7tLLTST1coZlhoR8QtOFYIUrd5XzYyawFKPdICtUKhVXrH3qtmKl8SfWWvp3BaS1c
wI6o2zbwfCMwJ1sCaLHGJLqyJY79TVVUivbyLqePBxKMNZuL5ZkFpSSiG0+8W79JJ9Jh7NgiDWtW
PokHG05EG9G1AYvPpKCnoigtE7pYRmLyfrefOrEzKWChpKrKzUt0i2XfyXzHfjjPYwjqiaqWLL+r
qTKMyJgGvuS5V8HSMrD6JY3HCh6agx0IySdedIoFPlYUVdHCME+aI3nZHN2ki+Rs6vBdOcXtqw1V
OPrt3bDQC9Sr9r7MhA1m8PRdw8ccypI0i6QnA111d2xno4nM8ME52qfO3iUGmiC1CcdCKS1qEwH8
06lOpyKfBlDlJ7HgvCpWSmPdY3hJZ5z/9a0z+I2x0CUV2X3ExSR9Y9Tzr/M6zzI+RfMTAC9ue+Ad
la9I1+XCbYxHyZX5xt2HYcK2px9FwC/cJDYhoLu7icvZEGPpADTi8BRsbAHTcNCDAUBImeEWelB0
zLcF0xPZjD9ag2oEwhviLyS6edhos6MCtx1UTxPjie6ToHDIzZipnhhmiI+n3wmbxQQ25tYNmBn7
6R187zzkXUs0lABcOMiH8joPSQjsiCzLt/WffQU6l7YC4hnMbwBhIi0MCnFuUXM1vazsfMaKQiP9
34vl+Vo5GA2UwNGC9yr40U8PlXoopc03GnCbj2CtpgmZ0cTsBr4H972Y2AOlTr6DmRqTGWLfet16
eBDv6DTXCpxTGBJpidfEYoVY9ysKzRTpYLSap10woEpn1weh7LYHjPZ7kiMy34Hw58Ed2Ms4sV47
RIEjxwWdxbL/KMDaHzbjHcUhvgemQhpBOFRBFBD61qm4cjGtCg5fA3X+uLYVHezMZC4HliX5cOHl
NQW+qjriBNRntXb6NQepIuVY8tXaaYm9rJkFXQjsDY/9dRpJKEzkukrjqVUs2g3OcpHeJh8YUPdH
U7F82B05WT5LK28MQV3BfGspiJzGfYTLy2JuLGQbp+f/LWMw2XvuQQklIzybyrOnoTZChbcKWtbU
BEAG8NKubs8nG5ycd8IvkfVwydNUdF1+16mLG3v8e68tNL0iilgATzeqOVVlBXTth0Jo7Q2izPmV
W/OIVwThJx9fvIq6LEYu6Qu6qN6bJpCAEEPHj95yQUOkEQp/TbHFrC2ja2QGGqpbZMbtUo0p2OAQ
7N0XeV8wNK55OE20BY5+7EGzOyBMO2rjBS/7ksL2x+JBaLk5m9ZURBNxNdDxG99x+FqNA+xL4wRN
mrARlSeWJ5z0mvvgxq0ROVMza1zMig4mnFbKRIxJhlpJ0nlmf8kKObDi/7mDMBEuNhvOtKnKg8tq
rxnlQ9n9EvgqFTwf3p0CPrUPsTcMDnhbh01nUJWSgl8Ew8HXHb3SasIwkYlGaf9ctdXnjtc1Blwi
MNjcmUXk3nhGB69IAt2h6JIYxnLuXmt36E+r8ajYWUP/hxRK/HMX9CVPctrDBtrQPS44qO/29hxo
m4QqqWUCLbfV8rT+Ibx9PGgQVm+JzwGSfjykAIelbVeWN3NL0f4lm7p6mCpLHyjS3XyS7BceElg2
VSu/Pfd3WxedT7/H/72HsEr0CA5/3MOcH7bfT8mTJmHjUB/n9VnEXu8BPBrZtdLX9oB3hjERIjfp
wie/kfEWDPb7PFEoQSr/ENjj352JPsKNgO4TrxiTUhctEG4Zr/GSOZCYrUJAE41eR0NRSoG6OG7R
HB2jrjMY3iVn9dGXousvQuF9+oF94Q3pTPpm8HyhNSG4rTF0xKgeISFEVgNinU52GCEg8e+5fs92
XUORt4LgZRKHK2q3Bbuk5gsbdA32yt60XPIBydjTRPIhgr5k1HlOL+x52hv9CYMFNd7+R8YiMsvZ
82DyvMWCbhPp4a1yOKgLYglufU2DmxOrBCOZM0IrNHW+K+DYnlZOytMP0yJesL2i0DNkrMTF1OTx
xejYkJgwtloAgbiI22I5dzlvnjlfNgdYqYMqKjyf0Dc+9VClYDo07R8oh4R0Coky2IrK/+947TAo
u2iA811cNm5L1aFn24oar/yjSTJUIDZuzg3eLX44SI4A+frI6+djRb7gMpz2hs12e68LDrwvjP5S
8TzP5CglNNQ0qStkJ0SquvDJnC+1XglKY5lMnowLDfM2gQcG3aQVPSgUruBp0Qi5iReG+Puak2+4
ipW+Nyr3xTWckVJiUF10uLqHignB/njca5wYx/eD6rzwfwVQzG4aziUagUraq4PoCWVpa+38zXPU
o4OTM6IJNKEoBQHY5kFV7D9uN9d80iI/K5IV8ncpXaG6UWZ/GKcpso1lOk89dxx5plWV48dgLmbz
3zyoPI1ZTtYpDAeuP772GWkWOtkbh3s6Hi434jiMICOlqF3LWkLY4FdPl+Mt3dr8+8NZvesGNtUJ
g/m1FqF+BN+wo062BSwSEfbqXaR/M2ytHq3uq39iktyCtDHfy7RiIuIMfbSTIFC1FukjS0mYtv8q
VilLk6JPPwGxqzginnfwd4t4bc5mlN8kqZSunPyO/QZs2ZQUlDy1NP0GcDguty/6dFMNSll1+aVc
0mmAmRzcYRgQonb6WdvhvtwIOoOhj6ec5faK0kt3lhEsLj9HNSTQAm2aEgswbbkJ68mKeqHSJ/Q3
Ugh/7cB5mvuRnBXyDYNt6ZZRhmiD2rI5MhH+iWGkSO99BhYZYdZtIIq8tUmyypbbyOIrqA10owEO
DHJ14F+Sx4JPmiJOhlMo8i4BnGqxCZOjaaKDmKKglvbcfOq3vRNFENidmQY/ZxbbSizxU5xpLWgX
8QwmzfFBfh0pS265K4rZ8qFzPXnHJHIPvzhqkc4Sverjr/shudMNUG9SywjCHLO69p0F6c/jhvms
0Tr+b6FQqop3RWCd9OzfCIQiLpRDfffGW+Xar0B4crOEBbn/5cwwlIl30WN1FK1XuQtQ2S7u8U+i
uRKTAApO4+0exgd7Ug/PVVDTkE3KS6uLP4Z9w2FVUt3m/TB6ZmI2t+RaWKzIyE0H/YZMlgK2ufsR
spS2Si29HwW686Kydj3JrrnFG5PqfsFKBvXmPTGfeh1jSUfSW6x9QA1Q/gITY3r4WD38EyGCldpY
gatiTL9J/3xv3dM64DT2g0ruqoxDsDRr22aSUIs9MAPsKtBj3N4Iilfwhe01aO9JZnM4QNCK82mT
+4BcF5bMCDILokVQhkY8rDvQXc/qUVUzyzEJ1kBAZQlrMgzbZaBZNC7R3/Hbz2m0/153Ctz8P/KR
zbJKDkNSQhQi2taX+p8Wwi8cS3jx80kELgJDRgn2t21hgupc41akSAzItzaylM9NbgD/S8gcSTX+
FbLFwKvU+Ymct+qOveC3I2LtZ7mszozKbRdgSOKZri6EWyPkWYswE3Gd1bNiNkhaTSavc1LEAsCR
xMNOE6ZIWEcrQgGaTrzMOiNxYvA92TK2jNzFC+gP9UTyRcNRi5201nFCnBG0dmevG8tkqggTm0BF
rseJ++ZGPfI7tSknrpOK5i5wtdTQGTLIZLvQX7SQ+ptTA/yvR+GVXmkswItmekf6rh8SK2hBQsG1
tp7SUSixVUu9gI05AaZ8HnAFdFk65jrFhzFCa4H5ct0nHI9vCJ9L6w+nWBhoaThYv6UFuCU3OQ34
w2cj+tusXSvnP6CDeg1k/FZRHI8zcUDDuogr6pXsDXROwEZJRlwwDY+cL0CJLb6+2bJMT8UH17lG
XQF1KwvE4b2NhH6YqkKglbWSIzpwkCL+ZrMDtj0lAO2cEcc2aEZWO3jpTk7921xwYO958V00idHX
zVFnsieT5YU5TxCU9ugF73tko6WG9SpxHYUlKksGue9zSGZVD/9+BTZG7EMQQHl7nzx9XPfO7jzW
ujcTyNMweVBm6nRqOLVv4to44PlC+X1UDBa/oTqzHFA1NIjKmnBUJOIoZY95ufZBhAUtjrmGYGfU
A6lKhNyHtzZ+9zNXXjoF9TdvpYg4b6B2ku0V8eZQe72kg6n9BgACmqFhjS908Oy34i5v6cZUDq2d
R0i6RSy8cx6CYzoG4mYmq6wOPugxbtXdv2wnrj7IVqUQ4Ndq0D1tPniZoz2Hhv24dbHGXpRmARW4
R5umlrXYUQ0GsKJxiUVpFAtNUlvIq3vGjPTAqEMH7rchJCIeLkYfEWNbxRT8LoCAJXfHotxBho0g
S2UlOwD62j79Tv3pDQ5ddyDX2LA92aNSg9abZGe5PJtM8IbDcohhgNLObakQ3ZFAlwTHgN7ScbPB
m8rqxeXxno1YOJhbjS0z1Er+OgOhgy0cW+2UULzCh6iKZHIf+4r/DCNL1nia3CIC4Qx+F9tO67CI
+iQXkXA+ldrA+SbHw6Zr9gwbO55H8aXLVMUUvnPvPQpS1NhTJ8dAYSFWIqmGGFA1qbbloj9oRPr0
0CEMRso51ISc1MvmtLCH9aTfec6d6gl7NxnoV6gnIkJ9n1wh+xm42puHoUp11+Z/GPE3Dhd3ITTN
IEqvmzqYUZfkNWU3WdO075PikWo+sPXJeIQmK31koQDtbfB57PFajnYNX0SFGWlEfC/KqZ1rdmjt
1MW/VvvPilFEOpphkXj0IcaLssgVnIxzEXMOKGYU74PMYcDjyHwT/h6YC7MerIAJ0Sv/u8ykjeBd
ZwxQrD42jWFlFFcf9C69YE+XKrBu8uU8LyeQ4gNNHrKRvRncVrrJYDMOXsmLvkEpumxAZzqV4ODP
YCek57F3vYvURHHnpTPInrUoLl8jGpahzwJ4ih6pOiY1hPcXZA+kE6jw6y/ejggfujHXJQea9/LB
B9c4QtXCdIt4g6dyMOuhYaH5CfAo1b0Gj/KM6NZjVicjkbr7km5hDvVkNoS5Oji4xsz4K50umbhy
NkDmD0HEK/eF/jvuioA2e9LQ8UkJ8z5d9C4eZydcJMoeD9TbhX7Ywzp/ShT+N1VL2U6YujNeqzl/
+gz6msHyHfYSNmMR519yfeYfmbW0mxhTOFLIsOnf5SGnO+YJy8Rgk4YpwrQe8XM9AfGg9gufPBow
YCAe7Rs930WB5+KC0mvnd5Y0fBKkv7f5y48lcvGmUksnKqIv1v9XJ84KfbwOMMB5PYxHTC03URza
0WFwfXWYpKaj/1kFvtj86vGQIvokUp9cyD2NEdNaOMC8JNFjKQQzrgIEsALWI5skcXkf9BhiEgnp
pSmDTZUdow0KDeT/A2y0qMPOsklQqTSq7O29ZhDzruYBAwYje5zZ7j7R+rX1Zjs+6PnFyI96eeXX
i8sOXmqYha4qpU9/eQ6Rq7EsJrfT95KJgWLPw14etQPYGFOIiglwszVPz2oxhEvNysKq7w80TUh4
goLsMHYWgIugPzJ9vowej5iP7DfYda+x7nO7igyFZqJ37GKxPyvitpjuu81r7f/FbUlERjpxYp6f
uQFnVnggnGxxAeapqWay3Gzn3asKCEs5R3Drf9Y+C/5C0e7Fz2xsOSG6ZHONpD20rX1JI+vU/DqR
kUOiEYn3vHF3KGjFqQg/C+euwD+5yq5gs11PcizRK5MdyWPHr7H1yo40Jk1fF7uBpM/+7Q5m88yc
Zox3AGSMZsWh9u9sQpbUEItxJ2eHsSBPpsyKcXN4RgrDNg2SxqXjok0DeudG9ibetk+8CZroIhvq
ZuoqjFno/U9iQzlAPax5TXZQ/0ZGKk6xQFx4QYxh/ueNfa90W9TXX6DzpmcF+P2wcS+VFWEP1H84
s71btonsDfOay0edOCyxj8fnkFACkiDglhW2Op7/5rgGUi5lmLW/Xpl6thRgONqMoEeOiUVvHjVW
fIObIgjEPqNWlOmjqSoC+mOotIyO1lfV1UDYHuRFPrwSH4YRzPbkPqwzdH+kkXEJaU4Uu+4A79OO
3m38uRBKn6H7quu8x/l6fnVtSQS0HSlVzJOZtoQbxPdW+Oku3E2q53Ucdf/iJz9WoVzYuFrWv//G
QQzZldFWZN6b48pkjFg+oYrzQjeDJ3XzkJGwN4mJDN6H52w+hKFGz9FMrVcHy20N6EUMibcMwSBY
ZPNOFoMLQqctDobB2NJ8B3sgopGB4Q33kdRTBrM/7v8D71UmlKkQRv1/u0gw05xtitu05YyeYNVb
VvM8n0ntdQzr/xTZGYveWPSOiqVXoUa3XJi4gDtoIlSB8wF6YRSW/1RP/V2z3Wv9fgNG0jd7gUDF
rvUPR8xDMdGyXBIoPyKDmbuBcJ7BUCEMO2Yjv9eQCgws6DPAh+SsVQSGitTbGVxbkjs8ppVjH/0q
eDg5UZsDFybhvUmZH+zgi7FG9EaXqGNGkdKn/wXywKftgG4DJRj3Kv3jO3NC4jnUp9fhlLKo6Avx
z/taSzSck5QQEDKptWkY7G2qUk67qRhAqqb9hb8xCylG5ChwIhyHopiaIw8S/36PQGr0pM0XHe32
Dj4FdQu5Q8Q+dygHv0om2gs/LkTCOp0jrYXQF+P/7AKUKKluJItXq4mjXXpoH1NjRyeMJ1bUUIWt
mVjUZsMxbZ4UQtLtYUCyxpMDO7o9rVLf0Tyv3FGdSh+/aD0OlIBweLKwFwsl9YkGk0WN8MiX5b8G
5FYQ+UBrcoCcerJmKw0X4i/Zfw9/m+C8VDQxMXQcTXceWFb1KybD8tfyBLhnq0t4XgFN1x9+TdKE
xDmbIK7DcRBtnEgJWxFSnNUU6Ho8SLu12XlQGw1Y5Y1zW+DcXWJ4URZ9JJ0KCruH/1BI2EnjCCe/
w9DT0pM7Ty46fVs1JsPxy6ShddQ+IXBkuIBndushJEklPqNyPntUWtqjfpsMnJZLLe+81yBRRUCY
EudkMV3Gk2QMmEhGE5DrYherW6hrGSqmTuhlW4bUEp31GAI/5oq2vGuVp7xEllyurpk8jStdK5sC
n3GVJSJryfl+SxJcBcW0pF1ULcOR5JeDynIaiyo7Oufqsgf+N2bIjw4ycCJGpZ3r2j4v7TuqFPjP
ZEqOBk+wzQbYAX0EAx1BGXppPRU7KZloq/w4Ld8DImwI2OBEWr4Gxv0uJpmZp2t/d7ryWItM/9j2
HIfy9inZTdQrpI3fj2dtei3gKkDnY++Yspj1dAQ8J2V3AS6zgfDa5QYid8PHp6gS+cotbLyli5Ob
Ajc84sJ4tECSL3lSqD5z7zIcd0obtF5j92JbBXQ5+2a+DpY0fiIu9PHNCGSX7f/Ukcyotlz/K0Ql
AQ0ouWjW1OOPzotEPZ8UlrvxqFv7TiqqVPmh2HOxUFcyVQgh8BgcNfhUvRSinVDVMWUBoMeiFbD2
he0wcbt2QJWZDoutGzHjMwjIaEMcN6f7HVdRZsHL8jltvXkuDqvJ2wdOQp+lAOsfCmv1rXdsjEju
vi11hNycuGEjio1xd+IgR0kH6Q2jNg88Q5am5axURLzJj8lOI3cl7AHhT7Ry+3yatCX5QHw/trvq
GiPtCUrx419HLwTEg2cllJdq9Hd3iqtth/IWvtGRYoOtmCSmlYah76GPWzJzu2vdiE7jXftYRJ/V
duSnR74oj2IxjIy9trbF8+N3z+eQpvqomR1dU93U2rg8eSim8kizbw6CH84iluCBp3colZniRaXc
uuJhFzc31pra2SjqloKxM/ekwIh8Y2HtPwbVhnIwV2K1w78hGgZb+owXov8OQsw0jg1Odj27taLw
vIufbbpzzeNdaElUqbpqmG8On2TTKj2U5z6sL5bohIKFAK153XF/qRODi7It3FAGRU6iDBtADXsV
g5UYsdI9b9RIXA+QP3GfoIUzszqAgYLtTUUliGMwiLJ585ZotRrenEHIdB7u+bv057u79OE1Qwpb
2Yy7zej3iMIpTrHcqmVUBGh48o8ze2M1vbi16rZsaP/mv8M+fCkIRjBGXvtl/2MvD9vxtwjwfCOK
9cM+EHmLYhmvm8+lM2wAGHZzfVUemdCA+xNMbFNdQSl0DXWEszcWSkt2jgIs6YJCfar3CBlqa1pF
BrA0Jysxi7mFxNuaAQEEvbgBcKJwAimIPNcuIeFoFZjLszF8oNOLrhoNJ4uRg21iE765gm4/7+2v
PdD0YbmWR81PoYjIs1Z7bhh3df5xah0fMycWqN3dVJ+vEQZ6TqgsY5gV6hO1GrvtMNT8rtpDHiiO
0/b9WSuaa0U8KCvOvCKzGpFzkppVsnQQygGh6vxyJBWx7vRgG/SouGaJOWVqhH+h9dyp8DoBcx/U
Ho2E+JWFBeOJ4QWxXGraxhfmZQd+Q+cIsP+LzfW1wL2dEBD+BsSZGAiX8aTvrs+7xMWxqK/GLBru
hEhBZOMps+Ab7msyTml6XtvmmBmtoNaWRxaB4gi8uMKhNHofKMRL3IKfz2yeD/91JWbNmXKYSFCy
7Qp7uf1MVvIUGvxWie+OG26/vnh3dEXLbbSrL85cP3vmiRf1YoOcY2o57WBneBc9jRLNdfEYj30k
0jK2b/NzQsQ3D7GLlLA2s9/LiQQjTI4LP2xylGEOqAKufU8dPUBmDu8LoAIC06dFYkv8ZeDITopL
PXrAObA6dmF8jcavdJgcqRj/j1qmpjQGqDsdc5WgB5SvVcBjqXsXRiOvsAThHPlRbOt3mDQ6RoTW
JOEQ+CgAwFv+UY4kENNJFHIJ4oPZPu8T3Z5ERqdSaVSfkTowvEWwIQugDQhCxyFIXOIkQdPt7ZNu
v1xVf7/CCq2PBprSZjjrGbW7/izeaaQrTgc4pInaiyK5vYSfcVk1HbD1MnP0PpzZ753PRXvwjSev
h6iD7DpZi1qGUNFkXA5MLpQu3EKwOfA8tCK7GGY5Ly8pQadxGYTaTKvrYHcYFsDc0c/o7V2GmUja
nqqigQw7a3XUmKMf2aojcYBZMKT7QAgr6bHaVek046iJQQveMErFdXtEUwm97zPKi7aJRu7A3CCE
mDdc/TZuiAMelhKMHJxW1MfFWsGs8aib1Z7IVu9v8xH0Bep6fxfVuJq4gDAnxKzBF9OXVw0LA+PQ
WNQFzRSj5G/SRVvO/5XQ0iHlpigGxfuA4bQUrWMlzmmlVqECzUcYtG9GchWfUDoVu8788RvXjDB2
S6+MT1RnvfmSyMdbcj4LTxcGsjutXjO6/dZ/AVFai6uocvBs+4PyORrBISSWiVs7CoBD0/9tfYnC
zxqRn+Sw2P//okAJe95rGciJ3Dbov2+oafgn1IebkULkKljJWCZ42Qf+2N+itgjwB2TNKHDNqbMk
VTlTI/aFZjNB6P8hsd9adsapPk8E9XgHCgS9yM5ud0RvhzIsDKR2j4xPmOE+pS+bNIXTZBncQfmy
MjUAYUF3Q77sDaDDORE5/ybjW6Ca/Jm/QDh8wjICNcICYkgrab+Cs6LpGxV94Vbs2Ejt/zXjoSeS
ycmk9HfpANrKqsgbJ7vrvqjtf72FHteMzBwwU0Kri8bYSsnQ5F/746sN9kuqWoZgcIHqFG1ZK6rH
8mx0rDgKGZWBJf2EfaOTmwTke32oCacC2gWRWlQZ7+FCI65lTAb6KKNuSlFufielPbVXZMa6ys1I
QwBnIisnNDRIOLrXxmN1go2vv0hi8yQC+gMMhBs/6U2KjWT5wxOcVsSYxTJNLLpgIUhJsHJ8DtuH
nIkeejTi8erQqMhZqoLVsTM5WT99zDtHRaN1sbX5sBWHXWd2chIR46QwUovIlOgHgSctaoYWUH9S
a3RUd2kudjhCIk3D26s9qcL4K/U0bOYdW3+pR0OlW+gZHPMwl0qclQTeGREhds8YSD0usEjW+BXT
r2vIaXO+/6igxksRaAzJhlKMp6o01dboqoZF5NNFbQ1Raj2o5K8yfe5vmFdlJG7bmuCUhJRPXL+M
7z43LhwUPkow4QSTmqPSAtzCCMHW2E7Kb5sFrPeblUuBHys+LnUl5/hSqlrALn+nswky+vVi28pL
mBdBW9ztEV8g9tuYbhjHm7vseb/LPGxXRrh4GFIu4FbVdeNMLO+i97kLgODWI9YKXEM1sQCSk4cF
SQJ8yl9q6x1Z0wi3CJwEv0noI4KsEdDELHQmR0WsXojtLEJp1R365Fm9xF7MBKwEh1m5dcVMm878
JT2vCUi57BwPZb84jXtXmJahjZrm2o7HNX3pyYiN5phXTFNcmoIfobkrDr6o6vu4HTIZxAoZgmAE
HRXbMk6rHVS0iHpoZkUciRiA+paLRXf9DAGcjV+5rEhk2QnNJA9cug+/vq/ROASeB6XJcWxa9bO6
M2A6ddB8PfZKGUc97ZfVhafS1nZB/YjcW3Byo+vzGMVDDuK7GsaqQ/L6yIZoqg1LDLqpB0A6w8lL
Mx5wx56uivs5C3QF6tLZwAd94+WtenhsMAsYJex+KAPP7BY5jpQdqzEsRQ16kAHpEWuJplvh69zr
plLEyw4T1INxgcbI2CQJKJ1eqLqvcwBHhbaPQrQAra4JR40q5jnLHeOU/Lhf/7Nm5Ed6Zar1/Us1
bPhzicxqUqfc23wM/Bh8rtvXO4oT/6glQ77JTFb+0ARBnNnCE6yZORPpX96d5ZTTpwiGOAkPw84a
0juFqYhLkBj9prmjm5HFtZOvxpOP44bxJ8fT7TJom4VugVozZGLYlS5OOHRBCNDs3pXyDMq2oCpr
Ys46gnC/OzLpCQaP/bCN4mkIDcEpR90f1oOFgNy9bnCm52dx6vgjTxYy1AdNatVyOp6e2dyVAgdg
M7d2+TN1Qiud+1AM4R9Q28oGW8qRXhA2tL6maTAEQVHbjieaadUBd59lcYx3OEjw1sOXXgi1zjEF
6ACIm5+HuhQcW8IMLjZCK+wotdrOt6J1HbcYNH1HCLu0PB9zhMOwaGhDyW+pRouZWv5+qovO7NfW
4/4d/Q1eFTbn3r+revR8qfWMvspSDtWyL6jisQReJF6g9qFrUGWPf1umPRh7nzGURyEd7VXyCDLw
7wZL5+GPFF7AUWf25ui2Ncmn7FyGYP5tjJle7IPy0OmUDjqYXyYRpFAcFf1jvQXMfDhBNy/t4fuq
QMmRjQvKTpyZJkWuKO+3WTqPxg0ocRhe6qXAe0ReDaASl2xtoZ1+QZ5744kYPcGL+QkoAgdZkEye
1UOdc1wv34M7RKnT778KRv9j6Tg5iHWyi0zLRW3R7FjAB83WiD2fGFC0w01on/VAqKysIUcfOkYL
UDOe8UGRfXr+uJv8FhXGeuhlO6izxm3Jp1EalyXsVFUTRWpiyq2I0xOlkflQmnt3mpftf4OxM64X
lIORKsg9ov+fnQnbEs8nOeyY2uXTO6mbmq+f/xvOEiDYOawQRaU3CjNFtp6pB5fqf8nknA0TwKQy
7WHKPWT2R6/NX+3o8z7O5KVE7zODqoxh2A2+SdivCjaXeKpbjrPO96jb2WrvTZsTUOkpCyAKqaNr
qT+7tPxDoJecPVFBjf5azwc1dpVA7IrZ97tSKbM7H2hCXYjKK9oXCTQM+guw09UtPcapZC3E5cAZ
8E60W4a2BET0gMPN6eJtL6x7MqFK82my8zGbw9dktRMJW1e0x2yZv38rqafZkSIru3U0zC0sHLUj
P0/Ryy+fQSbvII0v2y9DWLDyoWCYaYGi9v3MTRmGb6yuqNLLPwaXZuA5x78fvptgb5yOcS1pH8zr
V7tNOM0fOYcbkoNQi1wvu67ZIq2iZZP6ZwcAbiwuGfgK5iTdQTNcvRrn+WeNluHBeAYFQ2ySh8+w
gyEWDRunQzuawQfu2ei/5ycG0dDOS09tH3zgP2vcEIVL4zihNRVRtQlyQUbtG6d9czoOkHj/3R+R
hHOFS9FfocFv7vmBeAgEJP8AaabJzMOeCXlmxLKAg4nRkHf3IE9oNRm+QpIPu86W1iEKybHFvow4
Lotn8sfkyiyEo3ac55/O3rhLFGef2geOxk8S0sDsxvAnFtFjGTCrLvgGgYuASVo8cNzSY5XiM4Qa
3Goe1NjswLW8IhBaJOizvbFmU2ZiHJPJhC/haHIyRdimx2BK5Qgj/ftl7VROCCZlnmzieFh5RIMb
t6uC5ENMqjo4PUYv4J39myUJ2MvnMT10hVnO6ifI/pqLqyhHIE12jfb+SdSs0GXL8MrFw8NskVjL
GZJ70x+JbqcRcK4uU/Bkg1xBsldVG5uM8DI8tyNaQ1zW8bx6iafJkwjW/QT7nQzBuy8zLhHor6h8
sWWVYnGrdKQ0UajlWJcPK3OXXPmyNCRvy/cJnFK7DATDjOZG/QsUL09aub3AX/AP4nXfY45aHWhy
GZOCRWBzjeV2g2zCY9Kz9DeXmBIbGGynmaKznVbiDQxY1ip7JOCYzm3Nzm2amdqPSaV5NhRJKyos
aw7HxRgE3XXFXTTUej5kDeHw+5A2PIr4KEW7BS3WHRjcKFytGFH9sIJ06rYjEZL1TVvl2ZI5ESvy
AVPRS+C7+FVP37rK92hZ16D/5Nifd9Rt98nh+jNkJMLymf2EcKMMLLyJnAN4JZoxAKD4rtdMNRGe
LE2Oo5UY7dVZc8UwUj4Sd6vQm72o0EYWqYGgvXcPv2qMn0biLbMsUxWDGBhTSeROAcm5Lzzi8xOv
zmLlvFVg3xvSad4OuavwrbPlQr+UjPBtprhGWFS4ruFbtSSdePnvvPJRHl7pKr7L0qolUwdjf5wc
EQJFIICdz5/OE9fsy9s1exofb/86jw0VqBpSdsu5pOC4/s8HKvXeBV3w29cIbXROpxHroN0Li7/G
kdp6gQ+tplovFbrhaWKNyNyahbtEDxoqo5zQzT+mNo88lhKSj70krB4gRoDDHXbgI7bfuoimwA5P
wqHTFEGtYnSR4IVoiN1WTjevSLwXpOQZQhtvWOvtCZ8ejD0gojcxcoSAJHM93vZmN1RGpvL3iUoC
IML42LMKFamsryGN+cQCSACxM7RJXEc04fs6WAY5SN1ItuMrMG85rceFKSHsVjmOgp+YpnDTWOM0
ra29KQmvKRc5aZoV8XD4j0CCWoSEpwodS/1qA4af10ncbRWWV/5lRKbLqPzl0y9BtwBrl6igec1s
YGs3dVs32Vid521UXBfmVF03cow4WLSHp5JC6pWObiDkmsubgJ+ok2N5ze6+g7F+Bls6ZJKOAiQV
3+vigArqswpjQEpeD4R8NamLmZlDDYqYZQ83bMHYWCrnzMu+/X0BOz510w0h3xYyNMVQv4/HehSb
HLvs6pfMTIUWF10Zsy0s/sv0woWO8CnUC6icfb2+x2YH5CTRpnBnTvPRwqz5wfbHube+nxNv1Ik3
gfyWZafClyLoRPnfdzV+CBmYDyAGm7sm1rrQsL4rbLIhH3RoZSPEYILzkeP1KKCzqJBH2ZmDjEsj
l3ValfN8hN5sFS8/WID2wV7QqJI5ZOmwhQkUQgh0m8v3ak7mPimAIdDQSB032ztWcc3gieYK8jvR
4PF2Z9HIb/cqC/SU/5VcBOsKAZPNRhX1jY7brSrc+KypACVvp2f0FwLFPEhOFYRDPlYIO9XF0DQk
450v1Cz53besNtVnE3xL2XPltCtr3xNATVGqDyjWMgV7ee8o1i/EzMhvL/AtHNq7ODHICcBoIhWj
XW35/KAmnRaMJcC1yXAC9WitqnqdpkGEGurKLBtGPzy5ie0lEh/Z4vQcGdCdSinugmBpbX24mzIs
cV2i3AFT1TTNuwqSO5XoeWOrYKkAmy4itvXM/R4Bags5vqesSQD64FJf1FLC50dx8v2ayAATZ4Zs
RgCNe0RdDa2EooakA/1rrXCGANckg0P7H6UU3fGULmaPIWWiXFkrbbvctKboICUPxsngqNYdze1F
0Oqv+GbteAubcS361kDOGq66jdb09p7VM1SZ7viygoacLNngL6LrlzLiGTDEIrK/CftQGelYuZgH
3djax0axlIcenXjvBJbsSEj2m4lpYSeC7S38mxBPXNbz6bsXoqyKXiZYKukUWLsFvLkfGKHsuSwb
U6AkGJtVyBNwWTx/R4h5R7OyKESEFR7mBexEA0oJi8Z6yA8mDWPmmlN7qj8LBHpu33TdJ3uJQGCZ
voCu9ydLZTMxNDRsfNLH2Vd4yAXlQjxLXlIeYDHRxOzRLRO5NhLlKlTidPULwLyXR2ukX66baojd
cSkenzva4AfCEyhuImdegQ/jKSoC4pEigvwGFUIvzK043/mS+c8ft3hzggYlZgAXYZspi/iND3+H
IQH8z+D+81zPSPggk6oeczSJZn81IEe0WNGjpEe/zQTsncSdid5JIdMLb6Z7fmJt8UzZP1DNa5f0
L8w5t4mV5KF12f6EXiZs6qAkHtfTJ+K2lCmANcIMemPrBtUbRYLyDhWb9oFpV0XAxDOxuCSlUWvf
8Nv52t/OauZnEaKhhmvkMv/wAIrM3+z/84tewMXxKZ/oJkzDUe70VDkgdOdsILtWwnc8cbOJ81EE
bIp78bLT+RBb/8T13ftVXlIgiuJOKSuWQ7XCoMqaqBW6WK8UFggBQUoKDkHRAWub28XqDv1Mme66
q9yA9sp6jHQyROmYLIG+yaPXYx5BkuuGD8Elu5fliRMiJvM5xQ87npfS4cgAYEkXclnIZegrhhXF
9C7l0tOapHF8Dj828RQhX9yno8zFP5CqspcdvCzLzb7JTrY0tPDzkbgAPNk4Qmwrt4VzYquCBESs
kCyaQ2RoH02pLFyJfBdsfvCY2ywjeCxcg15P89nIzdqfndGrtISUdrg3ijRHCG/397wNsEojd1Rm
rcDUtNGoofhZZ2Yz8KODHwu6Gfeq6LQBl/bLS8BQwnXFKpSGBSDPv1smVvKKV4FAuiO0a+myvFA6
tzt/Ibj3S1mAT+0yKA8iCHBH/rWgsYMvkVdACaxgNCpxGYyRfAAW/MJEka+2EqMC82gDDMKUo57Y
lrz99bL9gBVaSMYxcc3CC/9vrNE7AT7sywYe6nvQkcUMkfcr58dWALzU8QYB32RrBSkBsaFAXKyu
hGzMVHbIwGXfCA9ijjJqrDWbeGYVExa4MvUsz/6Vnt1fSul0gRvT31tyAWDMnUSr8D4rIS6a65qQ
C0BBa+X/tqcT5yDHxxGY4kMRzaHqNAjlUl0hbV6DzP46BMbuoKhaQfgkk4ylPhC9G1+3cVTmgK4w
pnCZEz4DKSt3GLJ1g1sIU1zwY1jcsogSJT/s4YbKkOmYcdkPYKuTBK+U8mqd064Yy3NNRDjjF98g
GUsomzWeBW3+u2v/lArZNFbPSoIeWKLlwLgqVhhTh8/56O7KYGG6hwtBqcX4HoaN9cqnXJswa9Js
k/zlid3Y9TsKMsk7Kql/2O0PMMXA+BfIMWU/1eGJgtZMl+rFcoplabctfdWyGELTdsivGq784NyZ
NtihdWlrDdTgFfX4li/ei4edIaodaRv50pOVTswEk9Q/pBX3Dog93ybFWjazjhKwhlKvdkLQFY2R
ucfycJxjxfh9R0VpCLySAfZ0Zz8IWjMtfcLPcQu98+K6pgtKKNnmjXUlJPDHklubimLl9eXBqWrn
YuMVV3Q8wPqNJw9CmvkQUVPd6KmxeS1VR1r5t30k9hLHuwdjSt1/htkNjmIrPkUOQhAsBkMT9E/s
sU/BM+zVd0UPT/pAxKd6e/tTh8Aef91mdRXs6hHNAe3Fr2tk9PqnIaHsVQrwOdhUJuKXMmJUbbcl
i4wnLeiA2kJfVAMXd6XeQ6xPXVHlu8QQn7i2N2tOOIfZUei0Ui8jQzWnaX0SflAw52swPoC7Y7rh
QLZfSkvxcbJG1WhzNdqJIlQJzbCw6D2jxy2k0w8KecfN/tMkTphqjmk5FHZc/n0A/c12tEW2O0IT
DUoErCz0xlqzAp+67uVZbSuAZ6m0s04FRTmULj/t/0aDhzARMCr2GR17LbkNLkoEV1217gu4aXtK
4Uyvhmz2t+4R/ct+n4oUk1nNzu5HwCDHvad93+vFti6Ngui7MuLgrXeKHvPK627TtRRN1syNuzE5
nxqQcXCgk51TPbCsin6Wez2KAT+g+EQJan08lbyKDiKk4GdcGDeD6rM6i8/rZDTNt2ye1iCtC2uQ
+4EPaxWLRP4wT0CtiEADVbzayLnBKdz8qiWZ2TL92mPq3tdH/taq4HvszlAjFeXy1jTu7WvebbW5
uSyxtiJ/1pa0f8qEI6BmmaSXykOnbUAq1rI7YKC3fa6q3d9/+NxydfQb/K8WUKpvCRl2P6ZKmmK/
oDX4yl0OFhjRUFO2M5rhUqlWfrEzONzdBYDEVZyKSg/imXIWz/PA+7zNbYfnMPcOybRRcz2JeQ/A
DCO5u/z627gMmfZ8l1B18AmbAWvIA+Z8xC7IyrNl83Bzs2VnxiZkNI2S8Kq2i0ebyr8vrcIziV7W
qJl67f3gJjku7lw11OZSPgURXlLl3xRUgQiWWUjvbiNvTeDb9y6OvXPdRYZdPRm/n/1OpmbObH6f
0cuBGNt/wi9TMotiUtinQe9u1Gym+c2+wAWVz8O4FJrUa2+Cg4Jgb93Ng0415cjyQ1OFCpkls+4e
pf0G8lrRWVxWp96NuK181Z+1odm/eDRR+pm32Gc1EVsr4omikf1kiZSI5egGmP0Ofd8CsufrAT89
L4Gc2VSmtVragAdWfbBgW1jeeBKRPwizu6wDhFQzt5HJxjGTyo8aD8qcK17yLPrDeeh0haUhKGCx
gjY3+n8pzUOzkIp0gfgGWPTa8lByHJ4DWwec1BGp34hTtcWblT50+62lLJfb1K8aEoA/wTOnXEPX
ZrwenJ22m6vf4Vo+aon7oGbq73UUTF1QcGlkd/p5iNn+xpAmdN+xO89YP/gr+Hvqaaha67W8l8lN
kc+OYtWkAI61ReqM/CATqejNHsnNEchB8CfoELei5LpSoGRDNMkz5o0kTkM2y/y9vGe+rtEhCHSz
cdHEV1/CSTPSWKjlO2BD5nC3pg+52wtNIc0VNv8n1VMfyqh6J+m1VzJc4Mh8yLZmkv0NOIbELdpi
FqiRm2MVwHCZU8KsOb03nNkYSxZ/MrbhgObOCAkKblHPnNCQkh42Z/Km5dv6APOVxTZEekO4HHQ7
FQouwnw0a4E3f/lrSL7YbRk3jIeEy4MIXOZRIwqy6+er4jWT8Szy1bQwXN5F6kyV6YU1vT8Ozvz5
2QthTY7Xoh7TLdKt6ggEEdNzDoa33CaFmsbinzvqqdg/tK6Bw7yXc6svd87TrfZD16PwRMTjCPX/
skKaFO3l67v5I7rWzGQHPvIya+cvrLBQS8veGBQAh786733Q4aE4F6r8HEE3/F/PcO/M7YrUTJFG
Hfjc/URmOAryvJb5PRQxeSSIc6BBvWYy3HNCplSsWspzpgPsFFmhjiJzE5Qf12JeChuDlQGR1WuK
2KDgpHiAtnWpMnbPufBL2hwU/j7Q55ayUQCsPQ4pYgDK7UHnoJbyNzjt8B98LS//rGaqyXYd54S0
5X0Gj2LtrDqp14N9CSwphS+JxuffLopCKhkRG6VZa9bhWjibWk35fXR550TdSLsRW3ie2oSXAwX1
cFP82D0V5NWbI1KsuH4PCl9HyYXnydytS3L3AHpoDHfcYXUI1py/HHu2Im/OfsOAcDGzst53Mv9N
NMG4Muz275NkX0ZSWfK1Lhvm8zW0DAFR0xBQn1YG0X4YCPccYLXudtgrRr9tFlsgSZgZ0AxfKne6
ix58cimhKyBPvaEttp2ivPtabaxshwlGWnMi+7j1y/WfjyL9pWzG4aaOD/scMcUyJ7TBQWpWZqoP
pMwHAmFfYSwEdEgpwd5ISTS7Bpzqpj9nx6s2BHYQGgAYaQzGndBCymKDUE5c6tw4/xkyrSz3oVMJ
BnGi6yeYpt9+RbjdnZRmkgChnzSZL/6xp5OnHTeJjleiXQIQwWxVKQ+79Q9s0Dw9rkB7fiRPV/6f
HHwD3lpkvrhVMmvxvxx1W7/44nbSQ4ZCuNkguRf5w6VOHvzzWUkd6Sczwy3LCeiBv5H1JavpEiBp
yH2BWwyavAdBoshSlcwefLGiZQPlaODl3JZn2XRHcz6T5xfgcPEBwqeyjCMgm3EokoCQi8nTuub2
6SmLIT3V1qnPbkkH5/Dc7xXL6l9wtxulcvsxd+/8pENnYrcd1yK2zHAAzUrGG1dr4mDnssKEXJAV
nMUkepcapHF+RSblgvsAYJk2+CCqm00r/fU9+M5BpEbu5nvB1ywsXuxcxstaXbaiTbrF7NC8yZmh
mEBakvrNtnv+WJKag4K9j5WP3KrNwYK55U/BSucIpz4v7y8Gz7hieCAw0FWv7NE9q0o2X2e1Fqmb
qG8S0YmQlLUd+KsvTYOiPk9jBWxMt2yT6Eo7Q9abmMtZoMdKfcHtI6uMGMm00OCsy6YmLqzR4omZ
RymHLjL6x5+Hp7ZrXdXx4kFdX1Ic49YLqEwJUsl6AmwzLHVDG0/uo4OiZbg3wXn/zRdPx+8svZRk
vAjRfyRrwOY0uomz9ePVoBsrEyK1Hr5pW8BQ8p7HSBBp4kJDxndAa/I53JzlYMrnwNCGmihTPqXa
C2pPnQHy2UrdoCXdjjYHD4AbuEW6JcJun9OSfavKpPUyhqCxmyRXFM38+NzSrAVu0SqTVnmRO/vH
AsepO+nAFvrQUR3mIxRns81dKbupQ0mDm+x7nUq6IaubWhCrGIgSxY4J8ISw045VZsPYFhXMcdJ8
SCxAbatfzy0cyD/mt8tekkQYI1C6SxC8UwzKiodjfie7vLge7zZbbMmfybL1Bi5TTXzLHDxKBIQQ
795R/3B+4XEbm5uh05XskRGNy305I8YxmvaLVb+qoGIv4G8tEbrelyD2+4HKDeGrK9StYIToLb1m
9XBCmuevBlvQIOzaD8le4FYtHtpC2mS4wZxocT1Ii5SOLXzBgdu3YpeQaikL/QH7bfsKoE7uWSF6
wi08SCOGfN9gZEopfNDJiQVNCToqlhBPvDbX5KKRxBnxzIWJGOl5Gsaaibzp5PiDGzlesgP4sbue
l5cWw22Zzyf2Ba0ZDlEsDVbYcMX11dhVp0WaJLn0NafW7zzP1ORy5Y6CZc3Pj5M0j5qCIrOXB7Kc
+XGShQYTgCBXDV2Y429dm2imqq3cEtzGmIzF3xb9FUWIybgZB+pC2boa5HEhT6R6SWtz347nzuol
LAkeZ+lY+L/96FdocJfhhO07B5dKghEXMNlytINmlseuDikNSgdG3oohrO//v8xibhaOPvhekc+N
1VFKGFpwrEf7OlpIJLd7G1JSuoTPZvPEmaU6XLM63UuGAn7nLmP1yhWrHML71gL0w/KD1s4K1BKu
2zEmx2qCIX/ndn/7naJAx1WW4o0sdjnZ13OHiRVlwL17khb9lmywtnRTjtSMaPmoTWF714e3HJDE
97b4zNeE9ilx/vOgGyI8bE2a5pNbXNzyGVxr7zRw63vLBOBvnD4PxaORKxXSMGF98nPrrBkU3jqw
Uqi7wkvnT0DvwXHbhxZVJjRRwF8o6mzM6m37+wzC1J38DI4X448nAEM398XlzlE38fmi678pNTPk
e+pqIpTARxyAujHNimKrShjs+kFx8+CNkE4EcuwKOi1cU1FmCTYJc+Cra46CIhQpO1vJvou/KI1O
Q4Kt3eWGYUnUqgqWwZ5tTa5BOUOX3tnpb0JmrGHpwiVQko0rbGdTfXX0RMxxbboESl3thzaSLNrM
ydXKJdaBtgOXTd3S7Qi8sZOxFs9T7fSiwXr05KHKesRn2vgC16Daqg+zvaJGduLcJZqBj1z5YK6H
bNjKk5o8dKkOnknuswLFel7gsRNTL5ZnaWZWQNB8Vd6iDOCub02OP5JtyZUQwSKWOkyFIC9RcWuk
/dCxE6IekNC+cbcZxzeA+RbQ1+hD/fcZyxs/u8FemkMOnYJm+Uz/+nTp06dlEgetrMge5HRI5Pfj
3seiydTSxGX7882VTErAqV+8aqwM8xTUm0zILdHNovGTcOOzMgc1EKkzQgeIteuZPC+BvcXqUduN
MpprEQphoCcHdQqfZ+piFs932DWIrhxCx+FsGgaU1t0Ql62x4xzIp9MkufU3aC15xXvRtq98LlQg
YLrTappAk6+US2nHOzXoFX7FDr7nFkPH20G56mAQ8aRoKghSe2GhJq+4bUjiv5AdEvYzhDUbPAel
ysaXeq6NPzOjdJiQJzi60/jH4zLtR/hUu/iKeXky0P+3n6wXvwhuEihOTwKMyNrgnhPBgN12JgNs
S2KATWm10wwMI7p6fkAhz41sst5dY+h1hUDUgj/6xi/CszRFg9s4djsBsM7yF8q4JsZOJLeMnEQv
QF7MHQet4d+iFAz1aKPwyKu+crIMhZap0aEJSyJN3DbBEYaKbCCvMftaWh5hdw+ANgRmqsxBvw8D
cY+9+UWkSVLKN5lSHhyMwchn3xPKE+dr1EFwWd+dbJiX1yo63W+SbtO2GKHJpiBowMqzG4uxgO36
qcgQCArPiyQJuavVIjxtV6G0hu7NVQHErvfvWQi2isLEvz8CN/f4icNVTbvK1RQx3ZNdB0H84Wr1
hAU3ItyQtiG1cslVT6jI5N6uZoGtPp8DPWVtcZ1JZx4eMwUxw4n6+8WsOI79DEl+bFW6KQ441Z61
A92G5HNv3GssZCXOBfK5e1wRHJcsvqlv6kDJZ1T/ZiEGXjWo+3nOrGryiWURCKCEpo9g7Tc7H6CV
43x2DtPsgWeNrkm8YVMicHEWI5YFMbxJgu1obU+qwoGN9gYNAjdnaXsVZo3aXA11hOSQ8fQXKaug
rB56AHI+44BcaQv1ggfoEPmuTX1YkKPQX44z2Ccxsg2Dy6J9HfLSPSq9z6VUmHI05U8DhBfnd28/
HNRbxgcYcJ7qCVw3VM+jzm7Ep42HQpdxE55quqFOKtCCQvR++dAWD+m+M81UWVDmiVCNVtLi9vVB
m5fJbqVjbb4GIglCVVz8wR7EQT8XcRBloBAxOBstUsJxs8Rsb26gwm7ISU4uIAVMZnu8pXJcTc+x
cvlgWd91kZcRu6DYn0+EUpDI/tE6Q9a35b6gFpMi0gwdI/1bnDyp/zlWI+i6BQ9CIE3IK7AK3T2t
M7UDThlI7BybjLNjNSQTFM7q9aB6UnnMuNVgalDdIsQXzfaKrjNKfokNHMIziMzWwtwO0oLw3bRL
xS7Lt1yYeGZIFEopD3Rqy5dM/0J6U86XLss70VlERAY0lEn0YZdfHBk8qDy9MxgggwSTD+HKvG6D
XA/zuU2yrExYza3cwgtMPCu1YIaFvbFazrKrK6Lz7HS5Uaqg0HZbEWFnOFxzOJKS1sQBSMXmaELN
Ez4sbTU6/m6asNnfXSFZz18xaHetgVnGHJe/l+gf25EpkmLF2Qsu6kAv2TU+aoeGVrqwuYCUknjj
nSFRhreZBH8Sk1/dDTHpMZM8LRtnUSJqBB6TdeBjQ/ZI83b3MbMUQWxtNaAerL3twuOLdWXDzEgo
zLzWX3BBT6U9bNfwG1pi08A3FUGM/w75wxUuFxxc9nyPRd2PtMDhbcCSkPGSvp0TDiCKqLt+vIqg
0oUje2ERkmsOa5mbk90TDDFHydeyDLaALr8sU5LnvqCjUy8FL+N+UeRKyh+1LF5M3PknFiZFba1+
ETpnw6kEfyEUH9xaDjC/FC0cRWq7Bm6FD4c0tztd71azZ6wmCTCqYVoS88AtryeDp/Tyvv/yAxQQ
7sZXqhYeAtUNfqArXCIP58zaMYl9AAeRYUCHD9rNaxkU61IwdNC1SLrN8AlsTXVEFpkJFxNdAYuk
waA9fJEKSTjBmQgD4elyzcSZq5a0LxErRGSruwxcBnWI9lkyvUVGz1Nx1SGzoa023TKsy/yLQ1W9
9Fi6wHDCtIRP+wA+mpSrLTKmHetjjNuyxgn1MT+5hBvxt3YCRlFlDpoNy/f3xC54rxwP7MhEz5e3
2IT04L67iV8mewkqwxDmIgcjuapn84JL/TJwXUI+/GYL5+yNkufBlFejjzhXbrryP+QR07ULtsh0
msiANxZAc5sXQ43WsV+Cru48O8iR41iLqPILgDnL0idQl6OLVBgd4i723bLeYdp/xyOpYbKoaofK
4jYBzHgO2R7EUBywyZuBXrWDqnGMaZLGN29c7q+q+o0xBBrVYAKmkJg88Xyr1Nf1Xvzo6Mr98rk7
L7Pu3WQZZcw5C26C7nGaOQqv28Do7UBfccDLM1ZNqv1i66KX32qx58ky5STkr2ANVkjpcoPth6M0
SjKIFXPApIpijgFMVlUiPrWyUZq6p2HtsnwMUI6aoSaBTRA1pAhxMaP8SCgXgSzptHculU7QFFPu
k3Plqp9zI3DgCqVJMpwxehH7lovdDndFydeHCDebQlOJWPsr+iVPkBNbOroyyBq5YiBueEN3Ts3D
qZfhFyRmB+sdWKe2zkPIDKHmRS1ukfuaEbVOWCsZzmn4fy14DToUbOhJf5AeA7sQDDet58KyT2Ws
NHMrPbjHK9kpJZxSuG5yoo+Q3EZG+BFDDojHT082/N2Wd+1/dGVPYUAKCdCoEVDzi5BvwB2PWoIA
PiSlEul7F/p87qhqZkFYbu9qfrLJXfSfPEJGZCIAkZHdZBWMQRbiFiN/pd1ubyKzEHYQxSFx52BS
PKffZBH3Mv40T1agyy7cTRkwza2g8cElyYcqi35uRXzqLSaAf89DajmwQ53tMH8ejDQ4C9uD96Ph
aQmCzYV7lHP4d5O4gqyEMQNJfWok9JsN1Lq7tBvxLwXpuLpDCkgbOnNqD75VDVoIJ8QiMzzwmBbq
gzFH4E4jnKAol3eyi7DHcc21Xt45qdd48uBjF8yrRLN3yMlCmlAVE14kLn6OL8NBTPPPTPBpZZWk
KOVuwQeiJvy40eHN+j3L03h6OZIA6gfSp+HIDr4ptoxGykrpSEWkzW/bNK6zVhZwZ/oK+84OtoLk
CnkS/OE6l8epKkET3qmJ4uCya2I66X//bkj9/Z08KLAX8b3n1av4YIwRgyCdx4wm+VvRhpU7JuIP
wY9KF1o+3BF1IEIBCBlE64Z5oqGjy1fpqDeGOVqhezHIsr2m6PAT9zTUDT1yrmXc42N6z+oPG50H
yzPCkiBm2Jms2jKN6aDYRXZTjXHGwTOYlFAbd+Bk68/T0GZjAfx2BeWHmcHdiXXDoL9ntLxUudMD
Tyc0y+CCrSXjMQNisp6I568CzZz+o1UTULMfnsscLcqAYj/OKEixUMTbn//ncyPc0PNm6Z78vGRy
VWdgYhU43JAgRv5Detj1PLECxHBQIgugE0qMhw2JbogxNV8V7reHuRYTHWz3ltN805cDbRGi4WrK
CT5IDy0/Q/ZXMBU/fJqnr59Yg6i20Lj/PIi8YIlGj8YqpyapJAVVry+WPRA8TzZHBG7WRH47yfgS
B9MIyqHdZ24NmEtyNq8pvPm7A5z8Qo9ij8KiYY3pXTZaIN4obTJd/Cmyvuvi494qXueKBKKGYp4D
zDtXNro7wDk70XX/OwbiN2SOQDXdk2/1NFz+RIHNrsKvwYhSZ7RIxdA1M929XBONVn1kFrC/hVor
VcUFdDQa73GEtsdqeZaDanIUFl2d16ZrDKJTn+c5LPNIH1zr0fhbwPe4GGaRdnb+NNQTEJpqshJb
0eTfEj5VUiHWeziXH1jh2OkDaZLvVtppYzS6eKDMJspiOU2lBPqwqmFXkUTSR7Xf8bDwowaz1bRi
bJ6r2paP6y0z5KEdethluDkn6E4F4b0KBW0RtKp0yaHSF+2I3zosntFkaPu3ZaYuKRx6Xj6ylZ6g
wBoHkYXz75jqZagk7+FZK/sBzEfRsbKMz866O3VrWGXwitHaWRasLXkDsadAgoX7s5eZBRR7Bd2X
acwzB054Bn84fkbYXOWOZ650btHzHjXYJzowXGRFBqCUn05pTGTHGrK1vGwm7TRRZUmn2JG6WLWN
KbIuCVwk3h03s8T0XBf/94KHdWnv49nLFRqITngimeDBU+0cU8HsBk2dhpcwO0E7mDAKm5cJxfM4
4rqQKxMdHQwdxxoJtIVAe9O168XEWGIzmy7+U7JIcEgeUmPj1jAg8tB1JH8/z/KCyjP6+P7hXAEl
9EwYZ7zj78gK45cpgFoo9s2QeXoM/e88FlShcsmbgmAUBfhOJv1tvgZJeFCSG7xTg0CCx+mfyE29
UB7d6xWZbzPg2/2HhkhLY7sQJnBmZEmCqevNdIzEWO0hTcZe1b2I4CKcwwZt35HzEgjuktrGMcJA
2OdbhmnikWMjEm7dSkhmEF27zX0FdIdkHPPw/8P5MVCnRWbvqkximlRbtvXVvMqNitTR5Z5FcvvP
lEZJcoe3MU4oygd51hNIpKOnxcnui4TS63kXLiPrLX4QPtuiOWq1p6Xh6uz/etAorIEJ+5EFlGJM
XdBQ+tHwcJzpsK5ds0Hr8v5i6/3e218Qzb0YV59cUWKDsJVJPggy+nswzz5nUUyyzM/2GRyYtIpY
mCAmH//ppI+K7RC1yM2aWK5C1wD4M7T0h62ux8OzvZagbX3xpjti7Zt0UCN0dbOOBXXbVm5hjaiO
NAzEHwj7bJKCGoKT2sDt70n/uGaseCUoOXu9udyu5urdPuvKhmmVEv3IIQf5cr0Yj2j4+/RLkFeo
xJyGSc98oRUnHr5cD3v/Ya8yGKnPGBhBgFGa7FBUM4CG7iLBya8lEhMWe2VNu+otnD7KhtTrYELh
JTwyqHpY95Kg9pxADAt5jpskE5kXxO+gYszFv+F9WAh7obSzwQOts5Td5xUG9Y0SpVp+0+VCBIOv
ZFOHNMViP4xhLj8J6bJsqXKPiwbB5PZk0ujW2eZ5uFRywORUE0GcSsgO6jRopkOL0cXNcpNF2khQ
ktbGJvZcEMR5zlLARLdlrRlv3pqwfObTJIGI+0D480icPSV17WlTCrg5Iw56Ka+3LasjvE3xtuv6
iYlxN5fgxHsYRyIu1ZJPF+WgsQdYeaDzsPf6sDovgumtlaVxwczT0hqpWZpzni1C4HJG47r2ajGx
/6g4VYFWx/FmUg1Hli0TCQL4/MZJfJ1DxN2S+NWcdM1elSVOeBmgVRz0JJlCFfJeQ6wt91YDn144
+vmH2T8kECtAXDCql9TjGF+NCPaqE+5iQbAXteqLU7qPell1JieRt4Twrzy3YHVHiDDqmGaV26t0
+MI5qnqQ+Z5AuCsqZU8dTozL/MfSdB1OfiXh9Sxts0UoH2g97qTpWP+OY86JxgB4OM30SGlQArhv
3UyKutajJHhQEAhFjK4eQKCNPMzzkZ5J+kUsA9mdlOTyEWKkRC9utehuVcFg52XXo7dB+/33wOA4
jiBJj+K/g23qJ07iVQYTOyx+uMBJOhAJdqdned+0RF8+ohiE4hByHHJg6E5othagbdUzUHgUzbxN
+ztKVuu3mHvfne85Waj9x+DtsHkfhM0B+gcX0GWmV07oHR9AxKhntDqTrxtfMh9MQMEbgM6qK+C1
VqykqgswlDKoscPCZ86BKQU5o6cmSuFNE08LiVxCUCp/Po0swkbmrl//qP+GXtM0zGPOp2IJ5w++
06LMFG7KDdZ5henBRHifmnaU3qtIw1zSTU43x3aqSm9zQKSQadp9wXyjHtYxKyDv9clRifiToRQz
CQSXIHtoFYVLWj7Jpp+PvKs3T0zOGAgpsBCBmXDiSNglivSZfSVCTs/w3c3cVVUQYchro7mxyfdh
97c0F23Lbnd29hL1Zdr6zRGYl3TpeMArYvSUZnC9/aks2GNrErZUfKjCojbVxKhSSYfA+pC4NguY
eTMHWtCQL5aIaZbF2B6dPfwRuxJvyHMRRjzAqm5+479uxggpCBStSe7GICRFzVulAhAni0S/iEsG
LHqCVtjRsJbjNxr9yhoiYv7ObK7Bfa2PwnP1cH+OnGbGYx3eNOonTiJafG2UUkNC0oaynwCCNtql
J1bj/DGldDjtQQ+JgqC/RfudfvGKnVrr+up2UYly6GnF3M9idxMVG0mSRK8RjHrChO9fLEQTWVJL
iKmtKpBQvd5QSADPgbiAuPxv7JB2Km6zjNtae4GLTWDn9PoFjAVNPz4h1lxU3oitS80mHcwZfPoO
+LlZfZFwID5ALHpF7LKxKZF74ptPQOrumcdqnXq7bGZJvhKeWYT4VB7oB3l5lO2UTf3kevZZ3fEm
mHmCkF/VRZUvNIyP36m/AO5qY1MXNJmKOxm7APoiy126kOLVVavpTbeHQdj7gOcW5aQZzdYdLpG5
UI2bagFEBpWTg5zIwTDxjS885P1LUw5UpKdu1HpJMVLxwY935V5wTD+pk4vo4gCXzvZBKamYcMM4
E8RbR8wI+Ykiwt5+rYFaE0X8Ndw7+/Dei32PdHdDsxVY2JbvO+BmSc0al5MBk+WhlKM00j/I/Gig
2ZCeg/rcOYhBYVD6nKfMRt9r/iLMTmD7BanwJ/26dp4Uik5LnH9Opc8qrCTmPrebSJ4/u0EnUQtp
UIOLhMZMm2fBbMbyIdPyCF513mBB1fdRxIx0+AfiyZtb8lLmtT0saJ+uLUQA5UsrXApLnPacTHgv
ncLNIhi6veENPr2DG0CkNq1Uc4Xxa2bFLrHst+RYDE0MUFG0eZP9Sj/soNAxGKHaynSDXGDn0TN/
wbTu1/1U8/A44vdS7lGYAEeMaztTtsUBkdV4A3Z9tYIwbAH1fNmBG08hw3JOZscjl9Wz+85fh7G4
GTF4xouN5/bcGq18Q0vd55CudAeHjTpAkRU7PXefFFV833J2oka0zO8OrlgchMVtnIqT/Wo+0/LL
7noPm+kYDSWttk607PH+0asRIbPL4onjfgFLslQDnUrzAHruerQrplGX9OLJpiraxZsW8gidZE5I
BgFFLM1HoZ4MgTetN4RuXf3RrX3/XlsCEOxKNxisPaE/gRkiSfXetN77Kzzh8jNQJSsFqa7WRg2Y
66nKKDlkUGHPwt5/DBAooQT25eLtSZIiGgg8Hrm/XUdCH7OC3e1UJmiXNuN3s7EwBMfLGNXIPSF0
j8PqzeOCNkyQ6bxiy/icTIyEBej6VV86b1EfyIzhvYZucerAuLh20Zvzc1YTbRC4ULt/KsJ5o4uu
BzRbafvqNAHZuhtd/Hk9ApmkEB/HtYgiZfOTHwVGY+WBfsraLoH5Pgr8nbRnwiPmJJlG05qYuZ7O
wizduxbQkRyeW+uwgWYzLE22QmV3NTWxmE4AjxychrkGxrlByQdbNVJi5yziG+bc+bJ6AvLNJl64
whnvGclltjNIFVxmL42LkA5P6Qz+TMdPjHLm4f/64D6RDpT6divCxcworbTrAScdTH1+LwSI+ntL
TBv+5wXQtE1VJb6RSK9633WvBy4CoN2Fw6ZYfU9+2kjA6eB8iw19yLpyaTI7l4G6YPW27jb8V3Ui
JDiUl6ZLHJxjzZ4W6T1aCcaXtLVe2PHF4h+aQOrBfxSI8InDeK277t00BgwQGcxjOcCecuO9GMtv
kFOFCiD2N/TaIvgu5KTPWwwXt+f4sRbNv13ANFnKH2WMtwuif8IoOQF/LpXYAWKc2h5nhjeiOGkL
FmKtS1vnvHwBbw/6sV5OlT8lUqthjSlFVt3rhxELD2H51JVP+GYDF3GBE3HFuJfSF3tqq2w5B1sE
bHsqsobWS28JH0CBZo7qFkY2IrR/WZN+m8Vj1IHgJYuKHcOkKKPWzuexdQrxClQF9owJkjbJa4x2
VLLIvpRfW+IyriLzEnVLxUSP0MjbG7RkbQjFNhEVZ2yJOOIbpTxu6sfIKUrFcbCydZwcFvy2kExX
aCiQM1dJAtcBopAehXLk5bXXFKEf4XVC4b3+KTdjCOpCf8/ADVNYGPq8gHsgUpliVc5g6rC0LDl3
dUHRAQRD31fedTLCxuvM7Uj/fB/KZCiDhVg91a/EqVKU8el/g8T9uB9ggKDB9chzJ1yDAagnS2z/
uNsv+sOhlVZ/qaiAr6fJahWXdjVST1fKFP1aud56pm2YjTcG/b7OqYGSOYb2teh77aNUu68h/yIB
bN3jYieGQYUL7OmV/514k86Ld1cR5GjLld+x1Zzg8dz5JPp5gKA5EPSEoX6JWW+b54KSRNK62fEW
vANBmbQ06USMI4HSVda+Tyy5pVG1Yz1zid173uZ7n22aoh19K7L1oK5348UaRk5hSl7euaCSCD4x
rQUDhRYMfgignwuvsDnXCBuBDQksshnf6JIhK9Lj5ccl+4OyEb6aGjRL/eOS6SgwSxdHyWfxykvG
3NcwjwOmlAB4LyqYHcBNb/2gt8CVz0rIgRf0RyoPpHscf4d262YTsoSM5WBNxCZ8P0Yt2xPzkbgJ
ItrnitIlQDkHgGB6Lj6fX+PGt6SDeUCf7u3fJHDuDbac0BqvbXJZM7/V2CRl9Syyw1O2ah3YXaGM
3IUp4ZHm4yF1Nd9sc6gd4h8EjKt47mdR75PJHMBgC6M2C/qAFrDBy5W2Gqjlj3O/MAblzGrZ30s0
c3WcOxMEhzXvB+GfyloEkY3STCVtZL0mtWGU7xcYDNEBhuFXAFvfwQOY7aAAw/ULh/insjkUTmn6
KpQqYHUhcOgoKweEG7jg4EoNwZ2gTAPdPGJMntPoYgRNx3HUNterjKOZIQasd3mS5CryrgDXjZm2
UwOfh4hxA3d6dZ9HMXOlpvzNQW180Pko15KRQLIvPwp3zjMaM8BKrsHp6HggZrfcfF2HFNVL0JkT
1ftlOoUYZihoSOasE/b9rebrxCby9jlHf5AD193OuGmbZAr2FW94w0xjU+U2GYehdt5/8GnVtcWQ
C6nEFX1VQ9Ye81jrxwEM+0IbP3QwbcpAiCdyeRelawZyV4b/55vyliR+UvGNqHqE0waksqeyRxLG
KTrKh3e7rzNI5g7gNWAVTNBarx9VZXeGj0i+1tFjT3lfQoLEVyKcrXHefXHS/Dy36P/ZQAQiRx37
BCD9LWFDnbXwWhEkM2Ww+tmdAli7XtN0jnok5L3bwXC1XfF+0YKiTNPF0g1w/DnGpD7xRDaW9NZo
gJ4bezdPZqiQGv61IyutPgjC5hRQSEGLPFFvSw9MPyzYMr/Us/exJpBcllbSr0FneTTrMaUJttA6
ozVxLhHTQo4w1cWvwvtY3H2e7Feylok+SwF1iMXWHkDOK80++KB7I3eKApPtW4N0M4t41eFUNcIE
0y5v/FnR8TibNFBrAP6CojHES2OfW+zDcV1+jgYoASIUXv/dkEaFWjAwegbq0ubo/LFtWIw6H+vK
o/bjiPddk3JyqFfBprjGiYb7Ov4qNwyQMNrN7DRrqjVjk1HFfLfAMDFJM9DX18+4PSoJvRdMR16n
2qbDqRkB1I5RJ7kNEuIeLFZwmLqGU3xjzi032pqimoPmgG1wZpeih+BYExtRw95Qx+esR4QNyp43
8YmM7kROX3PUkYaxVetnxMCES3s/PFgxqsPjhalQtnkrv198jgMA63aVzsf9UqIacMRJ0IdKkU8C
s7+iPvoTWhnudUY9nCB+uhq0n9KlGm2COKgVP3jpiGZT4sKKJGDgi9xEKMgrT3nnmHyC224SHPtf
HMhpP+nA/q/xKDxwiUtWQNrpQtFDQ6l9dooFHWmVeDVYsRjRlIrdMPFmTrKyqLiYOzH7WAxBtr9B
6xEjYoUhEZy7MTKAZSFgGKLVVgroFc4Idqp0nJBt4hNtcEpUcaYRJUnNZj28IYpMTns9xN36J02E
ZfaStYfIjYgKwfKCb/6hTdyOf7Qd75Ymt3dU+Qt6b5eMAzuGGM/iKTwK94Li1DdvNi8yPfKmpwcY
P13Qzq4fKSBkYVmSsyXaeZIABhNUQH5bCva4+aAPCxDltCwzdkUytP3eU0Cu87A1dXh3ClkcoZX4
X0B6uA0pR3z3R1ju3xY3+0Q/wUnfT8hhaTRyAGSqlLYBtEVk0bgYY4BX08IkrZ7NyOkdkukiYyrr
3Q9AQT0/+BJ69Pjk348YGJquqagoOVwRNiawRKBFdvGGZ/UIAx9c6COmtvF+XK2xQzHSu84c6rel
9y0e+Q/QvXZr9z++Y84V1iWc4qPVjdyKw8mrjLsr4r1ozNku/kfFjHp0/60zpCS/N2RD5H2PI2+2
TVqmDgHktBade0Q6FeJPwTQvzNFM66pTZGLwad2vw7wKlmk/eVv1vUdXC4L4p8k7gRrMtTEVUgQ9
ol57qxi1g4zRw0asxv3lz9Npuji6tEfTUBCstlpZJM3ASDW5mQatfvXqU4z4TegP/8GHoFhSTGY5
KfbDztRe6zirRUQZ+TeijMlEyU8Oxo+j+8qMwNBV4UuXcjrTbE8W0uollFN23JVwTxL7nuK5cJ/w
8cmqtVoywHIyPtytBqd6Wda7x249qj0yBc1o9pyu7ppQqRyBD8N/SWMDUBBpsudcMuMyUu/XKBpw
zAGcNCoUhr6cKyM14k624+iEAHb1+Iqxpt9HlECxmzlIO7zpnt5SGMO8EdnmbKZuk0ww85vmRRIT
YdGNhrli71ocj2brjM1UNwGd39URBcceGU9HfAd3tWDWi17dv92OqkzQCE3aYMC4vzKle2nkOBIU
4JdHkDxdu6C8e573lXka35lG43nSHOxUxI39RnuwlbpSVjoJ3q7E5urSeZFVF2kwkP4SSytZX6Kp
JLzameZO84BDt4CK0ZdnAjy+wMNfF7IhIIj0btJTmu0ZHqzds7xOvtIS7zgkwoqpat5FElpISM/0
FqZifdMsuMCao1q0Inl8rNBTDY9gEiMJU7bH1R8HXu0cmH8bEwdCA9BtE0o8ysJOsDQ1ZvCir5WI
hOnvMvO3VBi3OL7zE/xHJa0CyuTFvc4OjU8ezx6BJsVtdGILSJdV/PJg8k2m0fnio/UAE7BIG/SD
qLoe8zOoWqMJY3EMK3VElCe6uAjW05ZQq0iLUbevynLwkupTg5Z3IhoYFXQ9ybYYnO+k+LZyvLgJ
KwK26U4uhZSlJyItfhjAOXFVvsDifoXI93thGw7OkcuKa9HjiygRaQejuhzTQ4g22d6kQowFNzXP
pKJLteHW7oeh7GsEr8ofv8rjt5rPjQVDd/+oq1FKldeTv+KGdKHyeKI99mOoMEGXfCNFV4QQ36jc
qFYg4NJy/uii3aoc3z6An8s1wxPbShiZHV0s3FkymG/IAT2sQ6geq9DTYJUJ6TBSo1OCsDNHbZkg
x2Kmg7gYFITRbe+YEDKAJ1SR0kMwps7tU7MTY4kS+33ucslsmRQv5InL+v1uK9KN8mGEycJk+qYK
9q8qHLq/HuAS1D38U1kwN0Kv7VCg6jvK6Hdb5qwTLbsr8J3QtROZwRwK7Js+EbNMdge/pBFGeSCQ
8tCVly9lRQsgrUgH//cJzY26YtWucm4SicDN+kmUfoKveLn/w8MFJUqITiyG81o7DLcZ51pWXBD5
Ke2eoTXi+iXx+2YTpBap4T8iVQuKEMNUrpoXX+0wvsrZU+n+jrbB7eudDFRTZSFdhaVO/bIz9lzg
8P4dL7RNEzsboOUOLwd/viimR82Bpqs8euR5XLzpqEO56P2veQY/PBCGerfZZhSxmZyuCmGXmXVa
wRxKxvw4P3DEqf+8Cul1/MUGoncIJEN+03VfWppgZ7j1Q2dhrQJqU5uDaVEkyNBMYJVUbwH1XOkL
CF/n6RisXaL2Rs8P/h7+mCs+NAccU6pPj0rr7yo9lhi2TBI3yQPqEZaNJsxQSqamS3+xRcafuU64
AyraE+0qzP6v9SbDle2x0M033lkp+yAeV7wBiuiuXlsTHidAUtTsG5yJJvaxudTlKci3LBAXuyna
3gcKdM6sy1Ce3LANoGPWVDg++aEzSCKKM4g0iNNlB3l41zy9yYRFKko+sRPM5NUM+c+sTf4wS1eC
VrD24l9/Pv34NQpFxYefZ/1IRGBfLkARhhwexynjXqBGlmwjuWCno0t1XYjrqUaa6pZXK5Z+h1Rv
SX5bkL9KPALoeRYdbJ7frkR8XoptoJ8b3Kf96r1xhy771Z0nQSh8PkkSzLu6ywDYujHixkkaNzok
HBG4HbK+sYzWNbgqcRvO3jcojGUHXYKa6iKdzSjEssbGPd6yXdjKDwhc/XXCS1ePoz+NHUnAv1SO
y3w3BLYBkn4mHOJOuBzHnykgJYytOaxqfNtPD7P+PmzFgA1v4R6yJswa9gCWvkCk8PENyt0S6VX+
aA5RGFPa6sCpZ4JG0QUXzo1ktEDuW2JWvsbXryWb7SaMl9jBS7sGxtfb3fB1LvMx/LR4SbGjZkPy
YP8jraFgN4h7aG7c4atgZsM6Yt0Jz+uGcTt0MsrIz7tbkHINI6CZiQjF5fGPOlgok5HM3DX/mkhF
aXO1dQvglUGRKoopOt6EXdyVWsewFspeZ6k6fkC1plbD5y1ixkrHI84AvbnXHkqdnAjRwS349DfW
Vh+cxi+/BGZrKTYUaDAzPTu11YVh7+Icb+vGvjAygk69E1AkpKZ4txdgchxhA0+PLNxFnoqBLyBz
YzbIiMMtiK77v71sIXegJDpfUyjIsxgeDdkfgVXw0JypuNTZMEac23BH8i771MOt6H73pXM4fDBU
nHGRAHVDFNqOWaLvMMcOhVhKaWtT5KfH08o5heJAmd4dtCDrHhrv9A0GJWUpxFomWbuKwKYN98ic
4O5uYY3EzOH7hz+fgv95K9KXzUSbvV6OPqizzFWCdO63uB4yArZ92dNsJvQoGHwlsX5bAnFKPiO2
krRpkqzPwY/31CHiV75d6rTZrF4ygDrl6+eURftbEbxEn5ddKZo1QgLJngjDOuNlUeYKTt9iWiX9
rahuQ13OT7prGagsPdaTuf/lS/7gLUZStj5BNCEaCssJxqlOu72R03kYem3vKSK+bubXnCQ4LTl9
qHPQxjFwJA3C72lCuhzi+TvY7bLdut32+C8NnbzwAejgcadBHD2WOQN/1D9mCzw9U0mLTst0nK0H
6ep9YiJp9SMb/RXrWFSWs+O5aZy5lI2C4d/cD0wnmssM7DTk4QtolNcB6465D5YgdIRg/tUIgu+3
ym4H7Xs1ATkqubFNwVvnbS8aN+0kM4jYEKsn/uOlGYwxmCeSD6FDj6+xjZJkliAP9R9aDrnm09nC
XicaanlBKO7POa5PLoxf+Rww8bz0NxfOkkhjSOK/hnUtgiTK89rLTo5JFCGlno+OV5NV0v2se+i/
Moxk2HtFlqrUikjZ/lmLWKeCtwKmzak/zPNxEv4lB6wyadl4IE/FWetwJHUk1f/MrSUFUD2xokEX
mjGrDnw2MlwCPuz1YKJ3kSsk8zmUWBmKVTmy2J4d91nwBcicp7z4LIuifhftlBXRRgXNR0gdjAZO
0Ua+bOouk750d0VzFVk0mTafnJBR0Apmz/zMWw4vbqWWMI9eJqlUHqRQ0MxEr+cLVs0IbhtpwjPy
99YyTif+jHCHqtl04eaAtJ8MFsF0OryEx9vCaNa2iuSdkQTGuw3/Mdz3h5k6crPAjuNTKfVHoglq
BK75j8HZmWbMAh43NE2rsrBVNk7lDhJOXO32NPrkec/7hk2/FxzDvf7UKaBN4tynOBmRy8PV5qDs
rbZTiPXxqu1jjiXKMsvfgibGGE2ZYzKC6iAX6x6YBj03yN2yqVb1rkyFjiKCtF1Z0rcIuw3WPN4G
T4LR/glLO40PO5EJCj8uGm8jdFGFZ1puAln2RUkCijhh8OoV00KJxwK8ngqGITHxjZ5DHHd6iX0B
4u2nTBqPW8QRRZocRQfqMGpO8LJEIL56clmvGKuHMqgCN5ed8qMAHW4ka6+uHeS3UZu3t4fhZ2pc
09y4fLP26EpvaQlCGAsjx2RavNhCLx7g3ZltFmbv9fzySrWuRWiSd54GvENmYwWIoHFebxVKVxIY
Wz+Xq4P158Yw6ObqZ7Rd+LCQy0WTOwdXNQION/xDi1riovT51DkrHAyIL4XvnE56U2Cycc4DRx8j
ukD/8mnqjgqTKXUSOk36UorLkm8w1c30Cz6QgtZIDmttGd8je3pm0ctFiV5MLmGY59zBzh5UFlrT
hCzWQGwmtvzcXqf4gcTzqTGxqTbQLPmvIiMKHjzOedHIbV66Rq5hD31MInbx2UIeNxXMcLPr1Y4q
ThU+B2436gzepcTPnZe1xo38amIPASUUtCucm3P7jHhRGExL5XyGwSHhF7InVy0CitqmWgDwzDXI
QfT5piIxCmWWil4I6rpdQNs/ChJugTolRMbquUxiycSzTPos1wpCmhoOvbX8OjLp1ssik7kfpoyY
a8YPuwst4NAM74j4Zg+7H+V7KP22fwcYo59FDumDVYmaC2VjujX4Kz84MWYjTzemSq4ypKmqCJIx
S7etWjBeanlkce1alPUN5HhL8vXU5KKbNS4W1VJBPA+m31CrffjI6Y9Z/8cFsVZVHKkjZqdhk2aG
ES58cFMcGl0FPYMg3Xa+GdphnyInxRSyDKccskDPqe4Osj8EbD5SJdEFEiKZxMJv2hGKc9L4670E
CjomvAExupa938NzmqNUTbVwu6akV1gUrJGrRB+JJXJ6K3/k9SLLDSG7StOhlMHne7d9xnzl5Rxd
/H6XGpgjyoMGiROalCir7eo9ircyUn5agkVdnIwQd9itPT+PRbl2Xju0rHd1jK9PRyk4ieBOa0Tf
rgpNmvrwribuLwNx22RhXMmCoNoqgXRKWbyflRiZ/QP+jcFddky0pyTWVD57ZUwTX3aXPcq3Cxjb
XCBElNRtgyTteo0+/MwpKBO2Bi4MreuToqcGtcU0fB4NKiXHweqtQcHuPdFYQ5lfTUeFqX5JYUNJ
I8JENBWA//ttYrH6vg6UJSbFIFHVW3mw9cvtJBzwWsPDaFtxzVUBXRE52uVw7BntXTRDU9WmpHOs
i1RUfDmtLlI4vF1VDKudrBYLz1cqW9SZ3XW+lr5HBquZESWuSmw5q/+yuB8Xh62kXgFClfvsS9/i
0FeUnetzxEGEHJwKels2E/Ox9/XYDdR/t1yzuLp5RbTMx4KeMqH4nQJmfMpfcD76+0aqZmoqJlkg
vSu9NvTuY5Yx36MmrUSfuVuSwa8xnyBAbTY9Prc1g9kKgk1T/maEE77ePpOToliZkCrXGyKUrzHM
al2+PTNjPjvODQlLhnUMEE4d+7Zo+rZ4Ka66lXQRhx03xUssjHnLJ72mExnOmEQAKGn8V/SLGcms
/Mb5O+//udsippV2j/wY+VZsBYU4Elojs/j+rO1Hjy07ijOMj0JBKCsbP8rU6Mc6UjY/3Y2+ELjn
SZ2a044rHYKxDJNEWvw5qWZ4S9cM6vjl7794pQG+BbeDBXFXLNQfl9tnNKv0bhQDHZ9s4+E3Y9Nl
H1Z8QMum6kUaeb6ufZiTC+oC2MruSwHPybXXIa+fGl3njpbozhbA77AeXndZgzpsadzpnN1lJERE
l7I/JjXOf6Ds/8BmeugRouCzCRpKNagC3T4zkpQannq0XdHMoTp9CNwa46JzfOtTP0AJGGogG5m1
mVgQbWT16m5XMD1mE30q3XDGh/xDBD8Q2YwI36kqf7VClViLNsMdJcggeABo761uVQcI9L1Q/kRW
UZjS1a8N9M2LWn26pjvs3zSFD3xTzwctrfZRy22amWStJqD+51t7EJWeDOvj2e2Cd4YGjSVQ+ucd
ljh+z0C+j9qlhXQ1IXuYK40/Crgn542ifUFJn1UODQ3acDAsW6Fo/L2RPvYs+cVIsPqi2xNth8fm
bRoh5Wlp5KFkz7rCEc3CCY9Ke3+KG8+r6DA04C6Ia91e8/cgCD3TjpNNjZXn1g8wXwZMcEvPaadN
thMFxW2hU5v+UCBnCRRFAOse2afwyS89+6Bp6z+2PIX74Flbh6sLcabYo+Pnd9EIr13dcjoDmsYj
BEiB98jNm5NRWxyAa2v8G6a6J7GQ4HhibMtX8764Ey7Lcz+LJkJMsMXSrnw7wPw2hLLfqKAmaOru
xKwL99N9oNG+qZwmXuznlJ556VugGEJ5CJCM+E/ZmDVC+h/45e0D8EXOvdVo+Di0WknvoucUXw2N
ASjFMyebv/X8KqzyBIDyTBAnIfciS7dsFSSUNPG5ScA0E58Ze0Ie3CNzdV2WaRUvn1cmW58U1Uzc
387EL/8zmvyxqHer/txe+j5aVOzvvv2dRRQDHUAigLTOffwp/Kkr4/OcekgVxVF4z5kufdA9DCnH
MS4hwpNUvqEwBcGW4YYYhevmzheroT+lE+rt9F7L7fUqpTd17BX3bQOFesDDmj3e7MbjihP9CxWe
/1PhDZ/W4/wS3+VhGmbdDv4GSDHdN4+RE7f6fMUN9YpOBdZYtTDrW1tyaAxDaLi60TBnm489S6eP
hZTU5X85CmRpD4Etqz60rvFEjtS/V6ORITbJzO8j4U5YUNvliVqxJYTZQeR3lZlpZffqsNhErm89
muRPJyc2eJAtgxmTBhOC/JxVp2iKVNzqaFvOaD/pzZsb7vIgV0gwX+sFACcUM3FqKLGcfbAGoFYF
5taVcMkVvu0f+JELButv8x5T5nVfvLM3c1x0aH1HKrIHqQNA6TAfHm0qNxwyIakok798PSYfaeAT
fjMRkO9oaHwdRyvxUfmnRrtv6ApT6XITIiAEFhyG6S2iH8cNQ/TWyCtexl5DVfVRFqdxgytKjFzr
rd5EiLVxgp6RbxM+u6yx1fefWe3SfQSIGK0qqvPwlgG9P+FCjgTXNIWdPfQNNbvssl+FdYb4J3F4
OrIXJhIjKOvucOX5m6U4Ubj3O4uGBcPJuscZwEKI8tR0Snc0ieSJim7zWGxNuiS5ghLDSQFWVh/F
KdAB6qu4tjzRJI7wgOS6RJ5nVpmzAK13O4/MQzXtaKEbxxK3OrbIoZt9/EWd9CaGT++hVkUmw/n1
E+p2a+gx1N6n1oDCDRlNx0sVKZidmRWNPaUkyowVA7PqUuSjgZE1wVBiMP/fp2em/Sy9YYn5S8T9
bZGYEOeInn/d7M/CFeGJlH/JZmGiX9HVCV1T+5uoKRT7zLKixkrDBiMdVwlZmIgR+CEk2jLUqHTV
IfDTnzSmzh3W676ptN6x+RJoIJtEA7wzaP/pR1xnm/iB2dUXSPVbIAYi5KfH21j8wTFHKmPyjZI/
+QKkah+7m2oUsTLW9ho+quYhsMVKBWgqRARY+dQodpuCqTR1jJg31Kmst6fm4mTwC/8dEaurBWVt
FOVTotSQp56YLOV/z5N9yVEQQdhS/bmNS7LjTyFAPnWGk+CG7PYKZ4gWBeeNQ+Df7Mhh1nMLiKB4
koUPQWeDJWk4q7mEVN4AJkf6Qwb0wznrP+8q+yR3YIBq8hkop9iKjeF1HgDf+O0+dR3Zmaryh/gH
UhFjEPyvihrqvmzv5DVdDb4ABUrFlKdX9F++fsI1kzGQEzzwo/DHdOMzb98eg14DTljQ6W7kv5jF
dNgGuzH8sdAuenBdbncVfh2N/YPqpo1NBVBhICM0wznF/VOgEb8nqkTKiMVrXre4F5mWEOqe8ofz
R34m2wtdBqb2LkQK1UyMV/1NskHB4LjJlEK6KvBn4JzkH/QQZxMX7jV5TpX8A5Jq7b3NTgBduod4
F3/05i/LjmffBybyZNrTGSDChc8FwSo16PurCP40qGgEmzXKNZsGp6BzgE7tLXEhSfLWd1NnSWTD
+nO89oQmmAqRPmKE+Cu2J7OtZ411VbU2C5GaJnrYbyxDTG6/TTWvs6kk3bDoXjrWXuZk0MJISstu
/uSem9U6Hz5IfEGMiMdP8C4wpNymY/i2x+EGcSDVXAybRV89Zy7Vmaf6/Kxlbws8Rm80eu+c+f6T
SwPYfMnyV7R1+zExbatQ4KESnfe1ba1RtUVRZo2v3rjljdQCNHrVJ0ca1LW2yqLemBJVwDhk7jU/
F7+Q8c7jnjzbJ6IB63S/JoDHAzRImg7G2b4426NKSuGjpVC/zJfDznRXRpc99LyuPiUD+KtUKoOC
aEs8CmgSbmDB7cJ6yWA5b/vwpS/0ZbameSAP8wtPi/0A+BAY7YAPU+gLQWIY/WG/wkLl1w6zmDGx
MqLHgD8lwLLZmYR9hH51XfI44P3oh+7uMedpk2uMsXV70C3eAfxdz9jrSyOqyDvijOopLLFWmNiY
vgjmaRuM9RFFkaZDpAwpOSkvHI5Lh6yeDlBP3wF0lV3J3UEc6Y+8/T96uSUE5ff02PM7/ZMOEu5i
p5pnlaK0dvbvhAp3TRVDU8JAYGRy3BE91ELAyNwe4ryhGMqRaKaRkKOwfT1tYsGJ1ErNNf8uUnEO
7LiT2VDtsZq3FPnWOMqjbQ+303KbLL1AWHur3g+01CxGDZtd31056rO8atAUVBO1WW0GCjoI5VVB
fO1dPWUJLtsbW9/+Y4vYnJAIPfcnxS1a0yRn5YHTw1GfxTt056YeCu+hbNQkvV/HyFLKvXkvv0kD
/SEHIg6XJtq5uw8IP2iVxGZTI2m7LWaR/CnUNx/5p5uVFvyKs05AUitHTw7ozg4IxJbCHKCT7Z+0
aY72cO8z1zTZ9qh6dOz5kkScJn6qlxqEwQ38fpIjecZd180VAPQsuhIF34LTSDQ7gJcnbPqFAYEp
2n+G7kK75EnwyeOUS0fp8ll6Yxb+LxAIpRQqmKxUT+uYiGvYZ6MBq6NGpE1/eFLZupn9mzkdXdgi
vgrJQ//XJQbwlJK9uiXbRvm2dJYpOsRW3kOXbRVgIH1ZrlMQHnSs55gbNZb+/zdopGD2nW5Ihq7f
Vk9Kjswe4hqKQ018UrhP3rtBl711BpFMNVCts3gz5lb00GIHYhYp1RtIQ+lyJPkTxZAkiEmyx+gJ
OGfeLZjLEdJYxdOTh1M3wvRm9OwcxETg/LmakfXj4d8rnNCLTV5yI/1LSL9Q4u8nge0HI2UVfZ6w
jMyZr6Wvn0TWdlYgoA9PcUcD+PKJLhRua+MhDny62pAVGQM1H06JtTrQJ49wqNeJrt5dLFvbOOq7
wb5YbQgQtdxTCKYm0zsITNc2SvWbNeleRhfrhfE8mePb98+vjRAt1FqD3H/7ew9MvQdu0E11H5Zx
CjQbSHtCGQLnbT0+uhkKsjFexvaaiMwXYbb21qsPAPbXYG2RuyRmwfvGJze9gXwFxvk9kbP5Sk4F
rGvEb4Qz9ASuwxFfbKBrQSuyarXyDGzjGtD+ikXrROhjsJIKJXalnWGe1Kexlvmff2YKAg5vdeT+
XCW1BAFcVikJNQZvQY/wW7PqIUtIU8O9CSC135vvtDm1oyiSlbFNUnJtXhBpHzNhHL5REFGs1IbO
Ef+47Fj6ahOX4R5si3JtXQjJ0+eDpKyUmmAkRF+865ynorULwInnS38na2vNLKt6qItH0aI84ghz
T+usMSZi5x7E4QtplDG4AlByBnr4r8NoSQU8fq+jRNmVCOtZUd7pSR5etDCqGJ8qXgV4t44v0l0+
n+SnZk77amxDAADI0Yaj0XlueNMWOG35Gl4fUHb4NEuD8BVMkbxsa/xls6Uo1e5RhwbOAHlXDk20
ibLkXWIENGREN8dDucIw8mS5P19YljhBE2fX7O0EIYP8c9ahbsbwvSTMu70pY3t6+TqGPyOf62bM
eUqo2HtDMSY8ceT0n5NLKIfJAZrOhKNlzghrlkiQcIRfHuHVmktXV0Cs7r4Dcwd5r96r+NC0uGoc
/Ht90OHScQ0pV9YwOvKjsQstFt9JJF3fWIEj5l/BOADYLGea2idPuRTqwHC0yXmPxN1Fp/ga87BT
QoWdlO9zoqwM+hiXPZ++KVHLqOc0/maSLbWbIxELkknSV+H1ny0eq2DlZAzbI2xyurl0n7cMa8Fq
y+YHFwDwyakS7oIF4UWSAg+8u2/7Xxl9kWVKO5VIkWX422NJsPv35r2vYP9ckz9gWSPHO5NFqE0M
ExVcHsJJZtfQ8fqqwYWZJ3nq8l0fUKJNesiz5YL/SMNhvIs47sbXLUXAx8V1sI30eHQp2EuEPhUt
gf8fKubxDD4cuWwQ3hXAH7Bz4IB7MnDn1fI7GOlBsIVLeSDv05JbIsq5SNDHjj/1F7RbMHNljiCu
ZGY0LhOBlyb0FVA8xUfaNXLZF0/Zu+4zZI2VRYbP3Nf13TI1f+jaSDypsNdtR+mIfEdjWYnQE6RG
dQuYO6GUEs9V1ydRiII3kypw876WtK1ybJWrf56fot5T0DSY/Jh3TcQ3VgMKzaknbgZYzOf2sqKY
5YG5X6GE0djBoDfBCfqj/gctg3ET5sIuEQHEbLOQyFX4GlkFAZI7Wtq2KRaLVU0FJgLX2n0Dg9Mx
lzBiddO0T5ytDE0kJ058zSfmThDZUXWJFcU44C6QZ//j+LdCLIqklG4JnvKFmA1mjhHJjkbqyIv+
MsKR30W4pRIiMh0mTCFQqS5FhqAbfDjPn/hquq2bS7XHff/f6z0ezOHsZS/60XQ6U8JVXFdDtYhj
1UL4PaV4Wz+6U2AiDgVjXsz4qZokhcS/wTKIRKrdBeuU7kKI2op7fbftrjau7aSdxKts3pmBDx/n
7YsQxQpUiOaTpcHjjxg3QR6LJ/3pzomKiTFVuDzeaDuGb9lHvRaMud3jgEdmvHDnO7lGGbIPJ/d+
TQpwRVqZAPQzhJBbwh+77NCU8LjeY+Oq+Gn9A9DojIQ1jejro2ayzmcVXoh8DyrHPI4M8YZzedcf
NtKZLt7HyfmOE0A2l744N81t2PVV8VeDXset0oDqRsFeSY0YilZN86tWwdH54cVvQu5P68TxSnlN
TcZeFBDl7Coq3ahz89xvSX5pTuPLQnnM+0MXJEe6Qe8qsMDwgx81HSg1/UM94MJu/xWiYFEAz6yt
wqj1CCgsSvlYHzPGOE595K3hJxFe6fR0BWv0p88PxcD+ZoANlHCYw1QRdFbhfxCZOsUEKmyMb9n1
OxjSCUSU9JrrQ6Amir4jZl+sqq8MMVF7uDL3YzSFUWLCYkncRTHQ8G6wFoISe3OQXkZ2tDqPVojJ
yczGH8YlCLiMzrRpiDpn6+GIXa3V/L3zb2XOp95C+wSn2dYPI+cCJ1O1+Bryhib0m8IwSQmYaDg1
E3KGe5rw5wHzraKvKgSobGfSP7dk4OD6aN7ou6X2qzDvrXvJ5+FbRhom+eioB+DbQyLVY0/7dC0f
3C5CkuGQWDuLWMX3JvVM9Irb2f4VS+nyqkzC3SngSjgu1OZwXTvpukYOoc5IHnw1VHjltB1pHBWK
1kqJcGAhuu1FDiqKEpBIYyDF6pWHBXRhV47/9yw4qnpILwtWv/aBHRQ0eRm6Pz9lXZcoTu7YVjVS
0394MM0HOKUZjjgs0hdC51CCgnJkcBaLtSlUIV9nHq3Dkd9cVhFzQoTdbDxyB9gEDW+Z24mbDNSM
MppjblUmEbp4j9li7BywlADZrxpvQB++Ksm+wPI1K0kjJEBlHBML6X1UkpcRAAv44u410jYKA1fH
6LRmP7AahDOsZ0KQdfnfLkjjLtTX0AAs7Vu7O9foRoBXEIQFxneHBygvQs0q72AhtjEPSx4LBowC
D5XZ/H2tfvV5/uz/ov8hoBk28HiQdyMgZsZT6xf5juYyXPUNba95DD6mtzd+ZXHG3LF2SQNmGJjl
JllYSOu9caaorLThl4625tO2kmSXSOiCu9s7UlMdeLmDCjkhqM4Y/CKkCmTuJKil+EkMIwUXE4sl
vfOP3WDEVaHKqmRcnNWvGwOt7wL1z/jfFdNiFx98OPTED91DtM0noWPhZVMEDhJBN76i9VAnlDCa
1wHog44BeK6CHu5+cOJEdBqv5/Q88FtC0EpEmOHn7hwrdbu8T7XGs2Gv1Q1kH1zub91wSt+hI2aI
K+7p61SKmzFWYMfyAAADBvPZq9r+iRQzw6RJWK4u3iWNPaiJBySO9TplAz0fmB8QBdQIiDc8eZK6
kk6VI7dsqHhfQmc2dQEAJpgSJDRGvxKabzXcVbUec8bOBKUIroup/Qr9yIJxyRY/AmxMBNH+mmzS
Uutq4aoDxhb62ooNKpwY6oFHPHijYo24O7t2vqE3LEfCare2aSBgcghkuh0Ss1vKF8gKbYb2C48X
L7XnaHv3w1BtpcLztw4E/UhvbXo0pM1GR4Xgk0fXOq9IuZe14vRg4JEGRDxMy0K9W64CqL2BKD8U
Dy34IWuczcJ5MSC80CM/+bn+lpVFdNHybYGjSOarD8sh6oywI2bslPQAXcIbmoS8bg2nAp14PDGX
bz81Gg7kVPy+RezUmKmufhWegTcitvxQ3x/qjnFM1g4STuZ0QO+JPSjBM/3E/XK3GRqZGAaGRGel
lnbk2RtQcJaBW3QZU76fAM3p8uRWcIps8daX2q1NoDJWoXT9/0G9jSiEiTY/75nNpKNgQ5UtALPC
2nTCZibeXwasPUzpDsxGwULUN54l2oMkB1fx1rCA7g6oqndPtvvkOp7+MNWourtq/s47eQUVjVjL
rzIXzUc+rcYMnaZvpKlvA26DfxpLal9O5PcLCdYWfHm5jI2PhyKlnM6QaBvxmKMLMfaog3yJ+ztF
8euD2R7k8SoXOFyCh5PaA/Y9H/M86UCYAiG7JSV8Fx1Y5IntKybCvHW9ecVh8A6haLpvVD0WVqx4
DO1Yov1HNUFeg9FB2E+3F4V7Zv7OfdtYBxheCXjrCTXDBHEPyUSOJGp+INfq7dBJT0lzK2mbWh2l
Tde4OlCouLKr9lqUAHRS2mFCtxsb3GqwIwiv/4sWOjhjWrVjOtrwwowxg4dflzWO/7G6bnFvOrWd
PC8NpkpmpNIsn0yhSII6hpFUcw2ozheGmbocMolGRSnU+lSybl1oVp40zP8TZJRw2oCPV9+9m0S2
Kd3xVxPZFNAM8BqaEVTsg/hXqOC2kiL/hQ9P1zqtTooZnFCqBFCpVwGMseUhXMH4y3/5rUfsE6XD
NNmiN0BamZh9M+gR3S7zWO442zrLFLzwrCrXdyulDxZCt4mRMeh3qLDpH/cpa8eC0WEKgdXP3fdP
rxDhDxm6KiunpBOul5aAZHGXxD1LdAFObi7I2ND4j1MACRsMA0WoofwxAwLb1CkyotooVhs1iW/r
h2tWysY1ZsQzHZ6VWiy8Przd7xtSdJLbfpFa1smrkGPBEJ9NVDCM6s1hWuboXkyO0tiRmGRl1qPv
yeoIX2L27bgrElQIhoKkznd1IVt2ho2unVi9fdQnfrrJTnL/b/6Cw5J6og2EZTA5M2/mdd+rZyHs
Hnol3+K6Umm0YlFFyw9DRe1n5ihvPC7JmBuNIHM5mwbJu1pet3g37tv8JA1GDsF3PskBrbMKi3xn
bRh4JUVqitcr5gbkeGTOp2YJwssTtd3UKLLUkIVLF5j/cHNh400neP9xKYG/ve83zgxjGHeRsXuU
nIxIHkqBDooMYbKYGibBVxICV7bKBI2RQ1o8skKO/7x/6ETCSBXFFKjq78jPbsX/YcSFKb4UfPks
nUUMIvJdHEfLHfkuuFSwN/CEuDwJl0rL9/e1EK8/UXRXzH2qInlNeKMkPK9JSbICpLcIgLxDtqYi
WwueSRmLAPjQwSya8pW76lA0OrEZ5H8I5dk6P7GvsfopEjW2UTMKTHvJzHpd2pe1WMQYLrGThegI
7UhEowSlOiSfL0+oPOXx9iX3tB/x9qlYEEllURGHwWU9C6ESqtLtL+mXSgRYdHF4M8Zv3JFVoah2
ELknY7F/EOol73rzB6Qu8snrVmHc0ugdLPy24FFRIOat31hTxHWO4DY2Vc8JycxPc7YY+43k13Xu
r1+ofOdw6BLIFQ9XOUjuvGU+2ywbK1FhoQ0cCllt4mGz40uNS6It50k80/3tNmUw8H5LpzKFgQ18
FmM5uZwmaKtrZednaIbK5ld7NQfpIEUWS9D4r/ZNXDGhCfdNuVoyMlX9uo5jPnSnkSj1cZ8fBKHL
4YoGfS+z9ABVzluiTApv1caxasUwhP9I+HTKzl6eBF2nJOM2g3pqhSpfkdwN6vrAaJDjwdBje397
dEc3yVP9i23iM+vZP8jOLlMGvC7SSUbDvOkxLw07nHnl5rwuZoCGwUY03kCDymTLGSjZ1p97OkLn
dGR+Rmmg9PGPTkMZeoSo3koy+hjN39cIkiIGoxVNDuU6yZqBoAkZSACgrKwL2UriyZXtyRqBMDsB
Cbcm6C19EvuqCDxZITyK328eflZUgvhZoIrvkQj8wlbEwlGlBaWLtTx+rLmSO1Zeo9n0s2ZA8Unb
jkcGY28hU8XXusXEMvzJwgka5v2vwLTx2FvZEfBJrAihk23usuudb88QCFCTl/Cpz+fEyUEjuTIr
YQLjO2uwqIwuYQTyTj+YQPVoo0G+KR+gO//B60/Wic0JlwtS1GCZSj8novJhU/foxElv5uEICOj/
mD1dYz1ErYg5dApCE9np5JolGC7Us03RRQ5vuSSqzuRm/it4zeh9ktFG/p8dg/bdlnKp1BM9ZsYA
d9yBkCMOdMBH61mJ8zpKvp1Td/YrRNeMNv7BPcBJYCyHBLhAQL1MYgkmXnV5SW146osoIJ+11tp+
DydoZ253kXL3A2ggFDnf+zJgKWEc/sAPOGdezF+/uYdTEXoSlUWRgq0ffo13S4LdRKUkHH4uwULb
8maYNbeJNX8o1QEnXvXEzL9et38T3xYh7mwD2zaCVldeeBPXhYc/2z/eyO12Z3ycdE5zg2EkArDp
syhXgtcHzJ5Gdb7VNbkG56NuzIzdLcurHuqGQZfRIESZvykwIqg21xG9Zsir23QRDmLInSqJ7aHj
/bvT17QnrlCSKsy0bScQfvh1Lf2CDt4ormXMZy8lyQTCcqSxwGKfEJenv05zHGh4vYlCSE8WAe4J
/p7B1dSHgJ4Y4ssQw1gAY7Wq3C17rQmcawX16Avv2O0gwF9XxFe17D9ORAoB2lQemEzUpt3BatqL
oSuOHoJKqGFTtlwy1KtS2lumfD/fAV8b8ghHHELDIrxi2k6YXRWicFjcZpYEUFx9xMRygcRSRR1q
fdG0L0JmdRZsFP57g1jV71a6HRG8SjTvQMn8HGe9A8IyoiHAre1fFrlrG+GLse6AdYR2bvrPQIU0
6IOY10k6WZmOpTYqFpd6ovYDNnQMSr1CjFUvMT9+VGwb2okj2VK5zDSLJJrgumLb664FqN/5UPli
o8fkyBFqO/LhB7PU5jgze8Z418a4TKci5ZFSQCnKSVOJGfWiYricCEHXouv1nOG0Uw2v66ASGWTs
34JoeK9Wrme90roTaNXSms+OOp435Nv3RCRzYBrytQILQPo9VGpYrqdfGscXhfNiC37KySfYguJu
q4GO8iuY4lhXvL0suIS9XvRR/fYfg8bBUWyNdQtcTW3EDdIMwUnKmWsO1WndooN+EsFd32iQVXFJ
cKPzZ3HR8BXoTYlPAYzcy658cm1PZWDNg5eF+pPULYMF8VHe4QGZVb9mB75uxK9PdRmVjoxQQtLR
NIVDV65m9KK3tSM9uiysozGDestAW6i4CrO736KVaZuY7pBCl6i9amZtbpommAII+Cym8FxXDWuT
sYUynIIhF9DwdvCBjDZdorf3o/L8IQg6bzBqXAkmiWQVcFJ1j3jsA+Vx4YRcazFcvC/0J+V5iXmY
K2U0A8EgHUEgJ2recGfRRRo+sUC1cw0oIi0pksrcQQUQDk0Xba72joaY19U1+bKZt3IopYNcOEZm
WSR8r6qOBbcP78+W9nyCRa+l/NCdIgF3G1oAQLhWnh2yD7NJg0WoB6c3sCfnQWtieX2t+ABVcIPq
hrCFK1oXImihkjxLO8IX0lwxqxQBn1CAzQ8aZwOVESnMD5bc2eKX9QaDRynfSqmNUobnuRa6R3+r
RCbwHXx8vLNJKZ/CrjbMEwxFZ2YBuNIJAW9r+1VkPUlo0ibQswrJgb/CmGls0r3Gd82QzGsJldO4
WLfIlwRxrzkXoICpP9DdA81S89pWJRZr1WRuMqUjkSaOtNHMnpgvzH1KvkH+r6rs6LfW1COgQRXw
m6VN4Xp2GMzrCEKFRWSPSH20uBCJQTyYpAtCcUDbBc1JciHbNOZu7lO20QyrTs8aV4PGfYtNuojy
S19pwComnYJxIJgS78WgVW/PSMnj5fppSqb5KKRefcNiqq7DSTOelWnMqxY1qdIJ6mRO/rgY/O+Q
QOeDrcLvnLBtORfjIFpcPQmkPNVwZ8SezBfNpoWYlcshoT9FMJQrR9wbuwsxCTOQ8v1Nvdz9NWk2
k6b6OmvR9uly9c/BRhPbdekhkIQx6m1W2QWcF5B1Dmv/6+O6gNFydmB43EeBR7F5y+k0bGmGlmwl
HpScwvVUTu8ALj9mYQftZ5wRunKLDEX4PoV8oLiCtdQZEB790oirKBP/mwBFptYNPRuy2PwkFQbJ
9hwn6i6lRoLbhMnlJyKQ7GxDDn9ze6wFZVXmSrsa8jk/skTdTFtQdZl3hggd6n1b1bObuoOtu3Fa
1gSOinmAUJ/6fAxVAEnnQ+9NLw1DIuFBjAk2loTIZlhoxTmjju100HD86zUCYEbYrcLnvCuuM2ZE
xgMxzb1otb8fbWgKEDLCKUOudO6ZSl7wCLkYs5lI0AuJ7k22FFecbmEpqSV4Ts5pxy+gYz5q/XqD
33//aTjO33BfLtRWD3/0V7M4Iv1ZuUmlhVJMBC8nnHTwCAu6j6w6od9oC2nmFCrolcKKH91gDwHH
dIt4kbl97HSkyGhDuAd+ddGyBiE9GrP9K+jcejJnP14RxF5NlKKqSaqf9gHsFmCRzIT6cT8v04oY
w9CncVWjSR4SDZf+ces05uz6rxiTDUdcF8ZlJ53ZpMURJS3HWiQpRjYkNzTKMlF6jAoiwGiNJZEd
47cp6I6N4nC6mCS+yq2Ozf2htjHuiNaxHiVi1oIPuOmFpQaR/NQxahHoGCHAhm9M2xJaGgNzSNeP
1wFZYqZd1OsWh81HAUMmz+oV/JGBdpzK+dZTDyiPzYAkMD73p6hnyS2J8e2kto+gD3Co6LjYh5/I
+6wDJWDrSTiMW7189UWcpUpUt5oVMjKJi+3uidFsVLDFGlbvMApllqTAV47KJcdm0+LT69D0Brax
jNzUBTZ7g1bhxLnJOx1FTkAoqQ0wjDj63g+e/KXrF96FX/QJpBWof9+MLUPGOmmvfGTb28TkLRHO
Eo0AltM9hgtrcQEyKWTRRO3sAYnPuGv06OTvRH2ngBS9FT5tBEE3FG3PW2ALfZt8sCuGYYIdRa9A
078VvDgueFZpLz5T7jJzvj9AASpptomBfg/QHhiO8sHXHMRNrE4Cn6/+11mF0QM/KhbWRr0zbBa3
XS8e1PJVix7wVON1YIVkb33t1JFYTwc8q7Ms5CHYfRS5SyeTFkqBi4EHjrQqJBxzX7LKfFfEiNy5
LP+TmqrxrQpeXTjdGDJLZJeEVTMkljFqPOCyqouwDVjvtustGOMJkEbAw9TLCxVc/c+olUVA4MNB
JBJqdAolDiUgupNKDKbHyffM5zRsWZIy7qKTfb/IlvjyffN1CHH6wimYEuaJziNGW841GfYYkws3
tKiE3kg8WGJV5u5SRy3LIMTESBvzj6nnbdgR0NqrQ9qLzlNMTOQCyHcwSN71QEXGIMycKjdhGvFx
Mo3jwsRmWzBGzO7nloB/OicJKKbXd+u75SQNlOrpFVX67Mw4ljpYRCNPROSetzGGUX+b/kl5XDDQ
gHIiniasbHhEFDqaxD2GoSQnZIyQu0gLxxP30wWeQ22zZWs643OIVpglPUYLGoqyIPtFCQSFsGWH
yqtd3azIl/f741CabOOnQgpEyl/Q6Cn1VBkjpEuaZZp61AYRULf6BYXIoawdYpZazLyONX/FvM1B
6aeHL78+edORRbyW+O6ctuYk0HIZFjK6ZtGwvwdlzZHsi270NZPzrW3SqNyuEgDVJHRvnx1zaC3e
xQt3StS3qQzcKkvbt+R1vSvBBvlgOlZTScPlHILYYhwHWINrFyp7h7vjVMu6NTHglitBPmQ1tbal
2rLISAE0THaEo06KdOXhLR0Ovn/WZ9sDRsLj3hHIipP3x31kZK76hF/x/MNfOedt0xZCaJOCXL7Y
pgJnK65Vat/ea5l0dS1i5tLedOpRbU98Qp94TovhIFLXe4pLXm15nrj2BNF33RZmJTJDeoOYQJYU
VEimROtW2LQWHS5IopAiY7nrHR+Tf4yY/+Jr8KcZFNmFESRnCo5P37DBuE7FhaEN3+c/7/RZJOjn
VQlRF05H8D4n6MtQuZp+g7zn2KMmz4dUM4AQY+8S0rcF27dfBnwFjt+ioJO6kl+pWiUVnGm8CFhG
A91x7lAYygx1AD3ldLxBpddWqVX01xbe3WniqifB+A+VbsG0Rb3svXUa+4HnC06sSQdFv/iaXIkT
Qq8uW/Nu/DdXKCd4rIVeReXI8Zjvdb7BFIfrBaGs9ZImxUD7jHgIRzr+0rI6dFwOMfdQTDbrXSYD
AW6DABhSTbMjKUamMHop27CbKxDUXZDAM7/tTcboV1AypghGIs3SC3FnAP/A6v2lPh5ecnWyhOXq
Fl8Ib470UYFhv8nBGxSxJZtS9vk+PPnG9rXpySV87lY95DqyDjGELodb8R/7fL1S01pdplDNkbJ7
A7U2qR1C7gF4HGyFGTpM6enfc9hGO0xcdSbnRJAUsJyW03OjLkKbz/Xu1EPsDY58T/v/DtIsTj6d
IGZ0w4kquKDqQndTJTVq0SwY/YZV8H2wLw1L0ygPmMphKaBcXJM/giZOOgZ7pjh1BHseuCTQQkRb
nspAiUsf/ZjuxQbW2cOfUI3veWGUYQRM/Ti9EJi6iMLGjHWv8IraCuaSQDDc2W6bB1C0w06+RpsU
Ta0qAWSRZO2ksD42AbLTUTAwfljWjktMcMKAZrykmfj6i1ogrwvNw+lRjqyPABQnTC58JwZt/HOq
uFKbCTQfusSGnVwvnPinCDcSffgJIfusaNeNLEIy0p7IYztee9FbN7md9eTHVaF522RtaKHP8pSm
xtl9sBhzDYiDjmYMYgUte+o+VXdhec/SC4mYKvfARmAKcrebBEMGaFJRH3fdC5PjOSpD0DIQUSES
3bOn1ONt+5OHe0izfvRROQn3aBCLWAmAXHJ3LcLV1GlAyc+cKaFJazrOJQnpZUJIEDvO3PWryzVQ
N6QSlXKWxZf+estzAWCrXfRbq2wMntDqN1TEIswdpVfP8AZ18NY9GwNTNUWhzF1SBkROcgDU7za2
72o53qsVcAzCbF0q724q+DfhyQmNY1zPVl8lgpc522Qj7xAreAGMmmvK1orJymIHhFjDjyd3Hq7g
Fyx0fURLQONBiTj8EZf4rOK31Kh8pvoYRDa3AbKmp95bRJuei8YjMtIg9DSKhs3PMoLXcRAkyKSF
ApXk2PPm17RLmdBkZNzf9greg/w420SxCLK7O/cAsiK8nIg9mqkuY+b+Cdrz6uwBqlA1MuEiGrTh
p7zVxclyJw9LUO5zjoJQJTirW2WEqrCCZP2WXN9TfEya3Nd9dihfhjSJ1roBn3fsZnrzZEc6VUuJ
RFsHDI6ikYX2npr4iUK5A73dyj9vMBVmw6lS8HnZABMIPzRWX2w9askZfC8mTRqKAEtePJQDa4SN
aRVb2Pzg9+CV2HE8SG5vt1LLWQjcJ8KqNTur1xuKrcZEQgbNMLPVT/0sKoTvwq67Kx+SY2s21jLk
Emm7syDaC5rUG2MNkhgHqI9Tfk4CMFurRSSCZBmLFUOdpfuP6F6Llt3XbVre+XdFzXk7CiumC2NG
Xclc79VzyGLoIGdHbqGE5p6r2LvUXG2/gB6iSrREGcz4wKFqSO2Ft1KscE+A5G8dHDhBm0v5URJf
StSZjQjkxumuqYIl4NzbBbP1YZMWwieQOtpbRyWELCNNe4tEC95WSanF9+goX6NMgFDRLh0HZvuv
lw9ChhIBoLdB/FstW8dw62cV6QVedsGUTwsuL6w4E8Vr3vPEjP1yYkZ3wlmpkUm86CrMNfacfIqW
MPaoHJClPJapl8ntswgoD+XJe/VGeYcYHrj8Hzegl4jj3Q9j9iUwSr/0y7975qVwTomqLYbYMy/S
G9xLxzxEi/+aaBFLsbuPGtRnkwvNLDb22+WxkfT1+n3HV4y260kz5s+fzL6ifvLPs06eCB8tUKAz
mIVJE94F7ZUpDDI/cu8DXvMkw9U/OU0595P3iXcsHMWrgcorfvs1e5boEaOZyfumQu0Hyc2QJ7hh
6og++T1vc4/FAEV/sGfyMa9T7iRDeXwmtJ4IjPl4Dstahbrfi/CX1OYPvjIm6NeAHMz9iFA1Yo/d
WVRhXNPd/ivXl/aKAhvGfbY7HUKFU0rOKyEfJMlnfGmNDROP4HOEDCdkHkFYYIP1EOsbxbAgUTB1
P4LRwAM0QUeh7QZKwhQw3IKVmYjKtM0fdE4H6XmxGG+4CVMAXbXNBdubVWqJWjnnLBc3T+BH4M95
lrR3tGO5sBRXZMuplrTEWDijJgeCUPTIFZACoJeL5Y+ecLhtXYDwBdd1Cer30xnRvkvp2YlGdhx1
CAHAD5z4npHCty8Ztvb827RNCWJ+qCGm/OC39a+NM3uhaZF934JwyURDvC3K+7ZxBgnN9D9o65Rv
It6+F+Le++2IECE95yKORYdVwlYDutC70JqCxqMCcY50VSkjegnqjjdsVRKyfeCmdIsVsjoAXwJJ
d8WbKwbnp1W7EIZaV89Flc2SThxuDlMnWdCJfFFvha3cwJ2pgM+P1VfxudREvPvXtZlatRiEJ/lz
XGznla3/qps4gsvmhDV4AK36LaKPNGJXEk/TU/bzLuLENTFy7nPqmzVIXMrIMgeIke1rn4FmM+od
k+uvvBXe9ScrZdgSjUmsqIenoJiAJ/BkTMqhy29rt6WI6NszYcrotlcHU1uuKJQUu5R74fQiP0+Y
J2HdIbXeo3mktphuaEwfWBbrJNw621EDRZXAmACtYOc7sdm5cRXPE3qBjT/P6meQOtTAFEdmsXAM
w2eJE+nJr8t7T42nr+kosjOQUUQXcfcxsxImd4UgZP4LKrmeU6azy5LbxpVfLiZPhz4FCGv0vsND
+Ftz6A5+42c4MqS9oFOFFPvZ7VDogavopsfQ+3lNW1KxWS1v79pQnQqxFJCtx5ofl+neqDwKCJxM
2Y0VLBguM2m4DOHr00R0DkNFI2ODDIfNs92qtmhTD8U/EGsdUk9LI5Kol5enlN91PuUPt/xe2PKS
62Oys/rhvJ+4NCMy6INMxauw6/EPgv1eQLyMuAwexSW/yl08LuHL5pLYCk6cUUuPkf5m244I/tm6
8ntNHn5jQngSdAhT/ucoAVpJwUtlUrVALJhkPjVxfupLbDfI0H9GQjwfwj3DJzGGpLQrz6tASel3
piqkJKJc4UamhSjWkbU+QawdR0HxO2hTmWBd1Fm5R2OHZhYhkVL00oIK+ikj8dTLy72QdXZfiqfb
I90NvF9BNJtDiIXwg6hQlYgqUrubtrdsnfudkFHZ3Tl/uBLKUU7VN6gfX8ODo8gNYOD6TGbe8ANI
8ORru5CPb9WbLL6BYCckbUR8GuZlfLXHPneyWo1Xs9Zj7W7/3x/kCF5pRfg5WmxqkcR48tIAXTUu
Xb5C0uWQsWJ69DDQhdLp2NQtAz86KiVQh98QSkDBSxZfLf66cZR/rm81dJ+BXsxfcuncYJ42cfNG
0STqD31RvuJ1l9AbWClpGvhYf2YBVp5Rz0Y4zuS269hvLrv8ZcAMZrKzgpy6M1tTaNyNPMXeF3yd
x1ooEEfjxeQ9ZuI4HjHAon2IzQJUqZJ2WCiatwENe9E5xgYI4bVDTCHeINJsxoKAgKXCsA0Ejcui
EJ/mEN2VjzLaIMt5yoaETQ8I/E3h2RE9QhNjEVe9rRU4nr4ysQ2eWti9vcWMLEqN5yoRKGUyiUzf
ftTGoNoqg10FyvJ8hPmatKzK3iSjcOjH4FJBMnyNH3aeeEYOM8eg2oF6PaYas9Ux3z6yV3/32R+V
JSpJLm6g44L2bWNs05kGRga2dq4da9ePTdQOdkmXshyTlU6xmnDMLqZy1tpWTxpxLSBrtb5Vwwif
5BXzpfyGwKGNVgyIUwQn3Yt5pwql9/SLLwhrBYraH+J7DGZJvyt7cHd+2PdZJ0nIbBFQG5q3FZhC
euMAxZeGRNMvYqW1pGJQvyEjw+xx5XHRo7hhidjTYKX+4OyKh5Y/UDbDO1KFckDxGVu3qsNq/n2M
JpBVHcl/1BurhI8htGUaBuUeHDggVO8q3X9Tgd5f/FWMV4bYCgzlI1X6gNJaWWZRw0hhPU0lksGw
7TO8Kwk7ZTBhKCesEZUkWVGTCMAlB29YuAgYscRgWwIRjhz7rhh1eokaK7w51nFjqNoRlo2oFmsa
zMLocA0V6p9c82wY+xCbuG7AHaW9knrHj8yqTYgg9gs7yXIYTFgIpx7WUWrnwr/PWyAGr5YFtbSC
zSSdta0GNqWEls68pHAnrvLyv9UfuAmWaZ0tlFYSdV0l8lxmGYKN16RPobT3lYyeJbsZBVkEHhWo
X20CJwV5nyFtULKQZjdfKu0HsB8aEp5ke5KtTUE5Os7l9OawWnRdPOEm6W0TggeBcGM83Qp7oQLR
Ngst4LJxa9fcy5VcdvbWHjNvbrqGD2D2q3n4Cv4Wzd+IDsn71Kffzo47Q8cr8yQgG1RyGNG9Tos+
Yv+QkL+epfSoB4c+khOwc8ejnVRf8X86iJJeSH1Sj2zVuIUUeooAq1b00lgKcDyfUwK8IGRrdsZS
vI8Sbe4/R/jS2Xn5tYad4RcccKbt5CQ8haqXkQ+znBoXVLJG0L3wlEsdygiKennTL2yKOdLVXLgd
3KDdMpL81tWpeBNDk9NDny53I5pleGOLM2ksIx2Rbysyp9c4dbArcl0xReAPcE4ZzrXvvu9jfuBR
sIIy/f9XaodnjUkrNC1v3XkHmBUClW5fwvLqhnFCC/jxbvKCLU7yYFo29Skcq/qyjCOzZrKmslgS
mcPLnv5wU9TIRlKyXZ4vf2sje6vuQ2s6uc33jlfQcAGb099gH8PZz6uZeYsknTNuFZqeFN4NX5Sj
+jQUPjChISnWRsviWFgzrhoOjj/3FgN+ovgiH0zd1X5k3aQHv1hhIOxo/kA57f8NRV/d18efngca
2lyZR4fvVFHQNF7Sie13z3xMGlBE5BY1Ms+7vPavKU5XjQ1mH01Yck7dOZVm1zV8gTx+6vhpywRO
D8RUqsx4KRuFimZ1WUexd19w662/6E4wNm/CQlUaOHonMd29qFkpdoRSJ1SMJc9Ee3et/xf5Id/o
85UFldy0OqP3l1sOZeBHTiE/KAx/TNNi6KHWrJgLN+mh8EQLrAU3X/UqzluidsGpKN25yjqF1Hbw
GcE273xcLE44CaOPQ0pYtTDZBS51vqIfhEYn/OgUHwJ7729bVnFxPSvSFmnl0QbXu09oWF1jBuLU
F+983pMEeA0KHw+5OT8k9y0eJ95qGPn9Tzl8PJHjYK7p/mPfbqlfrWAW6f/RIn/EbjMlwyyX6Tm+
MroWGDxMTsNYC0P5WbRKj8kSVlyxwhdp8XRiFbwfH50YvgcPC97Ibx82cG41Q9HOB1RZ3zh/dBTT
N/g4KTk0WkSBOwlcxYqWMBxGljYVBiFTVU3+GaMWnUGEcDbAkWXzO82usWztAU/4ZiEFqcOMAg7l
SEJtMjWKEfCrYcHwoiWCVOd4jB/jbLE74rzZdc+K48jpL1J3ikKUCDiOpOOXPx/r37WJhId70SHU
510C0o2dRo8zMHiSnIuFoSbOBWkCruPEpjHJ536cx0z+QooSYasBUDvwEKqqkTVc5jZSvE8B4P/B
wGD+DC6dQSB/lwEnwHHrFlNGSIB4NtGrZpj0LBM3mCRXNd6cDaivMeg0F9Wp56/5pSeX033YI5kZ
DbvZ+n1oxsaQrcjxijvUTWxFaeeqnlr25Cz1TQsrEBgN7kJLwOAw8SKKL7PxFXgRsPta3gywxF6J
5lDKYYkyZ3xON6TxdtHI0VH8hFKFGr/3VgyYLXOf78DVghLmKREXZvCy2tslxE+U2pQd20DTFlZ+
3IDzMxZFXGuj1pz3oS2KH0yoOnmzxHDnHtzku4NVTNWOnYCGtAf7K+vWu89rumAE9zHj11/SxzI6
SO512Kcc9L3qnZ5uva5XNsDp0a1cnLZiuekVqvI1jF1RH9JYKgKz1XvTjrEPOw2Mimd5KEbRhXRQ
yh+mYHYjxJ8OKayHhx/N2IjyiyYqy9nBNNITYV2zx8EQSXvmyCL/NGHDAo6fkRJZnqHwIQB8RWvV
69+t7efyZt0wrLRwTi+Y+JcHbTRMzAtPJYG9DVK8P2bJUSBarOH5jxwMjFbTHe7tKbphdNtLUzsV
inSuqKStxG2d8RnSWpAICMVxmABVRJGk+U+KwI1jk7HNA4HFG0O3PF646rPrpnvtQ4sDMdRvyEPB
Zi3osc/ks1kJ4h1bD3PKLRVHH6xhlmplpBeQccepYqpuWdRrJTNHb0aOQtUgCTQXOAq0ub73vTrk
8WufUFX07sX5BlNk5f60xv31tjBBfUJrAeZfjjizH5AL9v8R5IzXog7fqflKswaLgqpJyesEvtpf
CjTvWCKywzG6pKgSPAPyyFZPWCYPFoEynPL9UnmrRBJ7aO+yrkgvS+zI9FmEl1DbOydrNFNqb3eT
VTq1B4A3dMb5an6VfZ0T2C4jCHplEiqVLtuodZWhJKfmAYPr49fg4o0z8E2dDT9i4pvpUa2QpOjB
H/8A3WXwHvzBVo/jZO0szBnYX5wuORgT5mtpfZjvFDfWDuGTNrXvdKFwFEoc8drBg28YaacckQA/
9KF5Tq1DpyxUhr3gZDtXfBtF2CQBTaX0clkGGpwHBK6lP056YK4WBlVp/teEW+z6TjGSBmYglO37
rLWUQzOz9TaNRFNZ9eaTCs+CNYD+aRozTObt7C1SHBHVJD1VDcsNRj3Evkw7rMWbqp9fqbBvyV9B
WMIGA2iTQ+EhSdX4j5hyGWJnZ2k65zX/x0oZWoH3OICUjGcY0FYq5It8iKzJE9aLmAjrw7gK1Mel
BU2+pVu2iN+CJhoHdMc/y5KksABdgFrtvrZZ+wnFGKe1dnWpKm0fVRIVutOd9OUeG6aHp/nq3GMj
3zk7NvxCZh72jU55HcXAsxC5yMxF3dLITAD1hBSrI5/l9NjAXceybCaOpFOhTZyf6Q83KvVfNIGV
ggBRsNpnBHG1kuUAgYqlxwHE1wtNxfvTHgkHQWivmzcEJDa1zls5mXYc5AdilZyd0PV10GVXZ7Gn
Hw4qRplycKvFh0qRmxJGYnsRJGHpUjSZMH2E15D3AMP3H18LIv4jbN+3UilLqLoktU0uUxPGQyfZ
/Yepw3eT+Alk3CLU0Pg0TcHS3n7c07Oj5Jh29XpMR4FDcegwAR+dYEKcBln3cSoNdSvOcAqMBCQb
vydsYlXtfx8fVc2rpUTnSs+4wRY2ouvu3Z8HoLe0en0ioHjQC+qNHSmMqaY9ddsknuXxfuSMrLaZ
erKWxpZPwoUCmUKNxIw+yxZVFj9BW5JQfNcBnoboSasTlR07JX5kQA5sWbrf9eayYHyoCPkL9Yf6
Xq0RgE1Rtx6OfnVhwEXGNQbUKcJahruH7wH1LrtR8knHKL/jNA38krx9EKizE1G3ERpIM4GShag7
rwNNkLZcV5GSVn2c+Euoj8in/Ey61jltzvzYKAcP43rnLrpAOykb/IRUBECnpCfYfM+mfFe9/Ubm
bHWvbrJVveHEr8ftDyDw0qEmnrlvybsTK1MlCn4SbNOOLlq1kgl326WBR8NUkp4pcFlv/cNACeCM
hgoOXjSULVzGJGSHL94Sq5gIMxFKSgd6ms/fHtqVPoifupZO1axu3N1EhJwd86puoOS4+l1wp/7D
KXIyaUFR+NeIpQKZBUzKOblrTOPMHwbbs8BWvaJWHB+vQJA9fl8jNn8DzRqJtx26woeXx8m36B/O
sBtdP9u9abdXKiVGrqZi9VQgeWIF2mnkCb8a1/BlorTbQgb81CQYKcY3jd5qKoyXD/wqkHvgPuCd
d4y52+HT3+K5I2S7hJKw6PArG8BhCCdxp+WIEA/bB8yZLFvjvv18PGlqt/o1+tFkIvrog3JK9pZs
SjhnP5NXwYWXNgCMSH1GHrm71V9eLYrnLW0Mf6cI4sC976C4ABomZe/fgRO9qv+UZkLbqWA1kIAm
ekTJSzn8SEqmv+ser1NLh7yM2KL3h/xmCqmoQLQIYN8ayShHBgEUXE7T2chOg+GMkAKqOy9rhPho
lJFZhb9HnTzZNTJW5gE7AiN2sq6ftRLhbmn1xxu/rGGveYOM0IVOTw+mJWLi2d0mGKEmzxibohTv
IsUxFjIET64NaTUeX0yN1EA+E7rHHr+3aZP3CqxTtRXT7g41Op/YBHy1J+3sQDxVYsvGi78OSZn8
e65zQTmnOSZNZiFZ4p6L3Ouc1G1mEyFaH82Vx2bAEz8LMjNbe9HngDE0PH1uVkbFahann14VRC6i
P+4YdgLtnYpjK6ZtN27uehzDMLsLKEqCKBBs0b/7w/HyCyk4lrERScIcBGMIYxVV2YO4T9x2lVuz
bN2yU+BypNeuYCmbf1aK5yz7jZfxeIC9t5n7Xj98up8mPA8ZM870fgE/OXGQmSjB57OFeECkX9Vb
50ZQ0s/nH0k/gcsmezWXOis2Ujx2wFPP+jJrh28WeYyOjhHRKF7ZjY8C7UhDyxvQvjl9jvd5wOFI
qstOxPRyJrD5LVSw/w+DiZAk9/TadoDEOYbDJatIsizwMAlwUAJy2GXm/SmIQ2aV7PDEttInBE/X
VjUcVDKebfZNdU/xAToPVVOXetnPibwqd8NzuZeuKrhzmhz/GLP5dlQshGZiq0Y+lYxCyI1HTW+i
Mz6ZpAP/8BYVCMfkt9wcVoI/mPlbKvj0ABGZRTC1K7fms4+4XpgPAEKw5H3LGns3CIM5xSDxoEnH
NZ1Ci2rtJp753fdZTL/ptWJHcoD3nQkbp2PzPsTCtuaY37IADmjHl3WqU2gS14Fgi5qGCcYkYmra
upxr8M7C6S/RqoXEvzD9/43moaoAAZECZWekYwhvhBISU2fRE+9bVJrfpBJP8W/1Z3NX3A8gkAGA
0WfGzeI7opGeleqo2+lP7pjvD36ym/0vFf0kyH9mf7lIhZuTwEzCGTRXPSx8gdTTlky12ziwQRTX
iLQj8gicV62B8qaUq2/Or/Ad419VGasxIDPm/d13USHQrIc4Y47WQbZNQq2BzKLJnCy37ETMt0QJ
TH6ntROarW9BZsXX2KYmzlGhqB+nXexWYaHoly3U3IXBLUm6xtx5+grg+9z26oRb5qjA65dbrYPJ
KSnHdxWo+f/XU9nTW7ANO/EOVkYq/iVpmSYHibJwsoLnLPNycd8fyi504vTGFH+HY45ye1+qfyDx
PIN+XNrLoJ9PGnJeI4ba5tZPWjgfAgkNGtpN2SJsNuryyGJnv6yesVdDcTpHRCTFJ63Rs+MSi9vE
OvYgvNsBzt+qYyEY2+GnzbBlDJEHtcjSyC0hbm4IrdjRHaj/fN48nLyFQ+6g1r6k84nUaz6Uoreq
4kUqAj/aEYNU+GU4IQvsg8g7XKDHRS2AmcMXNVNOIbYKw0AxDk2IvgHraeHKhiMmoXTyRqd2vHzm
QjRlYvoIFFH8R+d+peIrfmVWqbha8mJggrwwl6QftUGwBfqYvs3+v0ozkebJtpohRUN2jRSDUpkM
tU0qdlDcwZcF4XDq2IB/2Q8FhP8kOgM64Nq6mTm4kBxwzW0SiY+M5jXUqj5nP0xEsnZNI7S0S7iZ
/ZlZFM65wtAay0Mt/oyrLTf3tWwAw6P/eeyCd0zCkVHlvDeet42lVAEzZGRHRVjFE0OCWwk9ZMEy
Sdnnq8sK+GYmfQtGlJQPNXp2nrU392p4N8LJBPDIO+iM9Mg9vQD4XMOun+psYE6WDnU2fImRqkkU
85jg0Rkk60v/l8sv9r9Nop3WiwwWVtaDMjfjHN8xLK16b7AlGKdNnAdmrgvXx49aED4vi01wfv4t
4mtoAuvE9lU7YvkzOPWRxZIYXObDMv4f4KbrsDbNB1SX4wVXuFMI87ELJq1dn6bnsnpQ7OXHIsX+
E6F0YutakO0CmIs6sE0LvTMaY4eWeCG25l+pqYM45/fXRPA8lAMzPxglIZFBnACG48x453fk7psG
T39tXfU5SPzts2iZjIU+pTdvwpVaxCoybXWhJQmDSEfbXkOKi+Gk4T5CGxIWKMNr4z5dWCnDmOBN
WZCWxOYYb/GoDM/3dvT+sekSJalBYG5kyWwlOimkv66v7KXefuydcojPhi0E15RnjP7TW57EJXaW
QtBZEmCm/8cRjUVBDOpZigMWLtD4m/bnAVJ+f/iE61I9YhxnhiIx2TUhoQW79vsuHktE/EYXEbwW
jxXKruvxTrLizs15bk2rkcbcbF0Di7At9lVwpIaIopGLN8Dxr4D05Thj17gOsCMfQ6EAis2k9sQ7
D5v7QGPq7CycO07dDKelPsqsGD2a+3MAIj2OFy8BsO7ire1BW77Wipoj3/1MUtH7K0/hDA/TkTno
4p6V91A+SdOp1+NCWJPlLiT0PjCsEHIDIc+yuUpsNyTgfKoPhFHtezHpbzE0PG4uQoUlbyW4VMgi
VwBwvSByqj8dEDgmiF7Tkn0B7GydYl6O28UH6SZ5AXcPfWnRPAtunEjo0yRnL+w7XlvaqhbXu72M
+KhuAb986uTG0U+JGS8FijMkFQI6Y3HBgB64b9w1zadHEFBZBAagTrr/BeWqvO83zhuJ29VIBSik
D5rfwNCs15VrdpXge7bznpJjsb3JmYotDYC3FwbO9AvCxtyOCkQNPk5zsLpdpEiTUpE/13hrPVGY
JJy+yPX0A2pfQboyQkNjVYNORglUO+l9yHPkFHcX1ZhnQTADadtDPQYn5qDntwpnb1mG7jXbAqL0
cAN/v1vNmAQwe+LPQLIPlXP2MonAI1kVvAP7Qdeyo1QPBXDJQ0H8mGqOpFWHkuGcC4eYPZ1PjcAc
ux4Wy1YCzN6j1kL+kUbYS5peRYpOqh0QbwDWWCGJaNnUxhH/NQ0oIq/S1N5nbIeJpBMI2UoKpAoL
rc6cL4ks4CHAgRFnzicIFt11nQE2Eq1QFqV9ulUZ/9yXz5KChYGu/YaNcDM2kbyD+89afRgblCeB
OwuB8rn613IfY1Y4K2bEloDxmVeFsdfiFBJL2pA0Bi/hTttEHJjLHg1s6zph7VW3+If7Olod07o7
DLF3s58+xvg1V0nRrWoUb+kF7jTqvztbnA//BzhxTq6Lg8orcZjWWKOLlTtYHRLQ/vjCFOEotsED
FnWL1P+5qjdhl7/wu79gUDPv9ybCIJfdpNqXsooiTEyTrY/y34J3DjUeXxh0PdcwcmLRBFqI4eb/
9Al8IX2KiG/kqg/uqbPpVUGp32q4XejVnc1TKVJnrtwcwJT/KRYKQ6XqNMmRuCddgVn+sJJ9MGHM
wEisjFbwAbFMTwU+2Rc7H+dzy51lIXZ4My/II8jHDsFEn0iWk+VEmezzpmn+BPLdVHgQGURLMSpy
rODXLt4eNm/OJWy21hZsmMiTOwRI5g8bgXT/G/1wt9Q8mT/aZ1blXhEjt7d4/g13Jln27VQsPuM7
zCrNc9PHgoPer0iVwtjDWQI9mBgDYLSh3XP7mpFsDf5YTqYMtAuK59W8t3SZF7OEw94Zjofhmq0O
duMQoNJBKqTiwE9+DiEPWUPcHrxebenCxE2CmBYNjcZMo7Fj1JPBzgIjAZf8anwtymFyt1sorAxo
ENPsjqRsV83YT/hf9BtYP7/AwjgjwDJV7D93wCkD8Fww0IonbrOAwBCqXET363tVlRMVyeWbmMbU
f7Wh23FCijG7yaTuEM/sZzg1CRfKg7ty3Nx+Hq8v1ZFWSuiM5tyP7c6ScCDaU0eWO00hYxPnP6kI
yfLxc6IYtEQLyQlQ3ci7Tv1F3y/OwJ0xpjt161TkBEJHc4hBV3PVEq7XGfJdCmJbHrVnKjUzHR9Q
vVXroGSMS7Qcc6f1iJa4LUywNoSYVvQnFt/4TX2Q26Rbilo2B5UVLPPcwCj5jFZsRv0xhsfHGl/N
8guS/WaOYkvW3sUfzbqrnOzAdOAN9WkMw9IK6pnmvaEdxHMpNNxTtc0yBb6YO+qjfR3cb+xllL56
kJ5wRHsk7RblPNTg27pVfuYLwattorTIVF/bzV5jrsnsuuILUf9+o118JnAGui0p0NM1yGO3Gfue
uuFURLzeeRdz8HldHBvsjlqxaOWfxzWifDLUJ+aX0/+LkpLUZleXtrPzLetNiSgbIM8lU3RzXx05
ThmcfPLR6OS+TVDTSRI4iWTx+Yu8shIyxc3iDYLhhWTo/0hN1Le9hZ3ikB4Zp41cbrpWNhxF7M8C
9b3mAdDBYbg5N1CzktmKAx6UQdCBE4Ao+EHlKu+VIMZ0Es0iJA74RIyo/3GUxoiqLdexPFyNdKeP
LXbC2CSzNbz05TkgBGUVRyHwYERqIBLFZc4TeNU8Q6UzyFZebmOM7QjBkwO96KvvxzMMq2gBNJH2
3bQl1yP2rCYGyI/XRJMqo3u0ZfwlY9CWh/Rik8MzgPT3e/CbJKwVLxKB6mNDKj1qm2KrJ4txEwoa
Pajf2AfXA7kNDWGncAInX4kygk9ptsJpKlcP9YVR+jPtgBll4Ndr1mcGMdDS+nz/5YHzYpXc03uX
hU2j8TZUtiCgcGvaRfwowmYFUzvEMMakj4suImdqBx/kDbXGLjfwVgD0op6OIJpU1qzzvLmtwIDF
H6smsjnHSQBjkhxPI/+FMJ4xCdSJiSI8gJMh186cT4/H4UzwkShqF9n3izAciK2UoBD/EyfpZIOp
QyxsX8sQ5GcvlaIGkXTBEPobLFHrT4llClCt9h1pBmWILGw2P88dtpg+mJ3GUSemT1EWSZpSZR9A
6zymg1/pzSboXoi1gHMPCwv8eCQ7ONSN5MwHSVfplWEghOQ2EPLx4lug3KK/JLS7Pu+xDcR7EQbJ
ngf1EpeMhHWEAvGuB7g3WtKG8FA0Owv8kc7jbZuVkloMbrItDM7hMSkk5O5sXXgrD8Yb9QrGWCum
nH4p5seL0Ux8UMA68amWJgyPb1L5qkAkfbixY0x37qUojBV+yzlorfm8vTiYPsDrrYImuF+vMvbR
K3Mp4tYarxRBjP5RkMW8D6TaHw+p4JixJdK38R/i3EELdDOfpmuZBWKhKqKJioRu7rzJNiVunJoN
F60y1xR/W3hhRLcY3J3IYTMaPsuVql6NELyyHFtsMWy+28tS1nISpvh0A3sJGOZ60uPdumo782Vk
U8oYP7T0cTJT6RT6QG8W+fOu1PQTjamEeQRZDI0O3luBPR/EZbWXDGbF0G/bHo4pzSO8R1sJOpL+
NE4ANHGkKXfmUEdwu6Wmms8Hf4aiICvzACRs7aYCq3z+EU60utXrZd52ViPwu2+LMYtQ6XPn5T2f
sbGSFuh1f9NbStgCFf94fVpal18qqmAeaB7KMNp7lLqXtQIVMAAzD+jlt5sFMptxcfRNGBjXEW7S
e3gx82/Lsw1AkHYjTYcRwwuxNtsd3Vzelo6ppr6b/LYGN+HgTcrPkIOcmZvIitLYD0GDg7Vp/pv6
VKGEzjsa3MCPrfbin7jPQ/JiYEfH3Iw2AoXUhbZd93+FJkOMGpAZhgZ8CNpyo0xnIcaWTOePWSA5
R0hlrILt14lpw+iLBW8TE2IlEDzHE0dClzKUkgzes9iVLHSU0oXg/vlIAEaWYjrfZwzG9gk4htaJ
ym646vyX48SJqH4ikKgPwlGz6Fe2Pmjzlqd2AI5ItnEzKtbrSv1eWP5IbuubXuYRHzR7Q45orDy0
QqF6OeE9FEeKlOzeaa39y2Yi2SyYlQ1PjPLvhMHF4qKKuog2y7Ma4a7iibbPlIsRriGSM866trmj
C+EIHLqolxXdn/33zSffkwOImwXfyaMf07MZfsqITr8nZZdD6Gsx3ZrAnwozKMPKgeH4VNcnmcJk
RgscE6+uyivdROWPKMHLS37I67DjAFzS50Bl+tMB59gjgCA/4ODH+ydPigP/hDbMG4el+EOLLVt5
z718Hz/NNHP7u5bwb6U7eooiRGGzZzcDRIIwEvNR0vUSHTS6380hs5THiDZ8B4P7oIInvAKfnESr
TWZjvNHuEDcEnqMvWEpPbWcFd8ZMRZQ0GEVGmq/gViA8ENfsza6O/obT/uWDwa4uUwD0q3YjgUIM
x0MiVn/LzAD4SnpCYGbbiFSHGZFYUpdiyxAfQGZeAG/U9ORdVNRUgSgJSyRugMeIi1wbKvGrFH/m
kedwOt90+NJBx4PSZanTkKu29bbN+X91r5kjllMrtyGmf9k7QgL1AQtE0cS9AWc+H1iYQ+VzmgIW
6rcNdeIZZZ3MOH2VWluW1RVwqw4F8Y6IvSFprf4n2+qcG49zFw8QT7HhxqgVlzmVgf/Pkidg4QOO
vsNPDM4DChdvY7Fj6ZSd5MFq33kkqccfvV7x4odZcV78mP4Blg+hX35VMGVAuL97NAL31Jmqhn6w
9p5ZrkWFrESOR4BJRgNWf4bt7SDfm3+fjoBZUSAPjG4qn8XBjsyNver63UL6VbHY3lfncfvmzl66
FgIo7BeUYzUEs2RLCIj6lt5IULD74JvY1CFjUE9eSleGqSXTqXY9XuZ3w+dKEw2QETcdMTnzBiK1
FQ2yddnkILxk4t1gCrtfAZUxtwjVIX2hPdBrA9BH42GlE/ouTCigT5eF//wyQY1pakPWxadOK3G4
tvD01Y8V5r7AI6Of+cr4y4PW8tqYNvix+kJpCsrSLMXdVDFr7qRLysxgM4V01lq763Dyn6VnQUwK
20Oh549k9M2B8C+6mLZ+MhwDd3ozzU5kPWEXNHBkutvP2uulUhbWZzI3T0TIUP9FuGxdzgA5HJxI
dN/YBv4qD3Osuo7WmFTE8dWKL9wZgVuZtplbjMNVQp+A4IevN1NlVe6nFooUKiz0VL3TpPSaUwyl
fcU//tskvbokmZDppya47dW/T+hxOLFAtBp0SEjNzSE+0HlaOQhbOqc+EbJHJssy3UjRvMEaoChf
9fPlFLmnp9aUsZIE+Fs+cDy6owQsdh5VgXRKkQnE99RyIgCSvYhJYBssAX5bp0zTBv86zazaUg+V
dxSx60OC6xYEm7JE1UGPg6Mb6ygEqPbHaaT5D7T+IBXVw20Au7tEK9krOZiHZvGcJzX2gMsuYsqV
EfcaG3JnxxgQmc2uql/W+qGwkNuwEuUCXcj5Gkp13+2olD1DAMPDI5ss489Mmnt1to5RG+S5CPgj
5sPJeMsfHCPpeWLObJex8HxcYapaYVsc/OYUVJsBYLLMrKsrUP40jJzIIBcXRIqqgKmhQllUpI2Z
7RyToEAsre0dfy66aErNOQgbAriFoQL3HnGMWfgcE/voqp1unsSYK1qyvlH+UXqVUMLDyGs6FzUG
YsOx43pSO29Q9hWud3XSarAXliqykM7CcM4dK1LTbW16w4D8/DN8exHh3aSzmP0GVNC+ZuQpipse
7VfajjlhdixDTszMrQ1GFyHu9Asr0m8wiV6/+yHTgneugz9XBgpgupLHV8SK9IljD7xZ1ExvwRoW
0eJKxVZgJ9Y/syhoHosOyfK1g7Lcf76kRdZOY0t5+z3yQ79fIxOO2THjgXpBJkC8KkAfimAfyBcq
gm7vwB2rpoSwM/2Tf4GAL9KsrnPmb66Z5sUwVdS8uQSapDhKBjvzLHjoFYnceRvC/fvMmRGe06hv
LYAjaC95gG4ZCEGPMIrAdRtdmzx0WDd0iiKxyBLKWdzDZLBR9PaNmPVLjU+MVArjLa6FNB+TLBXV
7zs2lNkE44GMIVFDTci7UNm8SDJu3jvJxYrX8JZ0R9bXPt33krifsBEPQ5s7dDUcX9p1fJ9jnmAr
So+fg2QP3XyaLFoX/Z7nEFOqYwD/THjG9bvGP5zDv8Ycc8NUVbOnkuTHIsKS6HtyqWMpIQra4qHp
0rhCKma4QXx9Nejcg4WDwwGXnaApm2p6X1qozMJgsanOXtU4ISItkwtHTUVsOiP/Rp0wQVF35AzS
UjOFu9B+iz96WOLYvFCME0txWoSiy2vmHnCihKolKJkJHBIPIYGr1ZPqIcolN1oR16synrHAWZ5h
o3xAO9Q05etsIOIIqgb31WUdegmN72xHHvpEKHZnJp9w/X0JqNU2uPeLNV8DuH/l69cpTyRAkp+G
HKVZ/UgdS0E6giiAj/Sh33DYqmERu/QgwA4cHNm+Hha64BjoS9gpwmjrhdAtlugupMir8xkpd5xX
dCu/lclUjSI1xULWSr8LQWqSL2VV/X7ITSFrHCeve9y2BpbWgN6PPfoxC1FvKBvIbxSldg9UBp3W
8z3MXMk9FsP+P9mjGNPhg6rNqHsI76CzXV2xdemPijXVY639efggNskwliG4ZNXHL8BWFD8iMkeE
TScCJTNDu+epOYAJlSsdChHoRdbBS6T9nECpJKsXceTgoi1z8zyb7PUgnw5YpWy2AYJt6tP0KJwq
bLSEArNzRl+4i9Gyy5WU9glVZ9T6hg56Z8VZrboUGXdCSp8vRzHNA0/M2UyMNKsk96R2bRaF6AGC
NAFtmId4JF4vsN2mo0znfy9X6PUnneZTO61qEdjbTVQ/2i/jwMwE9Ugy66kb3vl2mbHCBZKmUuRI
lYlX2KWv3dR3pKI5uTQYZ2UYnsB4hNFstrlHRpYkH9bfscZL6OOeZ0AvdmiC+T9mjfEDXOr6wqxw
Xxg8fdALNhs0KTR/TzkcqGvu4gp+jOclNYffz67DMdrWyKKcQdGac6qeoS2gq1vo3FdgOybrSJGu
YRAyFNk4Wd6N+Cp2BIqyq4bpOVtR9L6K+slK9yPHRm5Eh+1tHPiPh9yRxxuzGtnaUzBJssdmLPdM
r2qE/PxhuOml23AdS+JcvJuzcoGjRVu7c6m9zpw2oYj/abe+MrOUL+8goDEN7gDpbhRyM32fZE8S
YpesvOfd1i+/BHkhuf0WnNMd9cPaimOxlJCObc4SYaO56zgkWYaXfIlsfxkB2BTrv5e/Py3RwFki
SyP/KuHzpLT3W9Vao4hWLrdXDwiU0ZGgAipAKkfli8QoQl4Zlk/zaXsK/PtB4/fwWsxte0eqyU08
Ed87tLa+NDFKkhTf8Md7j+xJefRqnpMFQzOmVjpvD+sh4Pt4EkJ42q0QOLsTSqclBcqdDMeMYqwd
7gFXanIci51zTdr7E1ZWuGmvdTYIa6/2U1s4ndjnLOYodLaB/BxNP3ohhaS34DrGIBCuVG7tZ6CE
HRVE9MiwsZ47XHyBAsEZEE2Tgn1oATCcCFVRI+erOdIW1nnmPc68Qrr2QgqMgiDyuOQtNQdle98H
H/fuEB3Z0q+Xh1HzGOFlNsRT++lMQJdCm74tc2Sxyulglu3BRYLjbPU1FY8CW1oEG4eHxwjvgqsR
67ImfAFir8DTjsL50DNPsiiuA7uD5SdvkKb2RKo1CyhMBp0Q/d46fdtE5sU2XDVCgnPULttc31A2
krje2fJgUTQgXp07AEONAFRO0kW1ofBh7Pbb+o2QUEf0HW0UvTvJFuewt1Dt1p+8DKkP9XJCys92
9Gsl2FQ/Ml9g+SNCUq/UYpZN+tDP2G5YQ2jcvOSTLQg+Vir2ObHV+Y0Xmsmap2rN3vWzdHxm7KQL
S7F3Om9zKBaha80iA+WDS+AaY2/Y7WSbWUb8t1AmlQsbzn15Tfwt+VYTLDqsSmGbXgyAyf3lcWXT
N7voAVnNWEzVAwiGc1fycHfftDFdYUiTAvQtn2G++nuAp7gWH4AaZ10ikUGbFxirxjSEkSihUJ9K
DbE+NlbXeJ6pA6oDhPIdZyeBtr5l01/dqeWGBtups36DHbPyNuWsjnbWOgWEpUZbk0TobKsj+EPY
/+oj/YPEIEQTYcHO+m9pze2752EsRU2ZradJ/NoLqE9N/V/CmuegeTDV0Ds7we3jLFWb3XKJQsXs
MrMwRPbIXxm8q+QBakBeTRmNbFDGM5hEbj6kTM1uSSs4VsV3PxOL13n1ZIWJ1wrS+kWp2/SHxvax
P+Vde38nZ5T8GMK6V9T9TZcgSlzOOapgWO1+Dw37nV4IZTIRHU0K4O7bx5K09Oc8Ye2dPYmtRGyV
ElA4kNuAj6vMUqx4YMATJXr2ubGlZMYsHLgBYRnBZKykekbkxrCDopmJE+cupJbIBs1NRWhmxBxr
eY2eVql8z1zI4yCNI6Mf1hDDht2OPhe+zlDaL+nEs2ERLXNwDGX0EXr0Ejheek+nmFPErv629aPM
DtZnhIw41zZdd7KmIc5IDfRuIxgLpbgDNE4fq4PsgDux05j1vjH2kShqbZ6hAFa+pZWJB9yo1aAq
saxuU4zlkGtjgsh/xf0q47HCTHe/5jptfrSHq/dtFS+E4X/aLDRWIoTRpOEhFw7P9iCr0MRnqPOg
kVLxUF8FYEP21U6toIuTJFqpZ4wY7ix3/GqcCvyiXS4FrQrtt8YLl7jhADyoNbE8PVZ8AyFjgPvR
RwYK/xZ6EnIBBCXu6+imd9fFFiZGjlCEDXHGFyF2HekwVL+S/TnSr5Q0hJtgjAD8Coxm+yFBI7jB
Bageosm1e1FtKKOOvzjKKr6B2BGBv6QVtuSHenn8J3AzFhHasBqDB/pPU2KV4gz/gGrh7xBcZkfa
lQjenwyVFDDSX48lLMJQatDfxyINFIoVkGOhjsnnI/3K1s/hQq8T231gpZQ7ZFYjLwWTuNdE9Gr/
LBEvd3tFREofv7aVGvNaBHac4KeCxh2ohXh9NIseGQ8KvxXs27hfpna72bt4bhlaFKXTFxPI6yZC
IeE6hjATSlGZSonixGgQ+YMkcGIQ6FqBX85WKwhpKOeW65cVf3ufS7mDhdk+koOSidx4Qzni+ItC
hXd3MrCXS+PII9PqF7bsb1EWv2Wcjrs6l6e5L4jhVYgVc0HbozB8zal5IZkEr7thDKqeWbCQ2BSp
C9mSorKb9WE/XxyfppqN2KEwR+kStH24+4eKL5CUulEK5z4TrNoJwH0KBuC+IQMI24bPU9Zht0wy
vOPl//pIbklEztX+4l8NUkUdaCsfYhmhWKtpEZq9luWjPB9LAjZ6Rz2p9c1BdPo2TTlu++FKfHzB
palaiIfLB8mMK6TTNriHWfw+VAOGCDdPVOcQYPPmF4GqqnGbSM9ZfP9pOc71iEAVoJn/nNST6wHe
NFwnCKv+1PozMtQhAKHcukPC1dd3N8EEsTbuHuZqL9Q4DTMThltiQHVrbY2XZH0+JG9dRLzeEWgU
zFY6g0TlHeKtVVHfeha4UR4LqSxtb5HgZq2x6UmbbZ6qbmCTYsVh7KcZJCb3uQ83juYyjcsSNtTh
p/v+VNWhy+dz4tax1AP6Qu4AJSOLB6u3P23DCR5+gneRFSVdG2PpmaYjHnlkQ6gvm49xMxlFiUe0
uMgTaktziZnFYJWuOO79EB19nT2sTCMGB/h4vU/VS7BGaS8EWBl813AhD5C0gIA1CgIJlLT30DkM
4QSkXfM/aDNwfkM0hF6XCTuFq4HttCWUPF2Pi800/7EF2TQSFBuTEsEBppgXgqA4kxm0wSAlNh4d
zUSnWv+/IposVKj1ZSuJF0a8cc4+cx0rG5JthOjXy9SMS4UpCIu/hLkkXJxzE0wZ4Q32cwpo1Ess
DFLLoYEDjpp4dPO/RfipuRYYKQGn2s2CTZjiNLBLjH/W/G6C/3qQ+62FLG4nnPurjnvsojQeT2HP
pdt4TKXF6xufonBBZFgxYWd8mQkLvsDUD3RruNgdKUrEpX7mEPa1wA4loa6QuUeO3ezjxrD0zLzM
qWnqeBr2MKp+Od4dxck8j02o8jL2LqCzyRtUXeOnl0vagbFSQDrZbhJuCPHqYMXEKiqdo7R37Pmo
tN69Jtsb06XKdi/pdsDUfQ2I3MKVqMKo2yYP9oOd/ncrXbrJsFwzLBlrFc2+79uxmjr+3R+d80Oa
lBkodWv+4/bphYx1LbyRfnQtzry3Nu2RRUURFnovGel4xT8GkY+upZomJ06qkXtdL/e09hDdzLt0
Sisu6hFTkgZ5iojG+MVUFYmnIzs8htWIudnzff1IEST4x7Fd6XTxOPmYnnCoXzEAWaLG9rt6EjvV
b/ugCFuBOXgQows/u/RBwMuB0u667cJgfkQnEmjlYpwCQLhEEe/PERxrXXwvK8ZHQOyPSxAhthbN
YSKKqWfRuVXgNNxs4MAdRHyQj6Ke8uEeBPJonXMUAUwdoLJ+hbEC7rNzF4utMYYM0zcxdSszWK3R
OemDuYIA86Sx0hM7rB0t4cRx7qDynjo4uxSW56BJIaerTHyUybZ4n+lRdkToeuwDRKnLzsvqjR8l
QWLV1jLg57ENNn8F2cML/a3HdTa8KbhqIsc81g+8+b5ae6Ao5Bo09U+p9JIXDppZw0uOyER52GMH
Nrlu/C9uwW0UP52bD8ZTCIJmfTTJRP5T7//S/j9XK9calkQWX5Pic5KcM4w0O10KRvNj+MQFEwPD
okducgRtnZHxX/4Wxu4RDh7IqMBdl44XkaJtYuN+ITn0BLm9dFy+kDIaPOzkjOn0fkQdnthrCBGF
WM8tSbBYZ+kq3Cmspx5DGqf9QaOkb/c1z4m9n5SSfu3HES0/TFL0ahfBAMKijcBBesJmBjcczOy+
ypHJW6U7oNKmV3RlRV+7TBl2P72SxYRo1NHuPZlBNrU0tOU9sUTeMe++4RaBxzR9Bl2j0wCLR8fI
zCgaTsiU4J0Dv0ge3HQgTvaLBHIBX2vs5ZeK/1s5sHnRf13HTHDclla/v/GgWRmbrryLPcPI1OLX
l7GqWVbZqYLMrX2hAQLvSYJgQ9wuBjfpKnUnpuDMkD4rgeZv3FISaeVZI2rZ6ZNQ9a+ngbsBjpaL
1xq+8rKF1ApX90FzL/emNUwsDLZw+okeUZ9/0Mk8YA7JvtHYWZ7stjfaywgwFqi32A7QvDxVxrHi
ruvwEDAhW32RR6pmqI0mzfank+jx8qZNzet1IUBjZ9whrlvzwSKOWV9u1g3usKvRecY7UgghxXHn
J6kPfD5KoyNEDebcptA2zANX2IdnNtyN1kdXWc8i6gMnPOBADxlvjjjJjsefK/Y/UchSftBy3j1z
9WHh6JGJHWhaWpzGPZy0reQee+ZTMudC62N2tScGXZ/HvaIJYsUBF5SQrqK9mwYJ+zLzCtc53Ru7
yQ0yPy4GxY/P81l5Bcoae37ykOdj7WU7z+0sNvgB/yv6ekIiLfkHv+cdHit9TR6e1NNR6Ipf9sS3
lhw5UiVuoQ4PADg/M8FxWloP3ZerVC6Ns7a7YD43tG8WxYIjUEkT/Bg8xCpM1YIxfwzqPCfUyPyn
3v1kkhJ24aVjNHAouWWbAi8VNSSQO6opdEJ4NJ23/hnHfz00S7MdHrCorA3zIBgrgH+M2ZX7f9rU
qhQUgQQjxR+ntWmSAe2NlxFYsjERj2BoCH2iHM8Xc/T8xqCCTIjYAzVgO+xgd4t73qn/CkZLnDCb
+UyyX2fP/603cqYk9P5XAOOrBfbCZQiJk1liUaNsER6CG0Ao+PF/BsUCAc5cAhf02k81UPckKNOW
dal59FX9eZKN6fPopBohuaRAKPI+VNSyo8lRAgBBeXcEdLicXfjptRat1CnX4h7DIw7RWnMVY80F
Mc3GuBu67gZfFZT67kqnRgv/pipK3Rc40GsluTA7aTEfNya1fiKusj1lulWkQmZS6L+anVqTSayD
iURqC8VsWNn6fHpdslDPAwk8RIUMw5WXwx9pJlU3tP+dGkls9onUwDVYRanz/tcmUqfHFDmcDAFH
Be8MN9l+LLZ8J+EMFYcJ5UAPqSJi+cZDWqTUrrxV9cKTOKvvyNtz33yS2zPsWD5PVvPDDQLVkapN
f0I++Hqao3e9Dv07jtZ6cAHuXtopqt12C8OtsZpwhULp35S+NyaZ4GvpmX2D/tfZfJGls0r1TwSt
uJCpfuZ8CVLOsAC8gf9It/6ktT+oB/I/I2xqcs+g565MPnhbh3dkoyeU5SB32Qjq6zJg6YforimA
PZ3lXbiUvLDDSG+AuJcg473hCRTQ4ap1bF+dkVIdxSd/eWACJoJ2pR4U/gc7jESXG/yD+qAT3M0e
jRCrPBL2MpzpgfYVhQgsdycOPzZ679hSWZQB/9C/ZTpCIbuRSV/Vj4TVHVVzpOgf0KnjzOoTQZfH
HcVUIFHp559q3Yn+FAubgXRaI2ODbJb79ftGZ4EG8907qFadE5CpWXZ//EsamUxNEuHwC1KehNY7
MloJSanXlR6Mzuew/kGnbyY/gM22WsfRD9lyJgRnDuRBzFWscqUhNnnekW7ckqy5+vypVFYbr6v4
myai1GWYRqXje5jqKZmGQm7IHqaNuD6Ewa6pdkj7EPdJy0ZHGPpuMAT1IHaHRVon6TgUGj1oCgo/
vSUlF40/HxlQ4ivWWUXrLSgtKPUoqaAA2Ll3qycEinv5z0EQcZWi3s6FqdO7HQaSMi5rJaex0I8r
D4Ru10S38DIOagj0EQa7R9tkMna1QKfX48MdyzM69YqxuKbn6EU9TT4nTHuG6RNKqPNKQMytZiy2
znm/GEFV/mNiUa6wgV9YmDeizkAjNzvxgrLcTNzjikaRJPKMy40EqiJQrxjjb/CSTjRD2AnDyp6K
W4uIwo7Vf4YIbQLZK/kzwDuSylWI62Xksm+cQYoJx5nnSRVF5UMSpE3KNdJIe+Uuc2rJMr/t7v9A
tDK692kVzvPhdUEOVGC8EpN2Hm6svRwEp708ErbtOJ20x9T0fy1TI+zcIhjIqsJLAWoqDQP6mpsz
auMVKHNMEjQe1PUbjlxKVzyZkONBAQLRPK4/S8YrR/S2HZSMPzIj2v84pfWgWXLgzpf6PaHXOJHA
ZY5+fkJGYoSHi+i1+aKxJ4dDB6/biXGiSiHEtERVVSFkP4o1suygJ9I4W2zTWgKwBSLO/ouRnmwZ
eZjIjQcLlAlWNJQx/AS29ZY07F153sub9A/sMMnXHOlcLj/Pu6w/dFnNpUo5yudFk/4GMh6LA4M6
hSFF2sCtbxXjvlX13CFpC+b08Quu8FkGGVTmNbLPXglyjG99uF4DThiME/G4PS3NCXbvpNHvtEs1
g35VWNTW9jTT3ZNDDOJSj5B0djJah7fHiaboqzv98tMnCxr5bZGLywN2r00E9lQfySfd3x3h45bv
wXrfwP2idWFk4wSIKlVJvp/5bzGyEIAwXXtxOcaFVYZ5ToF+ymz9B4axLSuxxqVSvevygqES59S4
9iSDrRvzFQwKH/SpcB/nGhvXl5to9pXa4QVd1oHPHysF5q8AJgi86xTVPZjXb0yetTvZH38cMlh3
5cRL4KvS6Bm4OQ21+UY2qAKRuYc0q5rCM+KvE/3gd8sygpWtMQt+occ6pMQ9KmIv8PV3P5R6oDMj
5gUDomhcJbC1yTA8tq2JK0eg5idjX0glV7F9GuywfwyBg07WINuDZsu3TGJtdHRSdrzBIoe2Q/DY
IjzTdkBaAH3jfCLWf7urLYHJMDTKmW5knn/9myrC25b3+u8bzEclVDaRGOyg5HTI49fYUzw8hYXp
BBg05dF28NwPKTLkHYJ8rWobKXWuwowb/2xPudS+4Vr5Ah6qcZwaGZuGsWJMNvgzJ6lowE7B3UW1
w67W+rSmHMB/B6X/5oKX1LxQ8lDTlZQv2liwxR/DGQtFb7LYvyIUAYcuLe6j3Lbl65LTQTsusyp0
5RmMKq2NlLuasxrL9XA/09uGGn3zB/TWGaG2rdaSt5Xcjdxz9qsp2/QUL1ITFbgH20EZQWXhQKCF
qoW5m3md1YH2F6ERvUHPLewutOmFuWQwBnQxny+tBjZ6CZkGuKiaV88txH38yCUFqRNb4lB4JF9L
huCZFgQCwwmxzfv5XJpX7lUT8HAs1ozMyjMtIUTyVkwVC9Il2R/67X9OM3R7/NgAjHUZdqpwPfXy
0Oug5as/YNib+sIDqpWbyM7KnQrFXIRSiF7naRBycNWdY6hgg2pX/P1NCL7+SIL6On/QiYGzXEL1
Ri0UJc7Wgg89NXhdoMxl2ftuusDUybnegmPqxxnwsdSxsCz6B5e9iGqVXXjxKjaPC8+jaAahnqvE
U/7sof0apeOJ97+msnfKUOJ97ZIOneJOp8dSGQ4Mc6vL2F1yo6XnGKcXLijhkrWdWwZQKsgFLzSl
Ma1t0Hk37oqHj8L1zaz40AzHgHifFkqB8cWQtEVQevwJZh+OREEkz3mFUTPIebNyHNQifpWS03RW
7/GPDyxtyLLhg1kNKn5+JouguViu0+mH6GusxtXpWhHokmE8cCA7zFnraMBoD+54aZCFI4aqMmA8
ZLLcVF20V36mf1m/EpnNJ7bqFLUQVCqE4wfCmAaNXs+9byfFQK6612EhdLDzXFa+sx1L9dlal9w3
NTG3VcjSwzWp2rxezQWJwa/jig41byhUasgYyRUiaf7rYS4SffYq15dFIgKeSw8FnRFWD22Hs7WC
z/jPzcj4cnMlmmjfTWtMtNyRWqLNGmp/REJYrYbj6NRAgKb7GWLSWsn76Ms4qeQVvH5xv2g85YHk
qOMsIQRqwhHFDrwszPM2q/icvU3lKK2tTOGFrzxVzCA4gmNo/fNYqoDDyjnGnulYSXDIbzby/T0C
O1GM72UivrCMla/kq/wpxqN/t4WyYgEIaUqDoNLUMRJ+4niqoGnvHVagGN0IeMfnR5IYskwlVcDC
3iPlwsiwXTdCR569tj9vtl51uDz8qnvv65K1AUghHUQ3vtohogoJFLR8gllqDdXoaQVlusTt/heI
LJ/3zssDSAAc2+kIxh1MJtLD+shJsXFSlwOz9h2lHTQM5EFsB2sOGViobihYt6+H/xKzJDU2PS2u
fxdbDUrJ/CSdE89NoXiQB+3zd30kKXw3TKRmG2RoIroPBAdoGDhbG9HvvsOWVUlxe911hvqDsnCR
jUUHEVWRIGIEckygSM/kI8g2xfzbBnOCfMXQSD+D1f+w+oQ9JHf6Up9uAaCGevdIH+vk1EIyXmtE
4i8FPyllJAr+xNT05yElTfei/1SrdTz984sBU584UCk9sQZhY8rotXZIWBzsvBsRM2bSRWu1x4AV
8q4Y0LfZLT64R7RnhIz5ZHl/tF4/E3LC9ToTPtHq9AqsVIKwrdTjmbAyiAUkADIrRuDOBrbp678q
zUOjASls/fjV4BQ+Hgsql+ukxY9HEN2xiz+LVYFBOYz9q+JmHA3zM/mW/2/s/YAfQCpRot9CaHmM
4wo5CfVz9slRV38c1d/XEW0UzecoAxPzSOQty1pld0Slmt+TFP7Ph8cr6dDN2ZkoUlEHBNMf+TTk
dAaItckqpHR8b60Z3mLdUO54uscdvM2NMbdP3PhqcDXTZ1/th1EROXbshkCsLDiIsSURjEepwRln
2RcmqmpgE93meLLO1sYWuiuHoSiXAekVXifjnB8OjCy0UrxT83sV7nsZqAB4wy5BkBLGME8lyCK1
nIfVE4ohw0X+LWgLV4etCAfgfy3aAvXPBolWO3ADk3x7goXwKyDEPPVbSZz0VbpPJEpuX8839ncq
uVOSQaxa+XTJslY8f9ToUXcQDk1FaESa9Okap0/2SkHQKfHVEjICSuHcc0VZblfb5eY2rd7kTbFj
6RC/D3BYXW9C/+tPF7k9enxPqaQCIA1pyy2idniPLA4WEjHShjTqCIEHeujELwFt10C2hvP3YFxa
alkY0qatnGuZGfm/7pH6B+I6jaUhffYdH+j1fSk2bhBDtv1MKz90EU1HckRSaxkQ3ChaTg0INmDQ
22gnBXxfmV+AudiAYmjot1apwsW1d3hSxJzc+CvQwGPbDOOMakspEvZC951HdlCBngza9OOMj8Ra
wzBLTZpG6QWNcVA7tGXqImsFFjECbXlrXPj4atGOmfQuPNLl1Z7iMtdiESRuQDFQGwp2vBZ4nu0C
H0mXR2ABfiqesVUJFeYuxo8INB3UVv8r3VqRM4AYnYVGysm4bZToaascvHFji8DZZ1/UEviNFawi
B0efy3QNDwEPCllu6k5HeE3E7cHg6f4XS94iIYH79PqKrQbzTKh0ivlibiJNdYPdwYlbnznEC/8w
R1DaSGenqPB8fDCODbmEgYO+Oc7OoOf8OLoQcujsuFBkRS4+FNaO7lTwRT/OfEHEO20IXifMrUbw
VTRLQ17c9B9cUnYGTSrLYfUBN3KrBy1exFK5mfon79/nvnfDHpORKbid6809oQpRatYSAQlD+PD1
c/7/ECQEx+p6mMT0l63EWQ67T0T1Q4f0cUwjTr922BT/39PKD1j/ndQ8Sbn4IymYnMDZaWhWqe66
hDis2npLGAmWU0w9yHl5WgF84uDp+FC9NdZfasVGkk/S2L97iAF3Q6MA8L7mp3owgrbO5+WJS/RV
3M0lWG/QVNmjGoKQv6/Ek07Ku2eeA/zFo35lIXjLA8V7UjiH4wVyhdmvHAEE+vwUmbXOwnuRPb1X
bkOLAZ4m2phgX/fh6o9eGI3TKMUQP4cNvpMe/k7HHRgqAqmdIiehjmdRsuJ26w8RZWTlXollLc6C
Mrz2FvCS0+BcSbiSyyoJJwnNWBjQTWh0n5iCJ4B/cWP+bhJG53xV2xH/oMKQXh9D+kaO/jDjavx/
pUW5DicKQh4722SR7+iE8EO0nuNflUxq609ZqycTLnNh3QPLH2WyxH/fVWGrAw5KR+m+Rpq0+qua
rXjec/ecJwqQDAoUaWTpagOe0oInMFgrTehruaDup0nr4IQuMK4KeAo9bpPQyN8ASU4gcBQgwlBg
R5JfBYwYX7fHuRzchnWlzZuCvCjZ2xaQW1M5+p+aWtdSVEiq7jgLTM/TZmVUOuHaJ+BR9wF+8PfZ
NVNOLxv/tlJYCDzPwxggtiSNnqBExsn0kVwsEXxHLVZYZsP4Tk+7VtAGaowaf9T1VLgakseITsc5
vqK7rP4zjFdzkOC7d0LAVg0VVyTnUiogKvvomTWIpwT2sgdjRQ7zLKlf/iyfFI/kqO/TYvf8McPE
rVL6TC+pRhl81l1xABn2NX//wIQ8gcsQ/2Uoq5GPglsZku/FI0nOKnnQlgjQP2u43kUeno/A7JHE
QWKDw5ZUvHHIHWbFthQSGjrYWnEk2VekdewXF+KClWKqr+MSfb4MfSWK1lWMbWJAzkzos1lQ4LnP
7oPK05JIBspJjGLfVcT0G393MO40Gk/6DzVjCIW5il4RFFQ44Ok0oBQiEcA7znnqqjWVln4lMQcE
Vu9buiJpSlchQU4KiV3uP0hQPZ0T1piogz20VaVkO0MhDxHASF4I0CDRlDVBSmpUZGTeqlhIpQOa
hfljdNsxsixhMSgCnFQ70MpoV7SoEfFyzFw0XoUl/623DZKikqwz7VVxISqK4oBXODK3GGURF5zj
M9Hr7ZRTRMRQxLHZYReSQ4E+gOHpdCy5ZCLgVw0ckmFypRH/YEEXWohQeR0WbowmUeGTaPv/xS+S
2lwP5kiiCBbNuN1T+6Tc5CWTWRh7Ef1s4MmyxiMO18SRXdc8TBvBsI9Pl6t6t0Zt0s6ujJmGSg8S
MNUEO0GXmZwbzlCPdn1prWhwWJkozmeOTGgpG9KmPT7yHXL1IBMACSbHQVMDFoRaWvYHecZHN94W
gWzJ1a/cyqweUFXgSvouOaRWBQbvBP2q8/jrtkR3Ab/M4UZ6g5/gjRm10JMI5sdXaEyMWQVXgEjS
BUr2EJUn/Yll4jsueAo9IVfMzOkyHfobN7XMBGAiWzagq/PB1CDvPq3oOzFhHo0ZS7VqRFDUCS/N
YSoB78i+GIPmCgvmHFwAoVZuThZb0AsAxlD3hx91OaFWK90FKylV8xdHM1W2k+xvugwJi2MNecm0
eIkbeck8JmLD4GNmdhHb1/QKQSQ+mBDThIwbUdgky/h5/5vBBMfUTyYQbgNY4c7JwqAd1Bunv5US
1WREih5m218fCp50jn+7vI4sf7jkdMbT5LFDpWOK87UPJ3usGTHbB7YlAWmpQuxWa/T4O3V2YioD
Z/TqDputr57ZseZECoyshE1H6mIxxqcrwLj1DTDAcBL1b2BJcX2BZsxV+PKE0KEcZrPqE1L2VDVh
347WYTeVNnjRsEgP9NTlIYfeawW1JOIGnGM/fhDvWc5hthFUZDaQ230yiTeSmTl4S8CrSszSBlgb
CieGZLruQr0rhT7BzGBS5+7ULXlrwUzRCGCmX3gSU+OFOAA68Jbfpm3BORC0Qz8RCKIaOfaasJvw
Dsz6NWAYn/1zhkB7nZXM47WrlWrMVS1RQSp7PyKVsUss2BkqyXX5ETnACM5wlBmJqkeTWKcmoOTg
QTr4c/GPDv3wdnOJ5sZEgWpG+84oCEYHRCLMVPa/LeKjRERtDeVesIcm3dmjN+KqEIZN/uOXGWnG
UCs33Yin3HcHBujwrqFeI3zg4/9ZUQjzXKNo2LlXJsbURkqXXDWUuTyMmgyDmHoKRm51+3aiPggl
TlHE8f2/8a5qpbGmSnHGJhlxWysei/T81UiihxAkd34zKQg7FkazH6z4b2OK1UEo5hxqIiFC/Jr6
3c78SG5SWVoSQW864s9bGqK59md7I9jPwgTjUUziSkcsNPwE6et+C85WSkdRVFDL39+W6mhkvoOs
crWfBN4m3+Erg3jqOL05AFyvaOaD5OClEmuy8B7AeKU+UK0F3U+GZ8cplNo+p72EsppAfrQet5VD
Vwiyv7d/lJSCbUAAk9hZxzg+kGWRC+Ko0MeryB7iE31bnrK7MxT0lrJfdlGTkGqn5xBiTvv69TtD
vs48W8GWWI1HzpcR352l4RsI6nQRYrfYv+GVW+WxuEmbKLIcMk41PP+uOGpOVh2me1wI5gT6/pz2
HX5ahfUbdIrUuKTSK9nI2K3qbNs8FxkDXc/12gHjjjyzrAsxk22sLYSftmu9EF7lAwSc87oX/LpX
Iql4sdh4q4yfuLR3/bvrZXzOILU6DqXQfLg1ePvyW/Qs9YcvWqHzjZ54ZuwE7mBnVneCXfPtbyOI
NNlTdafA9/AnX5SZh/+7XCb9xoVNOen254hoC0jxSApi8wmALaKYqVyEEThW8qPX6R2H+KW826df
ZXfpikNU8HgziUuuORoD6oDus7eb+qY3XD6dJ914a0bj8RM89bXR5nyA0FaKjoCko2JxW1kmkvin
AURMFn3thBNnbJZBnIDwYj+HbY0Nwl8gJh2W6+AouVebjyAT1B4Zxv7bqwI/FsD1VjrpQyg0QJuV
Z7VSXFQVVq6T3W5dMnG7NgbQGrIe/nNNzDvC3xv9znc8ijmvlxGT5qboL813ned4AdAshL2fZhnl
X0XH2NuO3zXP5b4tQBi4cUFMeDuWD+KBW9XiLEwD2+HO91QX3iTfoMbhG7kisVQLP3eqt7Fx8zjY
Fei1AjNJ0bzYqD02RDxhvRjbmLtzojl0ETcYUcECaJHU5JoGMS+myxhuxmib67YsA50sPam+yFOq
HNw9k/GwXJIva24g88kYdC7Jt4LpLFTc8TZ6K2dpaxEgFKbp/2SVODWdPfh+B5N5XMTJyD/UWHL3
F3c/WGyWXagcZ3qJp5fURZsMM8hvZ9alfuaLnsJH6Q17BKbny7Xo1ifmSJDdTKCjtsjwlRBDToEz
PqsjNf3C7mqdBp61tudZPJylDdHMB9OD26T9ORiEkozoRjX72UPPFwUlGplsCA3JzxL9FFjr0QGr
w9W/O8wVG4zstWTsq0TDY5PoysJ4cW2kqZbM5bv/yHaniseVVfwXLoeHGcwVBTd7IOsDatawdFk/
XI7y/MD6mzfTJ3VadZxpA52fLTcLV6tNA7ybGYZORMqrk8fSK+XAM4Ob1e0xs1p3OTH6NR5LDgp2
wLmsyYXoyk3Huy1U/hNKxdncbxR/152eiNcW23keTTKhrmiElmlTid5vbVWVkTbqgB45WrDHl+Dn
JkgScO1JScApZs9ZicvWjITdqpllaWvYBz4voaZedGGeSVWV8EFQefjx5ys+7D43JGpBDOFqs4tD
2m8QHvxUrYnZxtatzI9NapaEx8cXu1i7NGd7FWdGVMYmZB8idku700Gf7McZBD9ZSoSIwg/J9xyq
ZlsB9ct4/+sdKbaOV+2SjIqLgCBeopPBhbX37OtCiEXdTu6Z82+YJVb5VqVv7ZbEaQ93xHyMM1lx
0EPPc12WsY5CexulY4Qeh+lAbsmdyq8R2yKAEBI4e2JEEncCK03GYXYfr8q5SXXDxU6128eT0ePP
/mmH5b4LG5vtiqVvf71D/e6naPOezwgiMBkj7XDXbQekTxJVWcHeAFz4DCVgNN4WK322LKYpDHJu
TRwcTatQXbv7jChQKMFwKt8+6aNvpxZg1Z1/QVGp3uyiTYzr0AZrR0OZJBHmDtMntUvW0K2k5Wq8
EvwsJvxkvn8JJQfZ7kKXTBBVjIDGCH1zBpmvmpk2vv+zsLYJHPeV6GsgFiO2qQr53VNWmsPL5Z/u
6arkq7/5NBy2lo23dVWzo8SHGZZO3gzXexuGGw0JCwlccTBlqBnVViSORe1adITusvWWUmuoGrp9
luD+RR+G/YINz4QrsjU4OBQpFnShFPEC3cYzxxevXpk4Dlg0RKYpdze863+NJSbAGu8sFP+iYUkx
GHducd2Hk+9vFVylKkiGxho1tg+yW1Tc/7/CAlI+mki80WXtX7v7qx1qyCepP4gUl8XBszh1EtKE
vxt8EgqvMJExcNobCcFH6OWeHnPeZQA2I6vDzJBylFb/k2avLAiWv2jlwAU/qEm8Zwbp9Rikyd+j
r/9PAyNgzDz+JHptTZ5SblvPdd2jGwWKlNbLJgNXV9pk+lJm7NvvEuPH+7SYX+Ltt/HNz0blmAYT
XTvfHcfCW0SSWK20lqUgjvQ6UWfk6KjAVYA6AKO1MduNbaijJnEcboGO7sx8a0n9ujQyjHJAfMwq
fGhHkjL+YTbgypPyC97QV8yq8eRqmpArdc395HUJcx4p7tjXqbLPdB1nL7gwcRY+6gEJ5bOT+9Hu
tBAIbQIbryZoPzuZeCv8fGG/d1DStWKRXfRA16frWDV32n976J5aRxeZrZJp8gBhgZaOtf2BZii8
2p0h/MFkgQ2NM0CqR6GI4HzIS0Ze/qjhK9RW28sTL2RE51gvmUxvfTUE3QkDTDZAUxyL6KewTU6j
WSNmMGYHUiZIC+pK+rmwJWjqorU7UKb1/kSDPsCkxMnSDZk+QrD1j6y5i1YYvlZujo241LNyF3Xs
S/hJLV0zIsxAFDd7ZK//AbPc0AGbcSZFHUtsKlPYXEfNzGs1Owv7JXI2grAYB8/PWEDDzR61ojNa
/gRvgppoHGPR/hEcyzsBk4loaVDaT6baiapgdgV6oFD8dgu++gE5HTRA8wNKJ7V/Xvnr0kedZIJF
DlPpN/DHXbZog9ToNG2/+98OfYyWb16187fr2npi5vHmPXILPAqNjDcHP5NGmBHoRBY7P//UzHW9
8Z4V1Upw/wOhDrRiu9x+cY7CGz6+xHFeMzZlWdG/ofaRUDzCRXcQykdja7atiY6vweaB8PRUBVmH
ClOcjtYprb5hGXZBp57GZ2L5jEChwbLEwDRUeE7i0Hs6Ph+iW4DElU67ogmKNe7xgzQOSAlZQ3H8
u+Z10eKV1tid20aVtgW6NKu1T9uAPftCGIq8Qqxaro+h0ftH+m96NwbsY46xup86NpxxWV/YEKOM
qaYMpM8CFJMzrB2GAVU2GYL0S/GKEeGb3nNDiw+45AiexzyBqRPanuZYpcGc0ZhkeXPXkvw6uF9R
7wOb/JOuA6zOHhKcMmIVy7celV5juOoxVZglfWAriBr9E8Ua70XxT9iaAsRbfuXigcZVMhq9y518
SyhSPcXchOv8qSWUHVKPAY9TMneHuFiEK/Xq/dEiM11NDplsqOGjlYNRGnz8M64G78tVMaKXs+VW
8V/iekgZm+EtpPjwjZNzYnnmahPcFIdjQafs4eS+IGneD4W0bAzxmahaKl+H0wdCK0SsxiAUqqqR
tj8UEA8CuQi+R/uKPUdttyn7PEaHIfKl8dhmyx9AJWFMA+0ouM0xh7ycLB+KeDlTDRLSSJExjABg
did5yjc+pN80gGLiUco6ILsMNV6MgfucvlIYxZmtw20c69WF6Kn+hLrJ/UmEi8VjrWinNWcEdZwY
hyWCLSVUvGcHzvIHFAi6fG3bod0SitbZ+wNegKushkENK9dYXRtBQl/FZLKNZ8VzXHuF4/s0O47n
CF7mGXVjqHFCDrOWWVbabNL2qnJSuT6F06/061lwqBCvJ2DTbnM/HbLU6gaBThQYN0Q5+NKJDt8N
hQM/C8XMpbJ/Yuaa9hXiVove0RPbfPXb0xeXQ+lW5iMaSDYK0v63qmLl2Tar2xTkAbuCp51kTq/w
HV1dOfKLUxwFEwxTXfVAucHiEmEPObZlt9oQcO/CapWBUKEhqCBMpUPhHXU/IAmGRwLKHzfTv7pu
+4WjmqFTFQ5iiGZSIZ3yIFpidEvKlwQgjxGPkrF0oK+h64D9sXjV2V7pEImZGQX7QPuhldbHT1BU
/bnYHtL0tT3NWJ1XT9g7zRgs10uV60vBfRMIKXjuD2BmG7/kYR1BHp6Wz4gTfM4l6cs7XoavC2Lf
uoiDx2R9G9/Wke6XUt5dmngo6RVZsPFeqzeuRqUj7aW7WUNuEJht45e9B5aMbTEwn6oDFckrxUqJ
7NXBQ+h5ugy6PnK1CKYACvI24IqknUK3nu5HHNk/+lU12kVA4K2Yr6ERygthpRSkX55TowHmLbdr
/PL5j7fi2bH/ApSuosSolM3SnnPltih3uNeh1MIzFJN+lONy3QNII1vw9iLVXWjv3mi2TNxnVTw2
JCErgsHUdd+RgYDmcOUymXFCNgMs+17JoUVhbYKhBgfFHwPQXPf0j5F83KsA/sA/fYteWXy8WNQE
rXi7TuE9NqQ3tlihc+Huy+Mr4pjhIn0iY+k6hsxw6kW9YnozFnWl5ta1TNQicqPxs81N4KhOgwhK
gXyKEuJ3keVVYL3+P/kzBEHkhS7g4/e/llCKI/ZcMdWdiV+glaS/3Qq7izyZXk6emNGYrllduVyT
ogIOjI1AgYOqKcvqgiGoT5ztWl/rWGFs4uTMB3wc/DZbrxJjbeiw6zLHwV8opiguuHNIaI4ru8mS
/RXffATljGtF6+hP4Py7zmO1CKJkGILeIdEjj/egUX3j5bjzWPwKbXUygVf+/zfEZN0Z2r01ONsN
3UurXgFpCxH0XKqPhIz8GxW01leI79JPlGdfBUYzRhrzzTjRMJoVtxzxpIfZitd+qMCBuc1X7kkN
eSDRS8AVdCYQ31bBiGban5rtEyTa08NPeX9fpOSFfn36bEdl6QAe3iWVTuxRCYHvi9VSbptoMKOW
Gy2Mj84OmYWF5uGf+99LRv4Ca4ZlnAcGHdGM9VmtwVnrdyOkg0udY0m7Tu8UzRGyx9tI8bKl4S5c
va2EdQv2DlZqVBKiGuu/PdbmxYPFKAXq/Jdb/ofksAj5kym+Xeb+EpPvierAekitPnXekbwXHZQN
JY0cpwtDJB6loIiiQ27AP5JkQZZzLA3Nu5hILfrpapZy50wCmok5VK+S0+o/E1X5sjpysxMGWHRP
0tT01oXX7o7stP+QGJ7vBDlHaixC/1YgeX1OPTcF/jR7yYf8BNA8MPuP90HsLLIvps9GV2e6p+Fr
EZ1XI8Ef80BKqhGY3+rSxcEAdS4MnHDPeb0hoFpXUyugTRwI0ZFnXeKUDr/vCFu2IiRg+Fjbmthn
Ud5WLQiY8xUuKe21tRXohpnX/jhIVIA2phheBDJxqceyp2cNYaPwIjuO9+TB2ztgkyjNZWduRnRI
sX4TMyUKNjX4h0+2YGxTRuLMhNqxFdT9ACvEeWWQQVa9Q1VaarOkaZJIq/T26strDW4zvdPjUq24
fkamJX+Uwmh8MQGjqRRcLTZnFUxYYY019MMPwi3MYF/VZpVZGHefIgm7ZeUZmu1LMbiy67ulrZGi
AsVFEYhgX1kY9uxiWsAd90GZh/0wZbnYTnERR+cqBTHLSHr+liDzR/10Efs5pDAAl3twJDNHh6uA
S3OXW3yKDw/pMPXuk1/V3VLEvfKr3wS1q65e3eUnyLsVVqEFNAo/+zoTzRNCZzE7wOiLFB4lreXl
VtprHMABxfuqXQIo3FrVQM13P2qiV4jv1GZ88G3VeNsoucwovd2U2GaGmtjSczyj8qKJ9b2rJNWq
K4NnaTSvmDfGPxXJMMESBd13y1ZD6RTVjHkS+yGq+DLpX4cbvVzDglnDqUTgQNP5QeQ9hPDKZdRQ
mwu2WMrxU8c5T5MU1u4plxrHkF3M6xu+wV22S5ij4kqyDSMUe8evCXCoGb8lF+JOgCATCy3LBgQp
PtC6syvgPbbNoJWYUWDZYuplJnEcLpTyJEIeq8w44gfHaKEP1ppEx/O6ZvhZ//VsgLlGi1bmtDfc
jNeunpqe50p8oxetR+5GD1GnOSrYMceII6plHDUZtsv6kRgQ03CKXcTj4rmk7THDufuB3MiLlbWP
/eY1mE616Yz3lN/Y6Hce9SZL4p5e0+f7wUQq0UmWWiwesbhIQoWC5GukcFrdrgD446Hqe//Yg1nV
5hcwnzGfyg+6kjtIYuFDtHJdCKJj7SPkqmF99PQBDjcOzAlMQUnJdpJj7Q6Dd94B1sK6dMXA6fgJ
Qc3B1xppN+mBLahX0Bwmabz+KloXVhSXM2rEeYxA8yG+DJzLwdBTgygDjvIeTGaXKVIdQeE7r5EI
7K9dtf+bl0jJlaPZqWXodNW7NXkKbj5dcq53Lh9S6teyMl+10+87uVS9twP68jUwbMJhIUwrwzsj
5G+WAlPX13x/vyeDD4JYEYkyDktNP+mbfdYBhSOK0cSorlI569yVinMwb35CzWrd+avJ7uUvAEKU
lcu+wYgz9+Q4CjJrdzCC4MDAp+RVaXqKvc64PRwZdPJ4DpV/MMslFKIbJ0FfUypdUJq4fXHvoDD9
jg3uTgwMyQ41RYA3fTTh/Ewu4Juwg/VmE5d4rf2GjPeurhV/X3FOdaOXIB9FPDHBjp/qkHtTjuor
hEbuG9bJc5qblvGZG7PeJRTO5Kcpetrb5G8MfMuL+SVYe0baJRmyKaMc7TZXuI6z+iPhRQAtbO/p
Fnui6d3MuKwXENvAT5/zlfv38lY5mBdMwc3M4drxytV0gZshXs4WOT0YoncVFS1oRLcO8MG84Mu/
YFX1nXibOcDVp82BAIyVdouNEDcObH6V20m3yA7om/s9PGJWlxrtL9xNH3b9dJdzV0gVnNtPNrrl
7wShfmnpwwErkcq0884wECTd8DX39jCIR5+zd1UNKGjFB0nIXNBCszYWZA4jCMryX5fnPVAxWAst
QDvhg41ZzfRuWxqcmhSemNJ/IKSP0uu/BIflVcKqzsRrZ8rAwd6c7A+GPE8R8eYDnr/J+cVhewoP
r55Io7jX37rkURVBsq6EwKqP0qXW+RwQ0kgCfiLdGkgoxMMM9JW9ds2cPsDuASzZAKZ/PYS3r8Pu
WaTpK2NFO9Au7uwd9YmcC5FDJwyN/ClQMaaGKzZNhbUbT9GvV10PwcaMVQBh2asoS4xtOXSFwLWQ
CM1kiBijhpw1NODLbj2ZXvdDtvZwytziwLXeaoIh1xhbLuvIxSr0WnMAtRgUWuA2hAV1iuGrwjfp
w2Tu4ZxHVthx2dQyCEkz4gvUjhWvSMHQaYOmnH0V08yrgfCuUaZpI0p1fAH4kikrUGI77VWs1eBP
J9eCr6jSG/skkS4pQ26nRGprWvJLmsgAOCTCxchJOMR0EG5N/I4uG0uKd4dYBm6tRCSUX00XlzwA
QcO6qblc14aTLQUl2LvIr8U6Zo5Wzlt/kXChmskcxpHuNmVpMcrI+7CTi2vA97pIk3xDXe+sf9LZ
bJEEljGAaJL9ujqy1fwxRv2PVPLqOWrGCwmQZqgKDz9PyMAkZkNITDjfD3UhrOMhZS+sYqGS1b1a
EWsDeo7eRR/hUThk75ArvkROm2pVCbEq7iXy5u/s90+rTSC/QlHojtouQ7T25JvXLQIXxki69yob
uB0mSOPYaWiB6Oo/rJu7wkAu0yTyvPskr37fdetRKUwHamcMdR3lkfKfG7gPXGaggz3zh47c1cB1
iaVbEf3qUWVzvGPCczUVORjZFLbGDJqBZbM2KAt2oP+4WM1Uky/NFJpxdVVeoDEPa5anx2RMrnZe
xwNNV2iPnMicbXcZ5kdc0sSuY/A08M9WwSA4O1UrwX3BjeOjD2LO9Zw/h+j9E5oFoGvUNGkKG9oy
TR1XzA1UFAzjFmkWfq/SmK35DtByneB1RFsMqX06mj2fWCs7hQIDw6TGp4XboKUQrkdhNYbGcahg
iA9eWPVxAL7qSnQ0+F6bMlKCPrqpjJnRdszs19JxKKSbDazeZBY7liyNJr6CD9+7uSkuXKVF3JC+
hPd36VbRWjrQaHG3cRU0FVa+df+KJGiB6gvjdKlOJvEzgGXGnD/19NyTpOsbQEnEEWiIYMNinjrp
J2ZJo5QVcfGRueYpM9ElQIxfmiUU90EUYXfgKnaZfFR4fNlZEFXisXCAvFYBLc1vynr3HABxS8Yg
tHmwjq0XbR0lyTsqRjdZTql9YHjQ3cUG4rYJuJfSNbSlEDarqE+GF2HhIlA+xMQbV6dxahs5RP5I
gcrNJGcRNgNcKyZjurtLGE8O65DTLpRm2oqu8SW9TjRVHJqmIeohmX5rQpf8cSCqErEj4dgcbOkC
ERcHzId5P63aM1v9gSe2fD6/dwO4c27OoxicuItCVeq/T6zjHhAIIM3tlWcRfHcoWjojqJuxce5/
BtRnNbE5yCHGQ7p6GCT0LeWbtogqNwOI5POwoImgu53PmGOHGe9Zqdq4I0xIOaBD1w2kZeHHiD/0
ldFpqh9mY3MPNZPfekFPeSwnLSeboh816PzdY68aDNPg+/c0EPC9fgwBnk38cCHVXGdk38lRPJG3
gVJdfGWIfIRz+YM+Che92qTr3ipth1uih/8chfh+cyQBLzaSoCYjbDLsbF/DN+ahvpLoBspWl2tt
hUeQ4JwP9wlt0JZ50ya24vvodN3U2UelM0EWi4hkc2qUqyyPaNJxGe8JTlbrlvVYUD0/JC15b8lQ
+Kt4VwOx2i7hlehfr4MNAd7W4FhjU4lTDsQJYssAgeaLDVl6dkvvmUwTuzwhwlP7xKgeRh+1wvYP
tnOqbCk+ZmUjOFz6e02ymbMisDpCVrTok9VkvvN/+8HwDbS4erhoohPCIztF0rARxAlN6cLp3M7W
LmPst71GUHSikg8pqergwjDIw0a0ZtEfyeZhpaWyNhe9rJ2N7iajCUqB8/g43xGcTDj8coNnyb1H
wiIZF9u6eVaTLu8GrNW6G7R9wppD5nO/ZW9S2dY5vCd1SnmSJbjkJP2Tv1xPS2CtjkcaXe+7d3In
/9ah4kzzErLlCRppgOqxSBBylASiWT0pNgqTwFU85TDYSlvQOrNsLWxbVCRsaCpU9T7Xhvx64qMg
YZ0KoVXH5+2YoTiM1Gcz8+e95gFCUE+y0PCCyfNJTUC8geX1V2UzzG7y3nA3alzAptzvz8KeFrLv
74uA0m+79f0yNgHhrdUc1ME9IrLGQyYS3NYAL9uWRkrxRnF5ELYVifbtVZtEK16DBpWJGq8fPOhL
J//9bbWUkSo55GF/UdAhHOhGamCsuOQEWLYE5uUIGfdnKOt4NkZdoA4sNfVAe5rZBdlZ3OnL7yKl
Bnj+6qfiJSdUQCl/wI8cnUiqD59BYpU1T3Mdg2+NZMjl1u17m+g4GEdeII4Uu1+ZtOmZLRyEBWI9
Ire1S+Ls5UCsPJasLAry5uzWGL3QV7M8VXTP2Gmyv0FlmH0lwflGCR8aRYhZHbBlmnI6L7x5RWQc
XXCPdHtUByQS0lnN1tcAhIl8BCIjFbaD6hwVFd7d4GNqMjlp9Log3lE4/qtmIO3kOiEXXgcWTII3
tyPQK9rcIa2BH9a2W0KwtUIAd3SYxyDY+mVrVvjGK/JgOJcH7JAxAex0t/qdBZRHRgtsjjBvLbdX
vis/cI8RYmd9H/2CLoPywcewB3Axp6Cw3exN68wPyhnTufXTsDU36cI9YfbJZPVZ0tnvqcxPJgB6
KV8qdL885kEHLH4wN6/e7kCgHET1mcupAclxLrOPHDxZu7xvmdXNO3k4XCNFJ/6B5e8lrKKmRnnD
TY5Wmg4wSvCDuyjwxt8OBA5AOWPs0pIe4hPT6dQaRcvfnTTf8jYQx5JVMJSW6l1Di1gvE01GgqNK
sLDbod/DFDDyEwsWJuZK6Aq3uNVIAt7aqNTFE42pa+hOscUNGucpcoMsdiUIrbqdBSD3MLmc/Kcs
HvlWHaut8bt92y+jn0TvGcI+EC18qZvp0l866MruAlTM8MnR+MlOuncOIEcaMcusoe1pKfG/2+rr
EWLQD4sRqxd6c0+59GjuJ09pM5RKMYoPkYaPzxtKyhjFC3EjhYuTldXiGIWUIxNttA/2xd6KSFDT
atoyCON8I0OH9uwMkzZzuw0Cb/AYJI3Fka7oZ0B02ln6A+x9co+TI/abW4gGmmk9jA22B2WG8xLy
4F+Pu3mdDWgPtXAwy04oJFwyEriz4QigKYyUZFq6rZ2M16QcwDR0FIBb+F6AG15w8phtJe1wNy4Z
Hl6KZdIrgkOdaXcL3AHKGMMf24Bay9O1mq6gTJPp0by7fbmPV5ZjS/tazg+W3cuZsLpewkDJ/WC/
5kq8bNkC85CEVaPP7QdZ/attmFZ/BCwrn3M+qJFgX+gB3e0REWhr96Zxp8VoxIq/stUyxsFkhCLL
UlgD4mHy/iPmIqtm2LTziJTJ8nf2iRp+6oC3Puw6ii2GYpXzPBx1n0sDpl9JOegH6j/reu3HwB/V
lV5uFdJE8jVb3FWDP587nmAF/Z0JPJ4gP87jLM1pqjf58DRhxYWRZ95zS3U8Nx9L6Ods6o29HC8t
wZ3EnsjAWtfsXBgTC5fG+0Z3v2FLRGtOOXwtIo5gMatX3cV5QGgOhRXpRp372KuEA1+7CUxZ7zIz
AHyv/fzhMw33vS56ZUDtAehlcu4865sGRNEjpUcHbr7P11FA4PbVj3OQAfeZ7upWHoGgxFJE2iny
NNqqw8fuRovyeXN/9kiszBlM4bl5KiWm+2EHJh1jwkmNDW2jQp+gFR6G/oRKpsf5XYHoeanaK1/w
/lOQkNMQyCgTxtANZxFJIPrfjn7i8o3Hx9xbMiPtJz0lDyRbW16t9G0O6ri4PMRjhkdKXEDIy0vL
H+MkEFCqi7kigIAaxV6I/wPPK69c9E2LR5m7OJ5yUu0OJQ1bw67V1HObiNe6fB8cuhMFH7AtiB1a
gAhjFmOTmLOa+SCitahI/HYHOMWGRVk62RlCzc8UT5zeb3s6RIpN1upx9QQ4npwYSXKkhAzEKLoD
g7klyyOlWCm7MHvMnng8L2NI/uCGYwoExJgUdR5oJhUX2E6P1Ub7Droup0qLB/g8a2HI0+Hjaxbm
xA7OdFcW9MDBoVI1YnIM+75QUEpoOjI+jWauWjf7hnRdvE1Qz/xnRVfgYsX4WEkAkKeAiV08hOVM
aUZvXGFRQcURhPohr2l3hRX4Ln1sCaDXwi4ucB7h5OEsFtxnfIn8ndIGophDhWGBBI3TuKgi3ox8
AqVfcQjGuGPNt4Vg/kmoHtS1I2Sqm9ekPbmgGFDoAbZoQ1VRmbY3yELvXzwtH9hLJ6Bffc2kEO9f
oze2CKKVxrCa1g3naBsJE6X5ButfKQDkkUvEaEYyDPVAinPu1WxVHr2bGMoDh4G8kl48OQMkNZx1
d2HGxXh4EjU8d02RejfNV6+I812oASwz6FnLKnz9oQONDDqOVsh9kb70Ue/JqHJ9p3l7ifFo2TWZ
bqFeJaxvPDfpTj4IEFiUd8cR2DDvF2bpvWWbItxhA+wUYu4w2GeN6VslngKSdfsEHrxuetA7i/la
CJqn/QDQjsfcTVukoslgjgEDMfDAJNNgwnlO++Y/0ek1OGue5rmx3a40R25Jwi7VcSwOfh9Sx8wV
nLSAx/ozRxLWgrv64KA5zb9uVyc4HHCZgWam7PAG5b+NSU9M8qhPXfWlvV5niK3riOpdSBSBQsED
CFKyLy1yBxoICcCe8l5THxAwzTCqe9v6EjApaBh/rapA9GfISlILi9n5U9jcj8DleW+cNRZI1Ma5
mSPoVVzDkkXYbg98Gvn7e42OTFtTvoJ355Gxdb+gYFcwR88rUWLCuJTerzyCjixYGhz7aN+M+VYL
SSV/QHZwiXmOVv6XwJL0SaaNN8PsqCoxUQiq31fo1MugcrEhFQCgmvUc1hEE5O2EM/ZJGaLipJOS
Qji9TIww1K/ccKLrX95nKlrqbQAL06H7cJqJsFCQ0dxpWA5KW2LoW09+SqgmmKJ9akG/jJtwUVR2
ndF0eBj5F5BzB9aeIw5w/w3WBHGEbHCvvtGtk42c/OMEeHWfoaq3DfX4/oFxi2Gm5d3j8eEWHShl
r6M17iQilpidZsFLYp2NwUEB+eooYzFCcSxtJR7PSKkBmMzz0387Zbj4qzz3tpN1rsEspY0oXUp4
8C+FHEG7q4Hg9S3UkMtFZn9jBIQAL7Wpa94J/ZYEIGfIYX/bEg13wfDLzxjyYOc7AlGtKJrlkkPx
5x2QTdneKx3eulldC5Iz6WwiUGXicQjCNIerfkXjPKbvsc5zPmB2Rq0L4EZ5RMVfkROsKX59XS1V
u1e+QYQ0H6SdTAx0uid6l6UqPdP8rNS7ynh7nyBuAI491j1WP/3koEgml+HivXerIFfnaWCZX+AX
k9qTYXhwLVlu4ZMySHRT9FQi+zvARssfeM7WmxFedjIG4q8Szt3XoaqMN0THy77qLgwgXwivAkyX
2RYphh6ANQJweL806AUIB9G6cOtm92PDOjxNQX8RrAY2fFEAC9urYEDCom5N7+/IAooY76FzW7gi
+IYKcbYeWBzy33BZMh+raUutVxuPih03bkqLTCin2n7c35cLwqYUstLO/tBFbVhjblO85UWJXUSC
bn43zJMrJfaHyzjwN3VPA8KV/jzWcETijPdsFjkgkEt2njyoTE/qboHcnkXE8Ndu33UI05JnlSAh
YQUCHHy2PbBb+HPOK3zgqzYnt8sogjlA+fKhcAZrb2DSLRDRqBK6j21VqZwgTICA0VYTQX8nXJIK
lpmFR/2IcxKaGVnRbGRA1uOZW8XTvhGVpM+q+SI2Do9pPjsfGZ3/COJS1x+sr6XOefxxKlx/jZmd
WxXbqnYlIwRSO0kBWSg4pwGiUVAWMPU07TV5FBuwPQMOj9hUH7H3NqxF1Gy7pxniJInUdyjZEJb0
1qHdP6lOe8l2xF57N8Xozm8LMbEU/CeIbs4ycPTJu955VFGH9gbKXlPLCN3f9MzDsZ8AtQchcD8F
sSxfENbhOA9N6bG9LbfovAHH4fPkoVnb5UgeFCCm9oBydfHM5W+GVy0thkNlmaGTSPA4IEjtRfHy
DuaIck4iBMmVoAfiyIyJ07mnWfxLi6OBolWoMZ7udwSFtnhGQaIwGo7qjaBe0suUYn2z6gUEzMS8
C6JBuRIjYmkxYj9bC21f/A9Fen3YZ0XgZaoTX/SFrYvCxOrKhp5r42W1Wmsnlr50Sl/7BqtslCaz
te84Hl6PjU/NiJmYnNjyp6x7tFUyOmS05LPbg5UFRyNGLtuNXzQmLOk0oa0vJLLyBfU6p34I1CdP
25AGb+eslNO3zYNYq61N0bcx6Khl+883e/qiCaOC+HWJiSniDNToj6eh0YKIzFuuB5eRk3PLVtck
t8ahmczLLcsuO53hREryQS5v4cKA+a9drZeWvHyP+TjJjx3PTA6nkpr5DDz9r29OwlDicD8GZVaL
LJz3xNCOrID4P54glB9k3/mZRobkhcCtpM6pPGOhvMjFK7C/5e0YrOknei4bxUG3xScCnEgaLmzB
LVqRlz8LC2DacxuhAXEuU5fbS6zhtM23oOelqiBY8UQL8jpBCGIJ+myX+HhQ6gZ6RbgzlY/ZzKcw
mY3uoGvF5+r5cYpzNyjVy93Yi0gohBuS708ePFl5WeD7HxZGXAj82N9dlzV3Z0JN205qway6YdjB
0UPJmX2cK1tcyhayvAvl9clzUIzowhZaY6hNaGINiu1V1SAvdmRfobieB5MRKP8vBGKzz60fGY3V
5Ukw8oSigffRW3n+PrEreWsLGEfgJqPrqIRX9KsdvX1kTNzEJ2YgMU3Qn22HNLAtuTRksNysqvkg
4aPpNDfvHDZRFsncZQWyDlnOxNZMo+u1pKE7DughB/VB+PGZdZhLA7J6tO8qpxpHIJAn+HxobOIm
xjpbBvyF+pikxX+gyOhl64MN4xwvoIS+m21paUHKBQztzKpaKwohYm0yk96kypB+TOCWgTaF1in2
e9SdWxVeRyULZOEDnXWmTDqX2u1dh5NRxROAuE670kw+o5m5EUXcGiO76pgAM0aMn0d+lqp9bnvM
CFnmhdFqRkklnoQfn5OuTOpUvHaQjchcDwfPYmlmvrslr/xHrH9qqDJs53Ti6qhs9h1U7IYu1G40
osaU+5pK7t+UqmYQ8MtD5H9FoLLctCd3tSXF9caIMbLctGIHiWRdvvkl4hrNRZzENoWNuqEXdC+f
Nw/BWn+I2MUTWwtFoL2elmkr9wEYVlUZPvHv9t1ANN5txs5jg7TArGEWefKMaC/cL5gZIFBc8auQ
Z0t3XWufVEDQb5tCskW7UXWHtqjmQTlnRSEcR75zNAZkFl87Udd+0AEjLV0E3m2I6kpH/W/UvoE1
3S7Jd0sNuWbLgHtu/YrYXtXu+AluKkuvgvvUZkONGI1MG2fjytIQzMAFC85vHYx4QyxU0Ef5+3Ky
J3cZbVPz/qlC6I5s3bv4kCVMfJTY1uCYsvO28wfK+4FV1LxVsrI6uDgqxttPceUhiNcqCiTb8vYb
hSzFyNi24dfER3oo+Q5OpNkclk0z30why7dihJJJD3hEj8tunrhQQ8Bzug2la6+zrRc5xJJzjJWw
AUoyKV/uiqrb/VxWMkx/0mXnjLh8MZRe/J0tuc0PP6W8NCT/oWeMWywNwVDKyRZZL92KyNB+5XQl
wgD9OD2oX+PWWglKCeOxha6v+ke4BT94nC3MlyEctBCilrwxecAK2TWOoDe2n4nW9zZVR+e8fMZA
lgYYdgGbA+3vbMl7d1hGDqhX3R+ZtRPmRscMoCXSG1F5GoPvgbcHa7rSXLsAkTAEZdLcYhC16ZB8
EG2Ep4J94KbEjZmP+otdmRdzg9gfIgpyXCFDSn3mbyUcFbigmA2eBXQe0/c6isixHf88hRPFCur4
JYlVq5Rsl1SMXxWtWthTtGeLbnDKmvFEhWWH+FfqawvB52lI6YGEiF2+SHJ/Q90n95zIWaHP+suW
ZwOqDRlQY0j8tVK2lnee/C3BrrFA3CNdqou5GxXsJlHMHfgH2dzRo0YjFUwme/VdwyiSsxq12Ej7
wAcvuJga3H6ZYBrGokMGVxihx3jcV8e0oDnV2uRV8e65traznwDEEpiNRcil6kIVeM3lx5iVfW9F
xBDQCzN0XzIx08fvghpv5Fdhum+DR8ZVBADF42uQoEbeY1H2i39LQsAGAZ3BhXLP1fOy6yUmJdcG
qZwtzWtRYuZALzo/+tOL3mUsOo9BgUL/FgHtYSFZwInACc+n1DJ6COkGg/MRiImK0E5CWsD4fgYg
nAqQOxp3z2ke3q0slx7JzZ5BilREYyoGN1cBii7y6SCuLL2fY3L4e8F+L8eOeY1OJoVhAizKhiAe
DqCSuaFzAcpUUcPLvQ6bopmruwRCy4f1IC4STcD0LJLL8F37UbJwU79enQkGinuCank/kDTwyziW
i6sk0d2cejwAnTlApMX0nSi9aN3aBtuvMU9lfw7doXTRWXJetU3vvPAnYd56OF3aE6IL4VUmS0+g
Vl5+z55gxb2QlBj6XmpPOYaZyYjNUgaK/zN6D6Ig7TZMnRB3kIfMQG/eard1OoE1vKfVBu4IxYhn
SwUHyUXzL4SB5aSGCUH4NcttR2pPZcCMMhNQUOr963u9QfALNJZBbHWHCpHayncW76CFIFBm7y8T
XNJryPNZq23zmTQZOoEMSjLaq6vjFxYw+th00aJf400s3MptuU5JS88JJX5tPpw8B8T9jBd52vC6
v0JDJwom25wSZnS2ZK7qsfHP59LKdPCO1/m9SSaq5o1+5qDzjUPsBJJdJJxkOPNGuT4B2TVnPgNe
5mdwlTp54gnQthJK/eNIsoh1oe0cY7cCA4Aoayp4dLo8i0GIBmYH1Vt+v/S3X7chdtOLEYVwzxjE
4jD26reRDUXHQ6gk1L+JJIemqIH2oKAH0s2CH4dj0RpzqJPWsU4jFy1RXKWPDs22RKodTSxS0L1+
IYokTbn4Dfhan9clOpfpw/WmWVmgkvawp9CssdCg4fGnqzt86unGuiw0uBpFr/STzMnLc9cnBEjj
3wl7Q/TzcUmEVX9fJxKTMbOjFhJSyicBIsdku3lv9/KaDS4Y5TIQw984qjHASfwC2CejiH37sJrg
YzJBaNsR5BbSf2oOHv7OzObBE/RB/29hUyNOFEVV6ZRittqSlxUYfvB643HwAGwvj7/QlFeeKAk7
GSoIAm/eBJO3K9MNF91tFVRoIwYI9KhaDN7njv1twFviO+g5uFH10L7FI+N7IJIsy5xuIgdfURYu
QirwDt3FoAEL3BX9tg1h0vFc6j2M4wJNmcdIQDrK7AIwjvsZvv5QtufBQzf9vfnMUOx+BjrDYdS8
n4/oExwS/0mnAd47BDf16lU/lJMBsr5VeQRouFZkgxoTz1dW56GMqNMgpL5Frtvkr0TUxKRjRFzB
HlhB77QEzGxRsgbcbXlupnfHvMz5E+uj30oIExhZ77S1UkSg4UlGY2axLUD8Zr0es6iC3G/4is5f
xmxzCRUz0bmImrXRTlgNnxSf6LBZTqB05O3BrVFV4n+DU01FsgoqMWaXwZkdV5T15jyp5G+5Cfm0
iOzqjMBfogGdOmmMEI6uNNkINebeY+UrIeVyqDXmlA9aIboC8Al/5HrGfMymAJzDkNeBZwLMwLVR
3N/Zuw/Rw4gxCzAQ3o8/BExH3yCcQRgZjuTQ9Fo471CiPZbrhAZV6dGlesfPelcggMwjg5FycOVf
7kXl6nNIM1h7AxmdQyU9JwpHykLEkSb4Y7u2Aq38ct/pCS7evw++7KEWPuJlk8MtSays99imOwzV
NRXrNNHscaCwHEzZ4OXtH5LYIO82lSV2JhhdiQKBqNkdAKK0Pm5DtyaZAw5SXDQ73iTByHBPwLvW
IfnIyDeokWvYP3I9Cuu/APnYhPM1Ktcrkwisid1SgkRGHT26jWqMEh72qh3jqmtfQLkLoGKTWyTg
L/iTZ5atGQPP/eGTL6bFPg6an5woO/wZdbbxUpBRMj1qgGgfHPidCNVVEcsaMZkPVDF4Hm4RrjXE
z54Zcp/zCP/z73G0W19orC87Wd+05EWeOXTk3vk7faL0UOE0ett/axPJDQxUSdV0bwgpE/UOCQwt
Hi5FUntyL0/hWmtga69eECLpicGi6OTB2hrjzNJ+lB2Nxl42+0uRNQb/Jqh97APaH2pGBmVV0V6c
MgmY+cIxrH/yqHh5kipy567y2gJ7zvwAB+Bqw+5QDk3PFUC7GMqR2PB1oriu1iizTY3/MDUJQJTe
1hgqwaBjFbJZl8r/YURB6ivoJPY3wGHbNKqkmvIfAeM/TRiuQHTthR8FNCZIj4CQkNFII/6Cs0/L
DKRmKt399iklITv1L1jcmfHDpPWbWEcZHWoC4AXInOHrpCPmWW6wQC4h46CVbVDyQ0mIuoIogsu7
NUGYL3c7HKupUEILd8JHnq3f97XgxMZfZWAy4ZtZybNvxMobFG9b7Cm3xNMqwv7wNeCniODmuYbC
1lxmWXhc6mdhu/1E4noi4Z1nWONgCDz1yTzcRyDcwbm/XSGUvrOv5gpXIWY/uCl2NSuN9x79cqCT
+cQv/jXHZBeOLb59daXwVX2XQfWBnlXnFDpg0MHg6MVykwT3GomdHG1Kl5j6B1zPsemuf3MufBHV
O2Abfm5WtDPDh8yCG2F83tTzYeM/8fGoJYeQ6lX1dVcWvBQiXkofDJda8avFDLLLRAgzAWHwLwZc
8Tz7CLxtVq7AJujrnl4VwuMUVFCB+/szkvx+LGL6vuLmaI1rILim0DRfhFRWVhqB8Rev/Kl86zxk
sIovewl9CcTgcJWpImrghza3rM1iwdbzxq4TlME6rAM2yKWXW1jvwWxgZ6IPh6yF9SN3RlPgNfW1
u2KloRX6B84q81Ke0OVD6huE11ocuU1wbI//dM2JArKUPS1h06DbKI0flvyvu9myz7clTeScyIAb
yCXrYnmp8dQqRO5IYJ13Q45REzN5YMwbgvPZoXNQqyeQuxOOqWEm5ifoYujRgKOaCIY6IDFUwGD+
Pan9a2/cHcLRNa3kC7uWPllshs0Cy8QFi3Bch4RG3CJve6QovaolxxqZ69pRsupXfvlRV/YNf7km
spEwDLrN9ZQWdvCqsFQJjOT7QSB9bDgn7ULrOq9c21eAn6uB9PJHPqb+qczHW3c3lc8uH9LfRUrn
fntnGYRPk4aN74d05ZWH6qOcQ4FhpFRqScWJn05smOaDNT2dRafwfQLDRdlVe2wqBBhnuQlRAnVs
za5y+4Omox90D4Jnj+n2lvhte07ZuPkOLGJZBD61MFdPJbawy8lPZgwcGDDm2HSbDHH5BnVjXKk6
C0TtRPFakeS+9TG1GLSFP8SVOnAHyyTQSvlOd6UEJWxdzXk/avlhb8J7teNpvgj53x30rUX5bLc2
NPHpNzQye/H96EB0I0Dv5A+m0dgYhTjK+RzF1diubV0nBwyWX4ov+waVdrvKTvD9XD2CAWWK6944
1O2n5vnYbMGjYiX2aQUu1XfbWfrJ+vJyOmgn4fYaP8OgfdaVfzgQZAPaiFSHN5Fi2ojg59bI0SPB
L+R4ClbDfZ3Crb9wvw2k1uJMwYa/jbtG1IyFN0iptDDjZKaVDVb5mn+E4OLkKCBsGyEgpSqeOVxs
/P/I98/JC6wIUIDLB3mcR2EabVkJWJNHEkvWJsJdcoIstR8l/Q5cX1ugF5a4GGVm90p9bC1cpX/T
Q9dNK39ALKJS/bb660dR8/NLoc6VVKirHr9S1Z1C7M7hdGVq2FvDLnmA0MvHFKpkMnOHdmIxiwVm
/EriYfo4P5iSKn/7Z9HZeOE+LSAGqnNYbfp8pK1DVn8XWnbOAjmR7NojE3pTyUGHLraXXYT88yGK
O7IW4edninaxhncnJD/2vnjvktmNiA8Q4JFWRS4ayq5dfH7+79yOzDO1tPZiQFpg1Dea844y9G08
laoKbB6otYcqc/TOSeepLi4gWXyahxi3sZi0KW0HftiOhNyQhKg8c0xG9ifE8fpqOabLhPFyxMcX
sUjZNgI8ybwF5yPVSwF3J+FLO7jAIfxkZNEHdb53CggWNkl0vdp8nv8jUSr1Q0M6OVjsBpHM7Pwd
WKRENals77DX1IdtyoQDICeO8uBlS2KScVyPBY66pw2E/W5eST4R8wSe3J8ZtsfxuMgicIZehioH
AwViHfGYRP59ZaSUIz/TUwtoWWBg875bjiCWzo1EmQjPW4EYaM3osdDiClVKLQZM6b2R9VvLo5cE
paYB0+7sf4CxK7r+QmzYVLU/NmxZguPwF5phKwOjVtBnINAzf9pbyuPJmWOesJRqZ6gEkucO7xiD
52hNkxRe/V1P2OqRp+khElPhQDSromraTBdledEVMiZ7Poc4uCCERP6hxA6kjJ2SABdtZih8U721
kMxRF0yWTGlodIa3ffcu4mBZbgDF/gKkwo/IHlDv+cV9AVNuAJtEtadwkl9YVSFYczpArRyG29Ll
VDXjhAqKUFWQ9P1oKs99876wj8+AwFK4Ju2Eg+XeLfRubTNA9iYHOc10IUSfLWNKk2o7N8ecdTj4
kNuU00idvVzAKN/HnfgcglL1zVkYjGG3sVhiU0LpVO/hEGyocsl52XeQSmkXEz96TvUVc+BB7dbz
+up8fwgrTuyz1Mo4LcY6I5KrZDx9nRDZE2ONbBdYtxjSiy8L8SV2VtvEIKTz4G4WLPnaDFFXGsdx
mNXgjEtFBAkmKWYtfqz3qTKcgUh08HMAdbU71yEumnrhNIjHQRlLaDMrhbplt8pQbX7MHiwiBDGc
GefjyvYoXoFluJHtb/CAISWiIzdZlZorg+NKJjjgzu3+b5D9atz+Xbcmx6FhnIlVCiHvlg8vOWzZ
3yGmmcG02J1A+XA6eym1L63/jvXqYvZuu+YEjj1axXgBquae2nK8P19+xQEHnmrwxOOycacfXbZQ
F/g3BMU0o3bBNYzY+0DcpvoSJaChfp66KJrbpR3dHZ2ORMBKnval89Vx+zg4gHOLOAzJp8qE7fQA
cAQg6Y/PPnqTOm6mTfrM6T6T1cYmt4AqQcb4QQc+vq2cpB2a5ht3ErRV6FFzuTJqE/pHi0xJlIbQ
C8QmL+/+zGOKma6Mb3x0zqsN2RqpRbT4yrTR7BUK3MgPSCqfPQI/wz3I1+rKEgiHlVcABHT4Y0l0
eIKa84nA3YtinUb/fK2p7oiqgzeQkWD8NjyXRmoG9y5clyW5blxavlCZw/jdQBMDtjDcENOSiIw6
VEh7HMX7BFT4mwc+RAlcRZhH16wFuB+guipUYwLK7UpZ/JmuUG5KeeWHkA1dPjKvv3Fp+A3xhADl
daWBsNCO+uylmp+LnH3BCPyNkEY7rW6obYB6oht60CL8ggrtcN3MBba1oGSXr2cp/2e57T6QMDJ5
vJw8XzP88AuU5qbV7xN3F5xbaVBnclgVQ4ZBt0HpgPRtofHTNKE8o+RKXvMxYHiF6qmu89rWkZ/M
pXav8iK2QSHm95ToDW31ok/WCu19lGZqAlnc+OjoFXQyzB5Z1z/qjw660eL7GfKH51lUBBSBpIOT
S41GHO116Wju1LTqdubhMz7VXJgjbYh1WuE2gM156pd4+P2z53UYgAGBvwAMYPWufORxRFZnpomg
2As+CxphuK1zkJUxd0owY1kSnbB1vQpepbU9I52Gvi0SJmOmZ7oTf4EefSEoXZTfL+7/8Pty2xyU
D81/WaNfokHwZ5b3XKKFddSvg7ivrVapBeaUtOqcniQo3FES44Xff82YQxch6i0VBE1lBEgH5I/g
2JsRRjt8A0qMhK4WwrELgWRh2X69G+dX68aFfpDU8OzC6621jvB1bchfV934i0goF2qyUes6rlxo
WbqK7mukcVi/HOuVnGTnNRiVBwoI2UrN6+Ef/7knBeQ1ERkzr+SaMlv+FsCE8CvlNiB030rp3BOR
M/G94LBr8iovzTPr/cq+IxI50gLddXjLIobxcOoTmsFu4zs0uYQGufPLzWoGv/tNIOGs9rWJ02fX
5c21mfhtVFT9LmSz36qbbzVoZhckveYDSlzJoEw36KDCmD0OKayz88mzfflcxSmmp08yi+N/kN5b
IBXsaI4EdQvIATI16ZwAJnkXo7gJYGTgo0iX3BSVHBt/M143fJfCQwOofezHI0fJUkSz9RY5+TwA
i9ExQVhM6EMf7owy3DxhASTSGY17UatLpvW7BVjLrEcGAs616MjY+ZqZRBENrL4m0Z4Iz2+Mq5CC
3GyTa0pELhU1HyVJ8max6GZO5k6Y1gCtcn057cksIEfpI5py7SuOIOmL+MTOe1hESkDBY/VHqI7q
cvuJQzCU3NNmrhAIroteQGLoFvAYQIM4ngpLz1RJFtlprEPUPS+wPCaloQ7UYSq9JCZPKR4uQONW
6te8MDc5hjYrjbjsRmgDCC9uot3vWyc8PkGFI8Xt/zaayah9QVX17uJtRVrqC6BqlIiBH4vBscGL
lmYGVCg4TpfLtUsMzQPKIEhC+2MBlyP+sY4v4PUe+dm8rnwgD1Yl1O55HVqSPGQWNMyyYEjS+UK5
GDq9sKOK4OC+SQfsHt48HJCImaB5tdzOOfL+IZAKpbaIF+jXhb2EfFe4r/LCC/GHu2Zx/zte4bVh
/o87PHlnj9UWOqJijyuFrsMw70Ld3wvGEMWa2XXTTeE/Lse6EiwTXh5V8WnXwYMY7gUjB8V+HhKb
rR1EunKTM+pO5jMjnrCn3x0ZzmGNuThIv4FDXGn7uxVubYUXqQdZ+KwXeE6a9CP2Z9rKVZV+3hmc
I8bxUEQfOZGx2ny5sfu3wO82eg2VFwSXfU9mhvh0MBdrGBCgnniNODEKmFDWYqgW/L/2t4qE1yq4
/PO+ipD62+Xn+bnZYukeyC3ppgXrl8/rZWsPPm5yD5kFWaSpk/fTcR0pHym7tLBZUrxIkjVL/8X8
cjJmOozsetVb+96UHJjp93W0CKVITcEpvceuVpYA6FhUhJvIi9dURpevHCbsXQCPuPa08NUwWbGw
7rCnYpalhv+SoPyo1QXjhg9mRX9Loy2srYQHUzUW6AJj/RBQ1ifetYUpwriGl8ZNpfOU1A1PsZfe
+37KQdaGQgrPNusaw+EQUJXF0Jq4VuURqv98ijLIwVVgW32PkZOTIkGbbBvG/YVyTlc3wt0XM1Eu
YzbBA+pAK/f/L6nncAYRwXR0IIn/uMDxN0SYXSIRzacXyrpaJJwxSH8YK7oMRVPTPequsTXxscYO
k95C/USNNZjErisY9MOlTmqOVtg3ePQ00gT9VJTKAQIQ0cs54qQwSmSex3sO0c31gtIQzWZAv5O+
g/3eVtZEdfpwNAoBktFqiqRlwjQfzJC2jdpZw+5+HyKVTelxW/5SXYEW7bHGQV7oAlTkh9v0/Qtj
DLLXJdRXNvOY9lGea3HIQz6y7IDxLGrP8eWx0/v0DOQJKpApVNgKvRHMXZHq0YPDxuoJzHRKNlKZ
v0qzxdNj4rtPjKmeDlHmMFsrGfoR7hwa19n2qdstbi21MyzirJxaGhc3BMr54k6sLgfBUzY9rOeu
Ff7P4vE1B0jvHO3ImDjkNhf08fdHcDLpAhCulqETDvSu2cieeVyNVyjt99/VVeyzwqQE+dnDwAfD
QXZb6+fOkozP8g6CQZJUIfdHd2idDkqAg6cqyCDzuMOJPX30CHNiQSLIoxU2RUS3s7eDst4A6MU+
kozzP8uT5UPVOYMKUUBkWraSx6DcEaGsqUfxCloIyues8CFsP9SUK8FZoFl/P27fmJOf7VL1i2As
qE8TG0CqZd8mZxF/CIgjtbzm9SpwRjDgRXfNXJz/b16esYaMKupFLtFLf4tq6ek/0vgolcWmDZCd
z9f5uXw6wXgk6S8J9MmY4CsHesoDphtq1nl/xNB+cRiCiW/aJZ6/DtRcAd/3Jq17AL9VJXB/6adv
Bi1BzjANX5LrKt4xJZicPBP2O1PZLpBDOIGLRbY6Cd4f7KkoSJnRiRtlIetgJ1LZFO1Y+89qxf7Z
aRnomGsW3rnycyOHcdEg/DCtxdL6y1dJIqKN3yKk7PL4N3CmnUhowodCSivnvdicyvJr3lWKll/e
yX4fDBQQDkZJ9b1GAMTA1kImWi3jH4IgX9jUE8sJ2ftamPfqOzryCL03uZ7YBCG5L7A+zk3oCj0N
p2YwVSe78Az6Asm4mSBlIxRBh5f+2Pm1U3WfV70T3cCb7UFQ5QWRZQ+krSXp2LSE3F9glvXWfUDB
0lnZIR58HAxIJ4YX9UJqyQ0ok+xqoQykPckUt4aXy4FCDZ57YU6vpOanDMfTh2jLbMMgBgm5h/1l
riH2KnNGOcHlanvng3kKxhilxG928iFGgv9WrKyDEiOfnt1WFlJiNNdPDSjXJQIYT5S/VvcLjfrb
i/KYEWnXS54nWoXSpQ+fRvHe/FEQ1QekN3orxErgo4Vz0U8LD1rnawTRNyEbUjL2wBTf/KC8KaEQ
pt34FoPNQrRqqH5CVemWwVUfairgIpW4tPQbXGaHemR+L/RQOG02/X3Hxp6ALZ9YMAYKYxkf4KzZ
uqgAM2bWhfpknRs0CyVZ+wdSDp3WeW6ubSloQI46Tma05yHwYYTHRBHsRQ6O+HjTWcvaIT4g82Qf
BTE1cCB5bucM6HwIoimi/WqXOsIW86c5tNJIMmQRZAwsrM9vCbKgnl2jjOe/DePpYrMDsDRQ0Nwd
M7f4UVXeeKr/rApKqXIh6HMbV5YgFQuxwxvG/oWMg3vJFeiABS/QG9a9cuoVInA8OmW4hPBW7VHc
Ccz8I5H/vPk83JlbmnFa2XP3wMp4u5mMigDVzHraIt269azuuP2OdObangMSs6RVLkTCVjypr0F1
hUp1VKfxDnlLp4bV/hglCOuSQQyZAp/B7n52J6vNwq59rznRSfINRol6aGcKYjXJlsbgZZxz7cb5
JAZ+tZOKnH91m4XrT97NhuigKER0m408gfQrV4AuTSQNfaAMXBBvr8x04FTqQDDb2BbKKoqMssd8
PTc2+MmFFa2RPahuDmwKZ669LO0qXHuo5SZt5UlA/lHtBcr6EpPD/BpyrxKdSCMcMsby++7OFjWP
0RuKjUNdUfpVwRsOduotUBV6PpGXiMqbrYsxbNce6bCDMWzAsQnwHkPih3kEL5pB8tNtGjEgGh5K
aOZbspOpRAgmua9IpTR6nOrInPhrHH4n54+yBZD2f9u8TJQLaNO+Y3nrf1ST/JdQ2xTciXS+wKSk
n9JbMR6Nyhu9/bdRDtOXgKeVxrnAkBZiSCPvcIySQG0FZN6ivqv8cxEYqfciGZky3bmu5CdIv69+
//8WRDIS8YQMkd0iWLcw8hx0V9CCrPWaJLJy3M/myAoeVEIZs+dcdieZCwnZOsnRAjNkojypd+gG
WGQpk60znfJ3Xf/x93ESotmklUj4sKMBfMQ0oE/AGIlWU++uCjEk2K6sWMpHFxx7Q4Ob6PvPBFZf
mStnx9JMp2mYFVtj2xVUwq3ll3uBaT6ysAP1ZbpH9C2fW1kPz9Bwjj5La1Y71xZYmubRm8U58bTX
zpV0AGuDYPd525myjNJq1RA75maRxX6tI++KZ7GHv/mJ+izOlDJaeAa6yZai43nw0kl4LBD1B2z7
//cl4AzxOfUm2q18dklVRk/sDuvoP4zfvvBxEcjOEaPUlGNUwqKWWaABcDhB97/obz1ROJNyy0jU
VzfZxTvoZJqoOZlfo7zutpacWZPFfkrUaZRtqpNnu+P1XavoWFdTyqJ+V/liI1mXnvz0N7qLtrjs
0TvV/mbJG68jx3xDileotiSYpdjSZl0Jn5N/ohnJBLFC1xt0hKCkNfX59AVj9Uxu7HnsTCCW8Ven
xt7Nkmf0KQUCFLM5nYt6oZPIhhTKYxWswixR1GfLbaldlPNZ1ODJTtmS6DxOIPytXxziP2s796Zr
uwkKlYqC/UEvci1xA94WNu0QqbN3zivl9JjmC0V1/RmRg5kz7wFU8TT6+J4FcIDSZvpdgT8yM4pT
FTc0FTLcXfYWp3AurZ4rTSJlOMULfU3Z6xQNJrbev0vLPT3wdQ9L2LHCGIULtGVwkY1nrTQYpz3n
MnexTZkT7tJm9D8AqfRXel0tsbb2B/c1Zb/JXIXMn/kPEoroCuHfmh9KMMT06XfwZZH+vNQy5h7Y
TMKC3vb1pj2JJuY3tRLyQoWr3lyfty0bH8V9YDgEbQzuveuJewT5Ybd/Tedms68yCgWGxLKO/U4q
z0nvNRrsxnhz0IDouTsT2WX3HRid/q3GzrjCXo6UpIwaxnGrOGRS+37GF0UnYn9DfPC7w0c/bYvI
rkREvsIL3Qu9yPk6zNnvkbiYsWOjVu5iXpKZN8yRzDucGypExjBuVHf2PLPWiMmm2n+2Q/3zvEef
xQP4TgD1aJgHMmYq4B40W0cVlg8+FbHxMkp89S5ya+PSRCmR4EPOoqqfcOeynRIz8XkV98LHPsz7
rJ+W+S/eq66AB+k2F5iHx+UerGM6xk4jIa83ExWjU11OeVWvzu1dU/MIlhYL02Guzo5J5AzSfUNC
s4NUjLpLhjdn+DGFfY+gh3ZJUIYH3QxSDlpnxWKWqH/bGdAztCraLLQZO8JC7QdRGfo+0xYAHDiv
fVO0LEwtZ68VIPKCSID/dgoSha6DscHoLfEDdsaLnABLZbRxqVe0pt1i4luKWyxhhi2O6Odc1Y4+
kC6BqJF8/yEYp0ta798ibEn/Sj2xtsfOWD63SY/G+P5plRYygl811j2Q6Ang4F/T79Ga2uL2zo/G
G8UkB6k98qTC1TfJYNdyOpCiJ2YUx5ghXa/r0zd9aLflAM1Bsg1tdidc/LYW8g2ONDmkdLNM4BMd
wZPEKK5ijtCWInO84QGyW16aFh6w4CPYbr0STAj+myxFmIehohuvmB/qvPaZl4qF0rsnXxLjrMx7
aoKwLy9JoKodQEKb6aQNXrIMPck27vElrJRWLu9HrI3GE1/oJ+HCtS7IFMYQdcUp3UpIiOMkx3dD
3voC8MG3Qt7veEsgG1l9c7aBcYnjhEoTCEQ8S84i1g+hVOB0/sKAgq/RswHC6OshkO26puquIVDa
tlTOnry6R39hhI2TgaGqez2DCBI3+bJ6Md9PIHuZue/ZkDcM7yUHa4lWUWh0enIOuadjoJ4s+Iy/
43kA/ZCWzwYnkEGwGx2Tt5rEyeerttKPPAZruDVbI3E0C4sOKZsvUQPZkHAGcgEPjcLTeApSRCSV
GPN7lRnvPLceH4h8DLbDK0Sll0pbgbeSD2B+tisWRudLX1Yx025Oz7AHQmHp2bcEq98bW1hfV/PQ
snEO8tlOjgOlJA8y0tUIR6MAbsReLEE7LE2HPUgxdrP0qXZZAmrSqO+h4U8ZfI8et+hIpAM0++/w
EJOSR2hAGWs2tUzQ64eWLpIbdeG+IpkrT3SE2yo03TaUXE5G2DI0yHuNkhNFMjjVacaXeg+s3yXM
UrombCsQ635/hKi1cWHJEe/JsYUt1zmG8hFqklFCCcZFRNj5IuLs7G5DUcGKuthOlzAXakEDssWu
G9NiiszK35JgOdmP1pLs1RPpMYtUGBCCEEhV8SYQS4J3KjZ+eXDsMEKUHz+bMssJsQnFEi3C12za
L+wyat6ClvGTHh/RELVOO3kKH1D6KQ8oWf3VuZTMKJ5j8//IA3OByLN8fEpAanO4MfeOHgma3xeA
9Q1MhqYgejYP6lsJmDmyW71cQv9rgRFPh8U7dPcaksHDuvhqXELzN7Q7o1zO16H2qk2Tl05slnQA
yzvMkxUeI6pWuBDTSO5LjAD9/R8nPNX824lYYKLHD0gHJDF1Nex8OSou894wU9a4Z0qi3StAJ2Ct
8BVT6zi4amn9ZJajQk4SQfBHxTU8CB1dHT6Y1pR6xfjPKe+xiqkQyGty2w0WJUview0icjov41iC
M+HrgVg7K0L4ksplkAmsQPibMJgXtB4XsNfKIp73DUunTdHd/i85s3gk8yd17IjMxpR645nOrycu
80PI2WpcZKGISBrlSaI7FJ3Avny5Atjx8ezKIxZVjIouQsFel98M3w5e3lUOdEE6X/rN+mzuvuwy
op4h+/qMy4otKMaZACZQSfbhmqh3MPkdalpxjqZvd18TvsbBmSD8GzGVem0FhyT/Xdzn0KwidNh5
Sccag8gDoO6aOiYAxpcyAqZGg1LU1YwJr4fm7cG71AvpNjGHwOaCrSB+M9Ze+qAPs+YI9USmM1Kw
ifHAE0Y937tjK24ePIs3Mt/YTZWsB0IHdtOxR+77lGDhd+5JCfVJf/Rg5CSXsaiDxylmnklPRmGV
HX0yWzVRNauR5ytfju6hMXw/6qRQC16swsTpNpgPyE3o8dlKtCtVtYys3Ir3Z9yB3neLopc27Sgn
xPRCQvxQqwaZ/Tpo2vEDAuAvqPXff1vAvlqnbUP6esSnMXpuJnIwnaMbvUREV2PSKxzI9x+JyCm9
zV6MvPyad0K40SK5rBdKJamgi9Eu5VRBuFWOGBrc/jO8lUn79Dr/jLZc+Thc2B/ghGz66aePw0rA
W+Zw9kUo5L5Wejdoa5RISR/SFclApMLIlsHuL7K8NIMWR0ZEmaYE+WFzfrxYco1u/OFpDgmLElz3
RcRo8A98rKPRetPqzFGyrk3vj7Bqej4oK0DljTKEgF6hW0597u48+AJ4bBiSuFPKdze4OXAnjUDR
v2n49iq1Q7PFUke8dijl0IxImw8G9CQoUK/fNvqEWCHjORHDwJGVeMsU5XoG0sZrrTbQqVpDup8q
tG6hHIJw5bGq1LgK3R9DmB66HKsbijlPJjKggaEmrV5mW9tLHDnMm6mbJGt7/KTmE8gkBACkGo1o
BOumDm7Jjv0BYNxM8WnvitKt7wTaatBG7Yg/XNGTH6ZRQKUQCJNdONF9tkrebnNPQ9gZt9jmCaDv
g0MZoIMgCen+BNXDyGSoUcd/q64TmZU9RVCs4Q9Lutnjp7fzHj2nNvPlKHRZx5xWjCvzKe/vV+2v
lfNm5M4ZrldRKvJBiCKJHtMZd1D/Ll7k5LuMq1rJGBO8QrVYij4e6gEK6e0rDVHzzL1t++1jFpKB
ENjT7biiYz3RPKGiQLP+nLgjrfBRNKReryxYntzzUWBA67IkR5NbU8r3T/fYMa7zszpIKn8FRjUG
rzMy/6/srFQvqNP4bZDJCdYGshuGhqALh8He3nRhwsHEM9thrkXIzfi791f+iY1MyA9Ihfs2O5dr
Xv1VTGwoLTcWKd8qam0gx7hMqOEAK3YDOA6+Z/8mQ/sTGk5q0WOZXxmk17X4Qh0crU3iWzpguZms
870khz8JKp3I7lbSd6jw43HBv9XpR+m31/j40ze9JpN9DHO32kbnYkZsGZ5GSXddYbo0RtD0s247
MOrAh8T5AHHimBC0q2eH8Cx6mBpREBq6fnEbLnij+Nk+fFT3MX5g/JqaT/VJKBSjMJaFnqqNeH8J
jYUL3AGov/ROwv/Kc9WwGGTI1ba2OzAkEvEU7MBC8I7f8SgFb6A/e0yWqpUgAmKoXlgLmguhIRaM
9niHGKNP3HXcV0+LZLLiRDW/2eWjOG8EC6ENao3MHSuD3Etb9M4NhBeFkPQKuMYGWIMjME4qaaIX
8sPoxqKhEkWzXcT6rb2dXAJR9FFeWHOYqDEVZLE2a6z6eLtTxI3OJCMX2+HkolEmuR3mPgb5poQB
KN44mMwEwMwBph4USTQyPtA8rHyT4at9SbAgJHgeuReR8JsBVFWWDxHdBcIcy7WkvxLqM0fuhxJs
J03v5BHq0BkkNS5j43BkGXnVpKBwVkbobTHw6MjHlABcWqGXd3aAk4L8xx82hDbqvDaS3bKxixDP
qxcExi9vQ4KNT/F5F1H58gIO6WR2oVeoVqMvKElqTB+qIA1MK5Lgo1gWwtWL2Z1WLzVtzhs1y4ng
DCPPBSgXErsiGa7yi140tZV65Zzt+2JvNmqqiS2f8wuqyJkGB16TEo0qdALh7Z88C4Btj5xzJpDU
AHRE/d6R+Jzha5Pjai6cvNXiZNo5YmldcG7FpcCVLAWlu4sD9e2ZC15KrcDqeyPxA1PiHm1A9epw
BSRmwDCA0/Q5RN5EHx5V/izm+9/6HbDe44eY9JpkG61yan30fy0CPWhZy1ok8TIDzhhh79ps1yar
7GLxeIA0ePR9rMQdsCFKj7bJi5CsgWuvGqtnTU6sU9JEvGLqzCPwy5xnyxMAgHeudf5GyiovKDof
nZIZw6tRqGfZnknI+j2aqUDXmTn1RfnFgj1vNA/3SOE3CaUpxroRA5e8Vv/oOMYFFN+vx3c97SCZ
pLKhDMzW782Lm1V3arTPzknvqtCr39+woBuEU/9zyHQ6gLoZH3V2DfVIN/VH2z+bUTibINqYu6w5
w3nLY4804QOjNyaj3qcKOcAoXAXtsq06lEcE7lGhErvni4xQB2gxcE6U1Qcu/v9wHu5IDgd21RfH
Q1nvshMz2M53TvX9kxouwZDIXYhar6RUkudrNYqld84qTrrRIid3gXIOv47F6zC2WWR8xVeEqOLX
mx+JLWKQhmNFilFWBZdya+0Q9sLzGYTwAT2JQiu/1MvPT55ZXqLneyN3nz8eLE8IDASPjZDbWeHe
7eQbEK1rAyH3nmeEYCRURuK7zs8ijmmNupmvqgdoWcxHPfCLt0f1bTJN9kqtkqauxNOB23K1vn1R
cKwLjChGIIGhhG/szUlgNQ6q+jqkugIH/W/dujeLbeE8bbTrQSpAALC8++MqJGFCRk+/d39uLt2D
SijTvfgHYgdaue+HR51i+c5PVhEgejXMY2nsg20KvpT7faUtz1VeIlryK+aiUVTXAPFAHNxE4u6v
mZD7DCVUN7qtBE2La7Xf8BqRAxqPyAtUcC2VYjWfTezf2fMjquwhSfofsbf2bj5Ed2kdfVW7gSxU
87jH9AzLobZbrFc+Xdyl7PypCeK9Omb4rZ9PsRhVNAen+mMSnYQgwOsgbQYBvN3zJTlFAyQ/nsXc
AeuLVFcVO1xae5S09L1S6axXfyq0bWUYaSSabVe0HdM0YWA7ydFK5ugfz63UXGHKA3Me6LNRl6yG
joKjAUb8y/n2YFFDoBb2cj37w8ODJrqvoYPLhCYgJJ5glZsLL5ZcbpkuR/YkimNezGxbjXOVYr5a
5LqsLYy9d4K+aTDF8PiwD9d6hXCWYFbTifXOoVIKASIoSNEr0sTpjesrjyVWmA16/29WtsVPTWgO
H2MKVQ4/TPwGoaK50Bl4r0fDdSeA7eyYMq9WVm1tuL2kujr8n4BB73x1w9o5GeKwWzQK8jRHF34d
IJsiTE+gUXTN/eZ8rX9mbo4y6IAAWCr6Rz/5hc2f6L+zl8vIS6cJDYA2LEH1+yKaetj6pnOGBXAW
ZC8TQ/sq6rO53X7PaY8AgUcyb1/2HxoTfj0nz11zhUE5I//PYiQBQClmaBaF1L6P4kqu4zrsvLcK
8uK3D+Jz0ZyK+UmwAJuZM4LLmqobZyAtnRfd57TosNMHz+KqvbEbU7DSghhxdQtt+lvBhAaIn8wQ
RAlh+dc4QNt/yVf1YWvIeCxAsl9AM9zbzbwbUzFn0gVFnEqk6bYclE+142V2WouVPAnhABy6zB8E
DCERbx2KXEqRg5HlGWs9GYWGiHHKFm+z6OF/c8ZYDnw/kswIBw0zCXcnxCC4eyZl4mVbUCqOPYrm
r1oiNOKj7YKw5pnA7Cyqq8MZOa8dDQyr33eQMLf4TtcZaQ7gKXPdq/HyPK3iTBe6iXE7ehPUMLMT
ZeBgig9GrJF3xxM2EX+rXP2DhtU8uUR9E/pbkV1pzH71gbNTuaWwi1uBzqM0DKG8ZXITIgqJf/KO
r3zqzW3safgmr/uNjBtwIKoFucqqooBVU+ruD+Rng3ahmgW7bXXyew4k8/evjel+bOsLK7G7sxX6
Bq1ZmXUlE83r1Oy0bYrl/hRYlFfuQ0OD7sPa/V3O4ZnpxXE4tetjYuRV89k8tZGas4pVwn1zlQkD
DFb04o9a6NEBbnqDsyiEGXKUcXeEc0Do4TtKQ9PDCzPFjws0irRjoAd6s9ppuxNDEA9EAYV8J3aj
moay0C+NldnCkBSwOyQdTVaEq0fCKH2VCpGTXTG2EbVyKmLwO/EAqwg23I3y+UV5Ivkc5IQhAldP
+bEcwdjhN8H+rk5+rxkFiG1hjXpOH23pQ7mzopmzKek6BnDpa1SHwUYV3k1V52Pb0LsMQJy62BX0
jVYLrWt0Md/J8tzeL4u78dbDQ4sJNydYvenjoBnJ2sWusG8aRxmPKTrI+HQ2uN/63W0nWrECP0HE
pkIDlPu9q+LGU2JdjIThE66tNvJLHkNgFL8BBO09KbOzfL+FUGd8noIe4DqgrtoXPB3ZmEE96aug
75UtkQPVUHygQ1Hio+fr2jE5rK9h/6x/5yloVrJx6+AlbR57me/gPkaf05kjbFK70Lcsz0jaQXkp
TDULowXMNs3/NTGH17kiaWVDMdCWIpQw0ObtPdZpt70PNneDdUZEFbw9YuwdhXqLb6I6M/x+r9t1
AjR3t0oIEJRI/xdW4/8WTAAw2O1zxn9Fb2joFkh6T3DUvqtMhps1S0RixT5ytvJV1JnLhNcUm777
Eza3ilalvaYYHE2ctbaHTvHroqC9gwQZFft1HERIJo6yZ5UoMuPV+30Jg/JQNG6im3b4tTNiULRO
dsyhDwjw8Szyr3ny9QdgBf5B6VfscKOcoepbPU43fxzf+kv0mMOUl7UYOFKzC/HjAf8UAa+WmmUF
PVNzIQ1FHCSryrSuTzrDpguCKqufAlrX5YdUdd3K60PRQxpSOUN2KkFvgWUXJ4f2/LYFgmpXByl8
ABZeRZpoyuosiXLjjwoP4wwz7wG+EprVKwzO+JK13yeEHmdAr5MrF3GBD2KgbFonCjdXC7ZLlVKN
LyENJQKx5Xdx3mbkT/6YhkVrqYFqLJGvm8bkA9tOBN5FVM1HojOPfHvBryy+LbaNB835WuHynbKG
uAU7ysqa5c7+dDwrtUsxhraOLWqnwPoxYFCh7B6xoDLgfR/8X4MsryqyhBwVeYIEpvUnanmXX9Ad
vqgZ0QaiXQBdt6QJ9/lMSAiy872bnISHYE8DEie9azGc3ZbbalftIG+38wvAMgQtEVdsYxPamtgR
6TLxxSfBvxbt+13gD+XkbEpyUaCTOkw9fMoi5hKqp90cC+bRvwBivL7q/VkiA8uJB2ZgPgvsxEta
iFYe00IO0UxxFp26l6mVHVDwE1t7fZrCEIeTb9U77pU+Z+oJjkUfyVM/vnKarNvcUbc3kZWfQsae
jNE2brYy0jG4yPSkd7wpjYwQrpDHiK2s7gqzlAelyjoOBXrXlj3tLBXpyAQ/naXB4MvRXzTd6t5z
3ux3qqaeg9eEVp9H3JOqODCcKDwWseUh8DrxEdymEAVStP/9oOu3+KVhQM0wPlO4pOXp6cmws71Z
gKt8WelaGSEHLCfbMkijKhDsi2/Mhth3x2QLars+piAjspN5FRkUCWM1hf+mG+fIt3WiUL4qBv1D
/W+6PK2BVy4jhk0VPqUUvddq2P8z/7GdM0/rE7Dr0uzyOzTRplor0ux6r8nvvsGESCTSKP7UxTxx
f/BjHo37Ts2xTH9YuIaKstTmAxAcxeHK+G7je35nhtunKv9T8MYCq3PviGsoXonbltiSDX27zW0m
GIs6MPHRuYckSMPIGPGOJr1U29IeWD+YfrsOKeMQ7IGIlflle9cg2H2+P5W0dSOa2qNG18rkXcyv
AOAIryvwOs79K0Q1AmjidlKPQ98GOxfXi/lTuq8KjLHNR9EQ7dtUUpZfDSfFMWOmpB1MVjXmza5C
Q88N5Ny5zQuPQRvGwXymB5NUO8n+k7FHmHkPBsXxPbvJ2w8pHOPbOvgKkXSARMiVauxbg0WNbQUi
mRCqNtClJS4bM5iLWBALNR9u4hXqloRlm3bgAJ2IOwPMGGvCLwMowk3wIhebWY+mB0XzBJGuC4SU
TZiK2IguY5uJ9jnx3JIoXraiMT3na69hzRegQDtxANr3xABjNuCdJLW9bxmHsFpeuNB/7Sm6sxnV
wm7G7sYUEbqQ8geV7irxZ6KNcd2NIy5FXHsu4EujJmskpMiRoSTbZbK432D4gHa95wpcrqxRwEEi
k/5xGTKkhUSrYQHhPX1Ew+gaxiH4JVI6pabXgHfvgCnXBqNLDWgwqXHZzzt833TGsrEJ7kfcz1q7
ZexuoxxjXAPdjVt4juWcYuHfVphNo2oMDtOIvuvF4ji48RglGh9cqPBcSSJrs9bKlDiXy1LApnZc
ETZ4wWl34LBnAxpdysEIK83N6b7O6qWCuMmKNU5JhsGGOLlzgFQbPOx//MlTPV8pal7DZMwjacQC
Zlx3a2RYcpVC59XFxWnQ7s8XdZC3I8TlyoGgNO1+pMCTiFv5zQv8Wc6rB9VAgW92WmHk1QXB1Pnt
XpwFWs83YLOxGNUTgbN/NAg9CD0k+l8HlnZhNKHUGau6yfMdUNOIjqhDg/cKedhZW2yKlcbc1HPi
JiNhirps9bbwVmIMVKmoeW/hAM1XhbqsLg1zPEZQJVrD6A5HR1FHSFaThF2vg1oeZLSNw8CDSCuq
wWzeASd0GH0pqGzeFHlx5bpeAvTfQUXtybo5j0aftr7BWBt2w4GdooRUeT6Qp4lhVq5fPk/9erM7
Tv3ZTQ2AnORIH58XnDqm+7m+ElcYQdL/Wv0iHHEmpqwL6eTBN5VD1sSvfG8wsrdMcCxS1ROF8jKJ
3yGkO/6haxmUrTDaZIJVEhhvqebP5HScE9SRooNDCIIKM9FUnmKFpr0SIIwePcDqYLcxlKe0Ncr7
SE6OLHgZOKXeBIXoQ1hw5HbRytf4xsDPEX/DUyS3EzZ/guThn2jbMOqtP0kSs3LhSWLr53VL6KQp
oVbjzn05r6Xuf3i3wU73oC02En42DxLsgEJHG2d4wK8HxmrVs3HSnuVcal4XitMGNvRIbrW2J42I
+6ArroZy1NC9Znf11oD7mMw0viuxdMeBkZ88cGgAitftrNlsXJjJ/Qe+kr213DOPxU4wyLGEGa4w
7+VIYeUNKu58qknWwU3n8pb3FGnYNhN/CAV3Exmg3kvH+cFk5h16KM0kC297ijpSYQa5iBrkRkf2
NNuPgWQli5lYEoqb0+9tj0ZMbr7nTTlvMALvYfsI6aTZPsZ83tykdzUUs2H69tXj0H4SNgICzd2I
HM91EPEWTynLMVlZ3g+/y2sM/vUh1lbM3ZwT7AMIWXfVF45Im+sxsEn7UTxNiL+7EG2D1dh4+Ht5
aSGiDwR3koQwZrY5jRppp1ch2pZRGmIpytUhEeRC1sN3hSrMpeurK9MbhQJ0ka3LoSyOA4LL3uaK
Kx44PbNxQupQvANZImlh0zCb8i0IZihmGZYfo1W6Quo9q7c0UE1K9AHPJb94THGKl4Qmo5rVkIdW
OjcAAqeDFYPYXC54THqjvTkkGkA5PqeHsyI2IR3EbmVN7t7lB06irMtSpIjYF+x7YtJESYUQ9VMT
VzFZ77d+C78uv/rjsDjCfSeDo7sL0runcT2CiPWKQoVTaE+UOe4c4X5wXgDerhiwZZb/q+OT84TH
eoi9hT09/xCDfBklOpMSwm2iiM92KhQauofqqCcWcJGZ4IxjsBDoZjVhmEqVaQIBWr4Rd5EmYuD6
6GKWz5dO9TZFH4jsQPodBoWIbMNrTzUk4ICldgJH7B56uzhxAjaxr0d7W2HRgza31Cqy6uYdFWD7
rnYb0ZSq8BTCOQ9oQ6AJ2qXKL6RoGzXNFireK7tzd3BOMk9sYuIopjVSWnrK0FrY5HdHiCWHBq62
/+vFbDGnOILpUIZq4SeA8sNz5K8GRNkC2vGkntU/aiErJMBGjBE8ebEIvgmBcvulQaDyhqBbvPpb
NJ59kUviNuvO/tapC9wYn3d3OMY5fJcPMqTCCubnPPycLp3r3dKBlfvaWnVZLRD3rN1N9X9PK+3Y
wZ7ytM3soElad45M1G6OuaSlYIiJsvdA2+pIgurz69WF9dtXW/tPFwUvtNK8wUXr1qgcvdsqmnBQ
sdzbTWkK+1GpwqfmERqeCM8norBF0S0fAUekQ8EytlJto2vq3ahxo+QZR/cjLFXRsiq2RBwQ/VYu
AmaQHzjjREHgPwc13mL7r81tC/kyqiHSH7xrb8e6Ob1I5RzfNSBDrqCzOOU7GoixSM/y34BiDuDV
yAnVuJx5B2vvMXuAw0+10LeLvH/GGEqmP21UJ753wauNImeItLjD78vD5bFfY/bAduw1oRAmy+Iy
vVYU1CLRlEJ6Y3oTl+BltOCX/it4NuENYlVlaGHYr3oqN+peKLEmjSaR5F07iTvdbby4RDKaa31q
+2+wfUQRpmT+GDdXFVHHOHWomB0kNAzCkrmJDXrMTgxmV4dUxxGcY7k/2CZFX81RQnTVeNLwQ+Wj
q6sHS+xL4V11ta1i+ZGvZd8b5YnJjzlgGRtXREoIBFBHn4zEDdoxSKvKxwGTnv1KkMRp+SRmL5SA
ASQXAXxXLFw+vBEKo/HGzIZv9wzw0aW84pqrmdSgCrHb9pY1z/UrwV48JAgqSnLOk1BpcOMY7KtF
0kgCuLX1Zq1JxJPSbUBHuAVW69fwRqt4PskDxC46dhO/WWI7/9n6OhFmj+QBoOxTSgy1IyRb+vnZ
qZSeIJ5Ho8HpD/Lzm0mT9Ed/co5WaqEEJnZEg97eLchOG3VqXDv2XQrVb2mVXhkxx/ahPfgCljOy
5cgSRytrZIMyOPCh4G9POxNGdAGhfdUXkb8MCytw9uqmUDKugiJ++813tKgX9+RUbMO/dnHIuqpW
QSzswduP0S4gEnQ8tsOoC3fNTqtGOvpolcUCjkrDLGATM6hHLDMpeEiy6iwd017G5N1X1aeuB4tq
CP+/wfAPj4IpwuhO1tU7a82tYXAXOXC9Pbg18N7Yb3GbMju195W+aZ1CPNB/FHCz7NZJ6Vh1zNSe
+NhyZRfk6M19mEZmzSnC4m1cnaavjlFaQK3v6CQt5rpgD+1zeGtZaC0BmIFitNmYk61XrEuRLMpt
qIq7OtBxOLhf06g8sSTzi19iS43oK0biphpK0LiNAcMTPFDgCJKtyWdjC0Cux5kDJ6FoB+Jhsi5B
B71dnWxn6KWXOWSeV4FpviCOFG8JAcsPp8/pK64AXQYLVUWsJcOEsN7iTciKeaLdr6y8QVuyg+rh
igS0jPxJn8kki/ph1D5BSL8Uw5IOfZTuVYgu51/XfqRfsj56JljbyFZw6eU50KPa3YBz5Cfo7mZu
kBJg5gxacYOZA4TXnx39GhNxdO95DoGHriYGpGiO2xan+RhfAaxmuEvbTEAibsUObc98cMS/rCoQ
77lCC6FNq436HyiyXWLy8L9ifphbHUTz2Sw5RQPdWjqCpUn52lZokcv9Vn3lxv6YYksjgYtpt7a1
lPkb/FaHquhiYeM6DRX+VI4yXtB06zrUFkLA9IlfbCrVGdqkPryMwWXnG0ht2gqiKk4zY8CV2TJr
xAhpfe1xXTSsIaVAPS5JNUE8nUkvnLkpX/St9mO5g9Ek6tHI1Z46HktLueB2xtPJxtiwX3pay/Vf
e/Dhpc7i1AvsnH1hgYhRZPsMuMHHHd0lzCI2ftIpD2EvjpeK/kz0ysEiodDSMNtAqPXwNNLDdC2C
DGHTpNzAUyUaBAlElG+vrosSnsDyqFEpgyEZNVoe1avvKBFS78Hjg7jLtxEHFXSqKahAz59vJQkn
HVx6/wbL1f5CgQZ4MphP840G/hLiZ0fdiQsBdnbq+SSswtlA040RgMsw0buGzUp+hgmrJwbcDzRy
dfW874yppPg4qEqQP54G4nH6MqJsFQbUEZw+vBJO26aavl7iwOly7kAN6rwDfk40nyMYUgfncRqY
1ZoXyXTfB+/CEyAJe2CShJa9tlyFH03KntxcT/x/G52fjriszW9/g6TjO/LXVcNTEHTBkX5ZZiJ2
aydrpxLwJUUsVi9n22thMBD0UHuX1eOR9jzRSOc0wdxL08XKYapXPvw1Oap6BhNykxLLYTtVJu72
MdshPoeX1PGnbfk2pZGOPv2PlVutYlZ+Mecb/SL5Ocmbo8lRZ8d5FTxlsIilbTYUluzFrJR5aWUv
cHdDPtTjxTkDAGYQbxoeHNJ1hyU3RyKwDC3VtNd+3cngh8Ge7sD9E/asS5EqhdEwjYnrUdmbIMBB
tdUBy7Fg7CmC00Kg2nqTPyV4Niv8NW10PIwVFPWO3iJQp//0b5D4/1I6lDm3kp5zdspcrDTJD8y5
YqrQyhw9pBhDH34v+pP9P7BXmsAKGcEkGZGtJ7PFGX5Q19V9p2ttFk4mS5quhis06cld7e++fVDm
CGnbfklZi++aQAlfwudBjacPFETfJ6NuKGmTkvBfEO3b5K6uLndd7aqZ//q39fPIBj4VbPeFZJHC
VEcDvV2hxOuitMun/fGZJOQCSyjCZMuhtj00INQY/05nubkOkC/b1kwg+mSZmW+7ECEebCq4FDFz
t1Hcnjjy2lwU5uD9n0Teer8UKhdlUKGwRA64icHHKck/6DIYz/psfmghIjE5JX9x4J6P5cBl1gds
hziF9abLbSsGbot+J191r6XSEGa0kobHNJRJnH5C6qif9mr/I0/AFSHSfCftDAbm6xdqrn3eDNxk
rT8bHfDANCePAOF/ngrb7r1Md3M3ZbACc82vktvF7fVD31b4gV1AB2M4KoaNOL+12O+sJoCqQ8Iw
SZYXHA9NOnuIqqVaKoMfvvSnN6NANSqI9PYgbn8ARFzj/X8b1nts7d6GY6G1IzH6ChLfv9pzH0qF
w9mKHfda2pqJNey4gWWEIaVQ7R2tPeSV33PXy+M0wBQ5yo8KW9ziKGz7cfoNEkAtwtLElj6PkOul
YCKMDtw141jjy6yUkslS0epVEd4ofK9KAHCuiqiGrMU13UaPSVuNBH8n+w+jSKSL1TnOri2sXO+c
sDAiDG2ZbRkXe4WA40TejxhGVA/IF89Y/5vVwsPwoi/DPyiIoxBHK5sYBNHEx+h69D7LclVg/SQd
Vo1SBnW0EPpNxgbThn0PPp++ho5N3nlk1lInyms7cm9lGkKT3W2fpOaY85dGPvfzAQCU3VgTWLE2
eEQnOqyWt4xKyCKGETR4Io+zRUt0ZEp4HFnVOgE1aiObw+IusHylq+ojoWZmudbBU83MIjUTkdA2
1eDXrt3eu0L7unlpe9Aw1/9Um6U2wAgNBGOmkFdBCNiieGGARLrM7H1nZ0QMLVLEBKzEx3jdvOO1
juJtDdW+2vzQ0UphjYgkEaExaa9ablejN6Nu5522Vlg9onI6jYPJOCKlhRhT26MzX2NKlw9uXUbN
4pZ9o46YO1btYJBURUaIsJaFFu0NqL2UR6f6l+oLyaCh/7lHR7L/sLuTGc1HqB8EoP1+sOqZfWEm
Q3ZmKo418jn4eqy/B5jOmaAcqHfdYqAHnWAT1Kdub2ru5glNjOxlKWwEZ8tPZeqfnm6hQQj6rUnp
ZSmOuSo+NIClPZj2zBzTilo/MfT1ZHgFDlkIWQsVqXyYcVD4ZIqCesDhpatq3ie2VlptIz8WI/7U
1sldFVg8/xhDv/hwHm7gCrYHah5oXQKpP9q2LNWZU83gq3t2Gi1smwrVcUAC9iAxBJpBbMWl9o3T
n1PetdnNeh94B+9prvdsujLB8FJkRALOXIVs48N1hBoqugYv7zlN58J/sVP3XDmxJB+xNl3/NHMP
wJtsHmqbDfUFABtVwcHg3aNQKbrOFRsGVcI+DfHFxCHXu9AOVIQpZIgYAAHdp8Jd8J/UPBlZmRi9
Si7CnbkGKIvahagP5GfXYKmK3STqJGKhs6C+7P+apST+zCk7nk9UHyJcHTKbHN6mycz/AHzsj9a7
DsIVoYapX5XZLydIdNZEkIFNr4BiX7UVXWa19W8A1dwLHPcTorzYXg8aoRFL2EMstvfxrTh+JFlm
vlpVJRh0QQBpD2z8O589x3jmLCuGLVvqM2juewPpeqr3Kg46NYwwoTpMFhZzaiqQdWJcTDyFMKGF
l8hJcBpIzF2DXGjHOgXydYRnxx1/2eHsiArJ98h/Ghw7hDMaxtr2m/O/QWYoJubvpNEpMzlJ5Ow5
kAf/P1kSFL5/CpsuZPpau7HO/i6QS8TDluTMePc2RqZ0JF+eNO2ve+gERY10DpsQSB5Nao9ERNGg
EZ8GgQINY2ygIOMiis7myt+1qMVLz3mAI5MAmIZNjZ6cgSQkEWoO/e6fj8T9H/sswATtILVYrUyp
ziPtIPCrHrE3vBUTPtXNmz5qoWm9sOEejTMYaMQuck9ZBanpHuz7mx5gKYxafMFelzWY7xjs4cG9
u4Km6JFibksS9SeO9XXiUmEp/51XjfcaFnPgB3ReATKn5TUniJZfaVkoFV5OeGX2VTMjWD2gfxH0
CcO1z+0xJJz4ZBpY6Njq1cigzP3mRlaTscJUzXWbZ9/VEWe0QVwVry4OUVCZ08i8HvIFOOQDpL4g
K2pdrwGlikOOKCW5bNBXWF2YJQOByu/obmgY/0ksscBOP1k6Qm2BTBNDhpWhpe9XIPEN84jiSKJG
p02MGmajlLFjtokR0gff1x2DaIDVxPKfNPYXwFfcYEyk3lBEdDESFxnb+VABAD5MPbVDxnDqgwYS
IEFxeqFd0I3UXf5j4c94i80LK6XAoCClbVSjovkj7vpDqPqdaowtcd+9dH+WfrcW3riquT+DjXgV
wuDvMLTfYOLH4DqRpo7RULHv26eOtmNLvTtdmAnFJHSXcmtPmdnt68BFkvNDiO9/qTfJgBxn66Mb
QT8lTulIvMI7u4C3GLH9E8gP1QVj6+2RSPpESxWpWTy2t2hMcbCphkEHGdV9o13piKRtrfEcqemh
UcFy2UsrQtgywwNatU5udDnnEY29rqDMyKukOLuZZSdA4ocSCo2kdqtzOGfi2THShrgsvKzy35nE
Bh7bpurHcIT1bR1qcFD+B9U04ulg1Q7Saow+E5Jp8v5dhiVJ0tD9A6v9Qsg46URr/Y3wnT1zBPFt
xQghhd6+OAJG9DNYOSV6B2sVv/t6rWRV7tXFa2KaSw7DdCPRE2l64NT+iVx0MQhJDd9jeJe3zy9r
YSxsfJ5eYDhtlb9B4ApNcqeRhFpvdzHxgx45QYUYoeCi+rJrzx+wTUF6figDyyB6bMLG9Dd7y4Nx
UOmv4cNgrzUTr/fvjf9rveqY9K0knDiQyy98adIc+rI5jzczfRr2HL0Miosina4Ms2Wh0QfaqcjS
EYM+K44Vb3uRUuqutrQbimpEVTcmcH9yG9or4puugtIkyE9fNOlw4ND4PBVVH1uyWQMTFc1H5Jya
4bJA4MiqHIUOpV5zh5ldQvzCU8Gs1za0tImadsiKNxJHHspmz4z0A8oL7oaJaCwJEV0pCwHMiXVx
/aDGQO80rgg0Ll6E2+II6YzQ8L8D/k7B+nrhRl6siVRuxHhvyM86EvF+zohj/gWEFlYWdXAqAmjr
OdevXyKNFMrNiiGQLxU6KMVawPBUSPsQTSoJXnhYGLVEF2jPNQkDwEEBcGPRfUk8BwsQ7+7OGy5E
vyVUdBhVqcPpISDzIT2G0XbusFWFOTJF3PjEmZlOXLM/PiHg5DJDAJM4zt4nRf3nqgwMQtLqn9Nq
3PIBfSIKggWqZqg+3Xr3MrQEC62hZ91s9h4IbhmVVthcXmUP2aRzoG+xgMaIQT4l57+7sx8pkoi0
G0fSrirjAbHJ0c/MAqQOvp9Dn3QtmBHlGC/UZfS69ngd/bc/wcKwmNjkq2X5vAKo9VcCEC1/QgOi
hnnkHSPjnBPdT8RF2Xk2xofvkwrGatbu33Djm34CVyHlMx1a0n5Iy+v05dpWVGIKUx4NHTeD5uS6
jYMKXFRC3G/K9kYcC+zejfWDgU39khzyLo1giEdM3qVwq0nQwYCqaF4Z4J+Z1x6vRdJ4DAZm5lHn
Vuz8UD2GkXw4aU/pvKmLaOhV/147i8SYdGZs5onqdGspgl+I99RYqdTHdR7WO7ct/bYq73o6QAPW
n8nXLh+eIJUUiRVeoIKmmRLP3Bx9hQ5CUxazxLoj4e9yrJB/BPMMZGB9p6PyVpueOcDn/WLiBl+P
8BH1vmLEs15RavHfCLco+MnVGg9u7XUTE4z7UnwJCq4hMlV5zc1Qg5ylQUBV4O6J54G91jfK6ncJ
y8UF2Wnfod4skrKZJ/xX1QhKWjilj0pV95AujMeZN8lYO1LY6yp3CoZnJrJ0Ssl/X6jMTkkVXe2r
qBs++818kYtny3K3tkRU1pk40rlACEN3NWLa8Ovbrn43GjNg9chkmvSqbYsOGCbd3JtcR/8cwwgd
aPkkytxxVMH10Hqty9bJagrsbZL4NZw5kjFt/Tfrvtl26QCFYpuA3qDucjtbG0ItSWv+Vnt9JOvE
68BhRqrxLVbRfTYq6yurly3eQnPRzP9bhOVik05v4H9sur8mwG1qhbAnMc2YW+M3RplfGt8bTUZb
3FXItVZCMFXhyXhHuaQfpVF2G7ZcU8ZIBzOGgaWHE/YW6YkjRjZPZdv7ZtP9J4XAl80u9ZHfdpd+
zkuO5YELuzILUb+9yJgVp3pCYE+sPT5Y58C4kMdT6jbByEFH09k6e6LZ23+FGZlIGxjfCaR1aSxm
Pi4bDh5vpoZQWWnAMgTN5kXTcpAgSCcjEfqAnJygnukaCDhjkubXgprj/nDHqjcyzw61EGV6z/6R
9wRByHfFzSs3HKcrqaR8d3s1GEdwpphXQ+9TfKIlQD6B7Dk6W5GIVQEduqXK9HoSwUftwMJEVWIU
1zZOcoeWrpyEYc+vacaza3Qe7K9D+lwElm61S7h3rjpaS/tfVmxnf2KibAglC9+OcIi+1ce8wr//
1clGB5D67dPUoDsGA9uORbfuQ9R4ys5s4gk4otZ+7iLGXYmnrqvD2w8fEkWCT4VMoekl1y5ilF++
uFDZDJ6790rzAn76q1ikPt2UHI7N+P7T1IpwMWvHWWXaqmOtGOU23D2a4H1HcSZg4CMlf/I9C4Uw
I6BvVtRfDtj+m9ahx47f8DSH/YX3JI5ZkQZdVP8g3kUr3Akwp7hjHmRa7qJB6imtiT6CNX+z+0ju
p8vmR17znjzrOWpsMrot+XJw+Xh/hFd4pXRu/cl98vRoisXUwJDiQhrO1SmX2IC4HhTcCB+QCyST
M+xRMH2R7huR1F3aVeQQ9Keuc6RnOaa01Ikj0HsQvqJvgGkC7ltxnfXJq6VYwWTvpXXcb/16Y6tm
H+AzpynjkpJBAQDHIzcjR9amtHlsOqKXgObgVF9cIUb3slTvhUEMTrVPhju/QS3ZfmjqN4ZyY03p
o9OjGel5mHfKZLN91GtI5gkLZoT/F/DqpQI2/xOfAMczoqBCaSKAakakBIBHbE2ry4t2HLkmPb0D
HOGqTqnf6vrhrRn1j1Dz9YW8E7hqXwZfTnQfN2hzJ8zQzW5bn1h1UB+MonFztDxCGkYFUMgOD08x
MA90frsswDK8iDatqMvoW86Tb5fIcRhwBbfUfZzmQv+tuuUbHayXJup/Kj9OVb27WL0luDlOzdeC
SOy/W8G4thWBFyu6ADSEQv0cyIBCcKk8G8AwrRnVPbDaNTNBoXyd3t405DNsBXUKlG3tPe8dLkU/
Cmn8Rd+pDp9qXi6EC8sccTznFjsS9tmsgGmMVqHDrwCy3P0cX17eYLXA4kro1dYk87ZybmPGHHIT
5k+zAotPe/Q29xflzcA/TUbK1STxMfvGfnqtNCLWON0Z4s2lT4UD2Fs0qV6UQnp7SZsGzZxs8Vrf
dJZWESYVCD//9wQceXU9eE3CayTMV8pslZ1KrxhQhUnSpQSg1zYHdhCO6Q/YKpS7rEGM1tzs2MZE
QYV+UaJuSP5YnPGtpKiTz0tpgyxMYo8MsMQwjhmM4Zx8y80405x/y0lK1qGFxbFS2OkEOUGU0ma/
5BbFun7J+kBoWFjf1FPv4kPawCVuwLom04UjEQCfs1JBPwGjiGfjhYMB+NjBc3UCN6rIqQ5MA52X
lomw59Wj9+5eDGS3Q6yfzZElrdUdA2JV6pmgoRxra6/DEtZjhAxlnVnup9fN3YUjkN62x6WKcGMA
/Y39mSm+HKQRoT5FWhUnuE6kWQjKYF0xlw+8U41M0bodYzxg0zN8nccaw7O0DgRchmS/FfG+Jggn
pj5A3qckJfLchI3z7P4tQM7VjpsjRgvo+fuDKNiWsDaXNiF/cVrPB8CJZyeaO44g5XsXGkWAVMm/
OHXDSVXkE5d1Ez5vB1EPcXjpaTROvXwjmOv3o0u6C0oOXKXgkDtCSCG6fKHJcCG3wPW/n5S3rGAM
lp9r2M5AFPsmjoZE5052qAY9ZfRJYEg+46/jpcUkUBoaHbxK72G5uPDnB43XcI3YqGRYKUpo5ZxZ
yz0+PXdYrokp4CBhCdExhscqWMbXGcX3YwAI8OHOsj9JdUNs0cOaR5FUd9p6hS8QDZJnHyJcgPdr
swDz7TDkwbBUwRPSYYkzF/Jhn2QI7htqNc2LvXH+5JCjkLJVZOIbD5167zA2pfigGNiMFxDvPGQ4
xUrUqYtlAds+U1txtt0rsXeOalhAwUqXIyXvf7camQ+CcrLjfab3yASKX9DhCKT7CoreqRxcpKNQ
FTkQS5mAvc3icLe+OYJpG0b62hSDNLBhBTMqVskPm8YEAbD7vq1/qGINRBg92ca8vvCnAlDoQ6LN
rXBj0hSsu2CimbHUrh3npKvkBueGw8agMxXxUlg875s7ltPj7uxEipBAHF1ZAtzK09VVGX2rPcFD
qNYNe87pjJc3N8JmWs7a6q1fK4bJektGaDLiNnWH2bbviuml//Fn6AfOA6UkBXbA5pM1ClZEQBK8
c7h6fKJGpjZWXWTIk0Lw5bSCsDrXUU2sBzeTV98UgSG/3fkMDTSppXmr6ROD7rHrt8Evnd14LDMt
b5nCLMkqHYnDYTuYyhxgijm4XYwt6I1MDahBIfPQKAa9D8m+RumIEarSX7dsxjcoq4kHWDaYYU2n
WvxeJrb1wgu1dYt2J3akXKUfi7J5FOe8VTUV+lQsl9ogBcVLD6Qt+TRIHPfHfekTC9F7cftSTj52
8+B8O5FX4kp6F6tmWQQ8GirNmQXObFNKdoUysrdPvQ3ST4CB75r9G8c5re7tFVhgRLCwYrAr//q6
WDNiHcsLdTx3qZ7G0sMmHIVOd3Slq1bXAIHkrFmY7co/I3jyiuEDo/vbknTqW0VD3dkLZUBdkCzu
PHAykjuKdC2cp5RD5b4MxydszzmjargnGQIbmPNzpMyqfx05na8uoHYpAOZUSer4bIQNTJqEEahf
0u8FCvEESnMhOVjZsc/sw3BM+ShCz69M3uhtnTYXN0WHHhYu3IXNex4nnTysw4/aLr1VisejvJEF
exemwC5uYTWTqVsbIBfEICTGhV7yWzesS2BPK/cOkgAv4by/IfXXmrIUEmB35EU7UScUqIUs6EAv
9+T/Z0Cv6pYnlS4eQW98VXmIjHhM3UelJzZvq/0h03yQxnbGwzMOMjgZQbReKxMCs7wfjJsZ0/tx
Js99yfJwt/tgoqjARCZ86Kh1+r0aiHL5hnV47aiUasgfl1tC4fKWfZIooqzLsLScJmhHq4QNSaGQ
ildksnRnDbKzMzxJTrWnFFs5OJuRyl7I0i4rqMdSiyJSXZAa9/sJ3yafeJi4rQzixjJtAxkhFHeB
ERZMsh4KeVvcyl+eioyVwACCjA79Tki5CDP/4CTZATMNuLOtyOxfRovHK9uEF4XmpqBswqnBajE6
tKWotz3KoKgLsalbIgn5Fg2gQatICzBrMaFvUBSjAc6dziNkKssZOyLcm1rTjDX9Y5S5bb+2Gqle
Bgbta6J4tWGsAcMRuh3QztPGArLIJIUG8uwxX0j6F9T/8u5T8u5d/OY3vkmo2S6BIZljyggGsKcc
xCxWK2jkyL0rPxTjA0DIU5kgnfXG5Aky7DDWiPSlh80CYIwqAGq0DjbTFB4Em8zRffausDDEgyt3
o1FiGvjKE9xz9krB2ygfK9SlxN4JZ4LszINMXAimR1gqyesDftFmeKtbHW7QTHACDa+xON3aLWTN
2K5PT8IC9A8TfzjkGJ0bpSgrbe4xljgPVPd7TLUVyFQhnytmUfJqtdtPX669tw/dKpVitjsea29Z
A/OzLFQDstkcBjJY8qDjxQcPoTQKjXLtFYKcyCRlFwJe/O+Z6Hn/XGdBkEn40EB3zqSiIAjvSsYJ
VEbHOmh0oAZeZsd5fjuEyNhar5eMf6Tos0uf646c/e3YG89kBoivhMQjb6TA88KulVP8GqFUHF6m
zqLwxLCYnnkuAfhMFbGzu00bgioFK1hASs1ckAA63uWr/+/rZrYTbXHXYadJaY6Gye9/UYkVIzrR
gjAHeCGk2yEOcl/qx9npVnH592OF8H1u4Army/gLzjF8msMCSrSAxnh/AZAc571z/+Y2bjzIlj6y
tk/gTrC18KSWMA8v+aGMY0iHeM8AFIrB06zAAJkhAhvJDbDiKByTKa75qZl/bCm0w16sfirDE/NT
CYGMgEIn6yAJeKznKGGYLwqVkEr1ZGgVZJzklJHK82xNm43wC+CvahXZ5K9QjZ09W6jldF333nyU
rJ2o6EJuEUHLEO0UzwxE5ruj/6qF84OQHDZwecLIytFT0BjeSbn/XGq9ThD7W5jN3Cx1m3TlpG32
X7IG2Jr9U0j361WZNyfBOK/Ip0saECop5gXfySUjMbV5clgwXF3Fyts/5FeGPM3prPpoVI1aTSiy
+O5BSwYPB+YqZuIRXTn4ikKowCoerIG/aEbT3XZ0rLn/1rz5mJYQB6Lp3a003FBlEFvortCIdbwQ
DqLKxGwXSvLMrm8H7/OBF5/hcOdG+l2PKxKzDhszflp+oSwFw24jvfZ6GpjeWebWJsF5UXv1kHe9
W3t2RHu+wHVFMz2Pvdwk/4ED+yfSPDFBSyRlp4sskiQsR6mjSOY45wtG9SmdJDyCCwU9I0ceb4+n
afSISYB9XV77Yl3ryXgXank+Mm0towGpmpQI6g0OxSku6k+maGAVQ8Wn7MP7csWoPGhkTATPbwFA
8/UWgoSHcrDdUNgbkxDfwwVunADSHTckXw1EQEwlm1N0QJ2leuCwbbNB9K/2sUfx2Lxc2upxP+JI
yUGtbVVpdQQEUGMk0JDG6rbkvR2aUiIaxM8itnC4Tc6eG3tPwzWObhnNsBxWTRZgyDetNNoLvF3J
CtRa2kyQrnh1THpkrsfOWEoAY+7DfknMHORtTGrx1zIRKhoQY9N+H2b2W6ENRQNHRh21vzxZQBXm
ZOCr606JV/gT1mVjrBN7S5dXuvl6LzSzN5YYy4g2thm7B5048Z1IsAUvvFrgW2Gfm/M1s0Q9Q8/Y
eBLHPV/hrRLt4hBPcB5SLBQGr9WsH07NFs8Np1dOf8pO0pxFrS+BryhIw1Sc9hoB0S6TBxz+WK0i
ZwtSvDv/d/22movSj0XH7soV83nw77fuf7GCwkypnvLNnNPd52HFUsE1VjOXhEiy7ffalKibbFjm
i1IdSxUOnJKUheve6z1qSSX89LH21ZCoHmibtb6dE/F3laPICfuwBn5XYvuoOBYPN32QgE5Vzm1F
Mq2AmYbKjgJEj4pnQ9TwqLcHmBgRep259CIaFh1PfYJlcfYJTMZxmmyDvmjMCPWvihuvrMSRIIS/
oQCFgHsKCJKleEKU2GIGhWMRU9bRpckcTGG3uA5vz79h1tWkNDtDEAKXdu8zLi+aZW+BDvPb5u5E
kiFi8qOV8jxOqS94YxUgzy4d89Ve9FytHPZctRnr7wwfrMpiVX5Dc4JGJVpajHXpwfHaMIVYEhRS
lFH91n+TwoiGiniDmwUzgM1v2qi3gDxBCb2mQQkbnNu98ch0IgPW8rHCtV3gLT+oInWkIFV2ztv7
WTUKruDND/XeacjOjUrcHYw7Ru3TFRwXnCWh+DK0yah0Nj8ytJMZ2jeorIK8gBPsmqszts++72Hj
Qa0RqwN+vfmbKbsKfLBOs+HHJksGPb7Sa57XFpa+1gkP5HFxXczGW4cChSjSttHmzbkCfKPApoFU
dYHhWwbQP1SF4nT+GqU1FPNycpeZ9PEcaRAwSfTDHTdh/MT7NOd2q5XMQ+4wZo0WkpRFcalQkv2O
DhSdWCTu9c/e0x7HmMxjAT4tl40iCBvSdS7MfTe5Ytwin/0jwFi5e5dlUh/q3d0O8xn1Xr7AaADI
NsaJnNOBVQ7ASJ/Fzi+b3WlDq/8u0j5cjTBYCUy1ILS9RJwI4ct5CMhWEfQ8+Hbk/+gUU3dOYO4y
Vr7j7QGmLCOvJsHOiRQLhicWEaCtBixnK1pWYiLarxGDOPYj3H8hvuhVaAyZbZ3e2pbDgnnMg3DI
vI7N8xPMvjgZyFk+21blIgKFXruf650lcpZTB4dBChagQSqP5CZ4YdDoZ4+SzWlXPRQXX3hfgps+
ZClDc8Ngso23G3DQH4KKzroQ5YRXPvHsL2E3TBQBqcXbummMlh7+g7M3/lC2gThgPhUxgLJ+hfJA
H3JuB35gbNdKHfzswAkRq52B+sBb9TdOhkt1HBOgGXbrepULVLlDCJ+pqGC4OnHSM9Hpy+No25xZ
3Gb8vuLLQCdw0DGldBGqFhDv54FLphmIWeaRkVotyg+vBiEIJz+Fzzy66pK2uUrbIUP+TDLNaqDG
yhW252L5SiCO9lofr2dwYWsZdKeZL4GuE7X3/u5OnmuCnm9YwkjNTFbu/ac/YyQEl7pOQmI47ErZ
9drkGObt5POdu6QQfN+EWgDt26qMtMovvMGt8YcJB8ApKUOES68C9RNngdWwCaMWo77cAjurRp8X
wyyLxzEWroh0gvg2uaY9j/wlnAGPsqkdI+aDFk/4lKiIKFbBexAIyBjLFjOG/HKzm6LqGpaLG6TT
4HeR5i3WUhnSL8+qt52uSgLqOa4CVejOoW1YiU/VMSXEVCXQ7IguX1PBJo77niBTeNZugzyA5SIx
XgedAfjnLbsVjsXxBOYXSFjfpoHPQjVsX++4g7/3VZ2wZqLDFblT/8nXNF+uMENOlqfWYw7775MJ
8sT5ZPL5MszVjxK0aqv+dyF9e/LbVSmoBmbs4D3IpwJy1ReIbGkCmsh5rrsYOwldUqFiTLOBu9f0
YcZF0XDGRUsl6vHyKTVkeBb/AUZFPhMKd1kKtHiM+csIM+/o8NH1GSs+VSoxGdptddOD5+cMain6
vv1vYHRUF7zKUyE1KYKGdcF3V2gqoUIFF3CCW8sHVgfxFDcDW4CYgliJVSAvdbsxRMT8VfYxcZ7t
47TCjDE/QX+4XZdYPPEZmRg2CSumWLtN2RiqjAqMVEtneDdN1wKfqcj7Y+avYGwhQMy5WZyQ2F4l
ZTrc4Sqlz+jXv1hh2R8XLlilXNWQGwKf1TS+6a8OqT7mwEGrBZzILVERZm9iBsm8PIgoY6hvvYaZ
2m6fdIj7oHW9wOUUJbvtcrQpf97r/5du+KdZnQ/z2ErINJROb3OmPYO1Ad75cvSyTbsHVp4F210V
gI8VnOlxtpL7BI3f868IP24wQug6dhhrWnnnVF7wKibvcBXpFqjgCqkjLeQuwWiiHm7nwobK77++
+VwgZA6r6yLwdwdQvs2W3/O2a1Efe3bqYQqas8RA6GIPQdu0YD6gkd3IUty61DyajwNZYryQEjCw
jFms8kWdMlbcL9t7UEfdvcGUu3ETNSmVNbUOnhYlVz/h1NTec73sc/0DtQsHeb35pfg5fpTp/k09
dOe8jDDWbu+LnkGtbAgnkKDv0opFbI3raJH40cWuA7XbMgf/OAv5L5okQp7Hjk45PdiMOJhBVnKX
5+D+CjqUl7u+rHkqlLz7PB/Dwb1qRW0uHQXMTlU1JaocoLbW+BjwR2M3w2MkEiAMRIahDMIiCfXj
zA0SoAVhOhIGM26WDuesyopXxvM5HAVhBIFEQJNLrZR65JlImyZTo0yAPEpQcbbdHbDBOegrZHfy
QMbKzoX5xmIL7T3ORc1taa3toOUMKMmOmU+tnfcKBRFzjoWS6Vnabk9II8AK/M19Ltes7VA5rPaQ
htOwndk6gmiYMNkygJn+bWdA9vHpTmHBD2lUr0oblUJ4Pb5zSeQ03TtF94XXFe37qpvYeNCmGl2E
mvhEzyJgm9Qhv26sIfraxYXK1b2Iza/NEF8dKpAAmCuFZ68P15i9UiMxbJAUw7E/5SrOMDUKQvVe
8T/g+ZIa/H5TkRY2+sPlp3g7R+P+N+/Gu6j/Yw12aQU6NkXbAvFTTocZfbl6er7KzymUeAZAoHnw
j3eRJ3W1+kl+jnl6ywaXr1wPGB5tPVY+jOol/f22xu59xvkJTmc2z6HJkb4Us3k3vov17A/Sm15D
23rE8vRAr80105WZ5y5y8T2pSPU1zitWjXc/miczdizoqSFCYwqSNALfyCGSwIbIOr01AOPG2h6a
hJaPLj91tV7u4Qqq73OAZxQ/G59LqXtbusZNOgHxK4FglTZ54q2LT6LGi1tx5hV9I9evP86WN+CH
fUlFF9mdgR4g6t3vUVPl5YhNvFzyL/REKv96I9YffUKCMCNoR96o29cR6YtOHARxMtKns0meWW3Q
uzCcyCFIsCTMS1IZHk2XtjIM/KlueOiEQ5HOLO0e1o3TpVe7bXPg/COZLQDVzRn99IRZIB+q9gm6
gr2Sjf5SHAuw1JJV0DudgeDuRWV7qbG3OWSTORQi5+LFdh/lAKsF3qPp6/6M3RMHblw/NbZgzmc5
rMhgd5F8jWwZDximspu+ANg27J+noY4xuF/hbi4GyTyMNUxHMjnyxhlL+E39TxPyQRy5YTKR11Da
b0sA4Zb8Q9CN55KWeMQoY5WD2bIarM2rEqqO4IzI8zJftnzPGJm3n2sSLIIrUhPuJMYpBoTii+Ht
lsH41BsLvRAUYqdDmmmeS6/jH/1XVzuHkkKvSPqpGjzDIe6SQ02EGTqjEmaybanCAwioQCQOKnfM
zxr/++UlLSpSezC4pnFjYF+QndlesspRuPAktP3RG76BUfjqJTqkN4ReHryB1XM5GvIYJSAA9ueH
gYaV3pHglhRMTYFycOAmrBm6AUL4YIaOYlG3LWySwbw3dCNyrI7l4Immju2ibbBAh+owiI+c8Qtb
9wKaobZQVeaTzM1s8ybvqinzBjiVKuOHjN3oq7UcL8SdoZPTm68wdi18H9Euw8kQJw09BhTAdiyR
A310FfF4QxeX2ACqrxxwC4gAKdgbVT3ZggL3PhFWhU0Wcs99dUSa1VGs83+2t7RpFU6Ze0CxJyHj
HEcws4X4sRD4K2JjjLEQj13nZCuH48yARlldi19NU1Tp89zrzyUPNS3B4JZe3lG+iUsY6Ci7K5ww
Lyt/HVj6sZWXlGQ3xkNYM/c+9nCByblceg/OBoRd5m+gexDcV6VLQvjwLmX1HwmPV5WSja1QD8sc
WmrdkHJ4zSnOrvuliLltmiZCIGbpEJFgmlL0BFuwwnrLcQaR0uyAYnTa77R2Nj/zRe8z3V35hSfF
N8z632PbrbiDMNyWMbIflpMkgbtRQjgjCE+pm6YX/EzSie+Yt4D4cCMu2NSQttcRumNwpZglgYvY
Qb0pvD4WJUjIr4SIcGeqU7DoRmG3dWQyGG6KGtupwD3OHehqjCvh2BQQbI3c4qvf6NkHOp/8sFc5
CRNXRESnhqW2D7JfccdTN5HCQ/0Jfq9tIGfWhatgIL9BiH3/xca09aKm4ntRqjbAbUStSy3xvfMW
y0RiMavs+F2EKJNmGUsEF9oRvI/0m0R9Spql8YQmyW4TLRnYnF1v6KNz76zMu7/2/8dVxtUT0wDx
G3SIOqo+bBf8/Zl0DqCKHOnb8Aew06/k00HHFLmY/l/yjPGX66V92W1IMdpHUk9EEA1Z59HwZOgM
uN6THFMPLdNVTgalsf8UWGTsMdMatJsTvDnkoUq+mYg/1e7d3NEVLE3iK+vuYKIrNkt0Kfxmg1fO
9/K34lVM6cVDMJkV8XFcPtSPAB8moLnKNVlGr0YHXSt1/Ven7hu8hHasSjh8dUfjbBWGoeIOgfqO
kTBlYgXLEScy8aTIh9xQMu9jWB8ZuDH0FZ6amJc8Rp2V71L7t3dZgktT1UYM5lK0I+RJ/5RVWAZ/
NTrldors9Mbikfs/jG0/YH9WZMNZHOQV6u1XDz8WMfvS1b1FhHZQ/JOxm8HOe/Os0Z/P/GzAXYaf
+v/u32kJR4a3cfEVI4Mi/GLfiCP1xsWk7f1P5Gqq6o1m0nt0EIovedcQ9BIvh7krX6tNdv1OU6OZ
/bd0D46JN4qblhf1KmnV58GTT1tP1HD9FhPotgYh4C98mAzmmjpzaNggNiXRmSjoEW8aJo1P+ax7
I5HVM824cwrsCRtLQOJE60c+9HzVTAGG5pChOoc9AOnclR/I0DOfWuTVs8muKVRhIBOlUrkTbZKr
huDTmi1x5vnoFiUyjCQi+GaXsOTv/ysrdKzPZEQahe3iTaePSMok+6T65zCgoTBhmCr1LaleDMmh
npOZABaGzUDpL8vk+bYmc6mP0uGrRpxbiqyxlE2CezAJVuIwn3OE5uGIbWjxSugcBpLR/rMSVBe9
U3iDnsyFdf9etxJiRjbEq5PjBJHT5LjDI78jyjD07UUl4xB9+WNKAw3SASpCSfcQLeSF6QL7wAVT
RUafXO9sLt1he9y4l/vyzKSQHb8yXPQa9LxENCjUzHyKXZOTVdg+ffNqXx+4UvqHgLARiIZqy8TX
Ng+6fSveMDzcianGtzo3rvTEN+v9MFFQPdp1Y4xJ/SlVBylTMHK6kSpQuHrQYv7gynprE3jbFdyk
TDrym/wU65r3EDgJDksVpjXxlxn28Nms1htv/MYquhn/2PwZ+lzENVRoUIZzTdw2X3vHfA3MwrKt
CX5HsoyguRjnMc8uvU9CGTqHd83hqkoPbH6YG+TkCxwhPtGGXUZPOrZ4+ghHUPa/sJlzxvfrPVHV
dI9Q/p9rFb0cjRCgz3u6HvuEiqbzoaibs5wSOvQpr8jEXs/O2JgaNlUh1tFewygDr7Jsw3rvg9s3
7T/bAtCYSywWRQydEQIbHxLoXCj9lNbqhSEvxt36kEqrEbOqoS2n9cpkHDOHAx0P/wqpjybRHVGm
9SUBK68Fg1btXRy5oG+UDNZe3NLF/G7My3oad9PrWWv6Odl4JfYN+W2+Iqw6cYHIUOub8mIzjQhe
AsbANAYRRuThLjowS4xyqvSlkjNlhYgmv1k+QhVEEN7NIFP2OX4N7StBXrKJlAObmPs5PHIyNbU3
VBqhO8RlVNbItOwf8sd/aQkNP5YfojGfwPwBs+I0ezLXjSRcDmuHAzfd9eJM+3RWd+yRG2ZKsZQB
2LjjkQIsSqYzceImGhhvvvHB+IPQGOapMwwLJEvqSBhtnf5/nUiabFYh6Hz9edE1leseO0okMIcm
CE2/JJ6L/eLV1M2GdARlXO5PlajzdwLnjj8j+9jo+Y1gHx+b7Kz1TIDF8HJcoupSG2Qo9XYD8zeg
eWekKFNdeiyNAA2La9cF7PPuKQJlfqsx7EVy6qpr7HYXHwBSG/jT+QTwCZK6Z2OMEF8n0xti8Hh0
2mz0RG6Jh7UlOInM1ctArCJUvqg+uchMv+uH5m4sPMczOnC3gTb7UFgz22LEldZIxOn3ySLBDIQL
dkPl4yA7hGffKDubsENdocwVovwtwrUcqFUuCveRxB+DHQvlJ7WMQcK8THpJsdwqjRE85j4JI5po
LidzSsDqkDPoqZ4Oh0I5Gd4hwkYB3v9Bnmy1dwNaiOpcL511AgAZ+AisLgFwYaeXAeUb88aFRmQZ
L2Mheom6dZV0S4UxsxByCYdAz+jJtZTuFXLuzL287Km1vlePeAhdR5VLDQ3k/gjhDo8DwEja4hj6
8WSBDQHhF/0dctL/KQeBrqE4DT+u7xrQ715pKV2L/i4Zfnb/czdCCb6lmr4xwRAu1QylUC8aKGdj
IKOI7a0xJ/+YA9DOl+I/Y1YrXA7IqyKU33X91fIARSUNquCJBWxVo1JUh48+DJ6nS8NUUU3I2cdI
/Gs7xFlktgcJBCTm0rxYq7e1KUlKuzcMeV+D7ZRAIhMBvTgENLnArOEhU6TdgaaLvnVtIy9glMew
/0OBHSWjcfrvTxv9nLNEPaxjS5aD1mLE7cLDuxch/j/32s76O/m8ezaZ90g6jHPTVPlOtX77sKQp
llp/UGEd/UF7ggBSBfNzCo1rsqQduLm91iRxxkN5D2FgxS5HMGMrEyO8oUXfFH7SOx03w193N/Mr
LYNDUVyN6FEtC7Ae7Kjsb3dK+ec0NuquEsid9kRDhOzu+10eu2ryljHqbEOsLyE8WkMajEAnGZ7/
JuWGHRqP3Dsgw+pXddVf6PjMVP1hiVC15bhp3pJ3mHY74FubrNA8Fte5P/LoniJ4pMPiKavZuIA1
78bauhdZFOEWRRqtReLq5Hby/VAON1283FGm9mTtrcG6VDDhGOgK/fUXLoCBhC9zYfNczcoYmu86
YWl3FunVQoouGObYrhxLkaKN3WzEqV4HW+/LjWAZHCthdqrdGpHlONJD4zlxgWg6BSzx+Ob8+X+2
xvopRcYPmSdVAhdUjflgRDeSE8RV1gVXUIqsA5iZM71nIlVEKScwthCznpqc+imHLRBZDx1vOD2k
WrMJlWIcCt44zUtK0ugUxtIZUaOa8CamBUrKCTmuUXnvsWB1cRFy3uHqmVsrUYwEJdl0MrmIBfYI
EN2AGLxodM+XKoRddIMF6mNtwTbGkQ/wrUi9J6P9AZQX5sXej1tkKvZ8rtkr7TnCaAN5FWwzVICZ
hc7m++SKEzYrePckGRlfZb+eekVbX6XVnupqbh4VhbAhDvK8PmtTyHns0IL0AQm3sO92qDtnZYxo
zZ/xcxpHAJ3ktAjyaxxcveNcX3Marw9vd9KdWyPpAlCmCTPwZr2lyKOIW7i0afhZC4w6JHWJb+zI
Or6/dTbLraxUzUN0tC7xijpRC7thuzLHQj1HtW5w+tOra34UptqNrZnUaoKDcVkfR/j/fJO5LmR+
hzhAhnfc9+RuNISxdFrPhEhEElG3PDCUe9uuEk7X3fb8EYY9iD2uIDPN/GnUuFpWG8BLHWulKg+s
wOQqMP+HmwjYkd1SXzxZzYArR6ovPahaMb1/nB0+6BSLh1c0PCea+ygGmV/9FqWMFuoT7uufj96G
cblBWDsncf2SAP0uHKpom8yPqmDz/zbe+9+qFGseWX8GChxN8L+g8+xdjHthehahSGXoABbRZC6T
l+pDGXBb3DCeoR4Y17XCxXtSjDu62/m/gCM2nfKO1FDK8hMJkXQAHgfPx6yjLNc+7LQTJ+1PchnZ
/gYHbvMJY6RaMNhHlxFNttw4NHXXNLUDAv4zpzFiS/7H5RCE65CiEfA9VmiV5OMkxypu3p6LjsxO
j/3jqtjk/NnFORLccln+mgxweJ7vLV+kqtSchrcvsJx9QaBrCgDpRooQ9AUlf5e7v9ZSC5Y6hWTj
tvyEmYuM8YTKcGumy0f184pfcdAZNAmXWuyzjfaVzHmGQcmTj0+A9dkNDc7uJrJFzdI7c6qLL0XC
Qyv5fR5EtExBA/+DXtvRtwIv9bQwz2fTD6yrsoZI+rgwdQZAniingOOWzMUpIWXGgXJi/JZ7RrAq
tPSxJO5d3T4GRx4ZQEbRFp2KpDBUInw8NYA+snlYRTGCZEfRk2DZmsQ6J+3cexGPhoR3vrZIHENB
7P8dhpbR+zQhxvmClFHsTle1TiwilA8Zu3k1lTA5DCKXgXLzqsH3POs8s+fITI6Bwo+vAZ/6JHZ9
qQnZ3fOKFa9wKFUvZI2dP0q/imXHREB5JqISjEcCJGAL6j5rYynFog0xe1T5xlazlo6KZyJvkvq6
VFeUb4VTzBjMJzDTheNbz33Dd/B/sJFWdDK8lgfj4NsWi/Jt6Bg+MqTsRfNFqnlTTyiuWDKNKnKm
6Y9vUjjNmjurKPHLgk1Zb6JyvnoBao4rbi11jwCO46w7t/FxyfVlHAFj8gYdB9pnyzKb1whnmKoi
64y1+eoxZrZQPl44IEf6xgYtBK1B1RF7Wpb5SntZjxpI6TVRkHmg14EJfGHcWmnRVWGBjkzaj3nq
irkve/BW9KFWV7vZDFVWl/8tPVv93OD2WDVXV3sLGB3Z4zKEw4gdyUlUrV+kmxNLGxiR+0Bnu2lQ
YuuS4wsQqP+BjNcYBaP9pyolA30gi3EGtbatzuX/ozm5tNWwLfZzHuRa7/WCy27MPGKQM7pdpaiP
QZYcDXan1xxUxWd4LYoH58XYiEubCePkBTvyP+1XSV86euyEQq9GIL2UVGzlybHbR9LYTNNNIyqi
z1KR92L7NnIx36T0KrNWtvYCONX+e7Aqv/j8holvdpqRH/ox3mXFYtC5AYO1rT6MAzgA9zP9YIe5
oaWpX0+9EWgG8iLQ1PCzZvYl1AS762HoW99zySKrBXz2QcTRgW4Mu+FAMBPXMCI4unnAxDzhQjyZ
3LhbgK+O07bseHYp745nSjrcAwOr38zUMRRQITKxDMNhqHChJWqrxWrzpmdAcnLT7n79bamWyFfJ
wqTexQjx+JxuWuS4CE/SvNZcddjDoYstN0kZzi++0MZjgV2j4Fcn9ZdSoeDywYEkIsDdiDbfNBot
1hf7WJcFZk6jB4YGWHVRyOr7Y1dCt/9PGLjjvV8JRVVJTa484x3l5yF5cYRqRla4AtY66b8CCvzo
GF8LZGEMws2x7MHGM4Ly4Mk7Q/6sfMQOhRxybIWDL/scQoQTJ3r6OX30iENXENMUcpqOqCEdCu7X
Ffk6T01cb88b8XPL82p1zImKvxLc/8ho7MgCM8uMRpYxw7ndErYjCNwMvk6n+v14NpLbRMhQwvYt
DpmIiDhfRNSICLAFxoUyKgBxFW2QLC2rvCe9DL2c1eTwdIxPwuffHjFR+DPC1Ks5tYcUbIkoTZzf
2P15k7m3AsPh0nBa5SlKD1cJtosMg/kz/qXlzjaXHsJLFEAMgmGZfp9AktENeOLQiXBfQXqwJKpa
rtYVvHoZXxobBZge3av9QOhzP+F8ElF4QV8WCITbxQ12Xuyb7o7SL06+fVayGVrBm/3rLDjtzYZ4
KUs+RftTSpeuG8mw7JPmVJstPgy/bLOb6GeTJFkZCrug0ZF/M6IE7mAmjL7qDBiwLWUEMBvqN0eb
TIvsfm49hO6JRvMdOJRLtI/vXXZsCJT1GMDJyuIv7NIvrzWWVxKHB/p6Mkhd5NhozRcliXtYlLp6
vhRsNFFOYHJH8DLio4seLVI0Nt8+qbRLv4b2/i/vD3oGoDlI363oe9Q2gt40MPnCl6TORyx6B5Y1
3tAZMqRi1vcEMTZm0WWcJRiUgLf+tmd6wVvJoGbpi1VD1Yn58KsPGJA3EvC104EEbwssNV/Un57Y
8mDrC/831K6n+0QhbLoiRP3dt72FF0JVIA+SkJ8UPSRCSliV49NDArJwAQ1GR+fL4RoFXven5O1i
8osjtZHIs0k/TFXr2fxf3iIkWwBhWAl2hZZ3ZMU3IMCAIcU9s95e+yh8N91jqzyz/7kkhRan4DAo
6MVEiIuxaOC3NqTarc6Mv7h/87+R/L2jDiQyrPg+LDRdrmCsMLvzwxLB2bSXZyLKORQIoltdBv6N
79pdhpiG+g8013yQu40CLH6D85xc4dG3fQ3+dT5rJwSJfexc9+nVjNLTrQlH/Jnrto2W0d50ShsR
Sm6QZ5LY7eJNZ0xnCF9oq5RdtLjv5+XegPKLHJ9stdTYYUYbzX0NAHSf7W5RfKJ4NrLErL3p1PLG
Wfwj5TFqrcK/LktfjBf1kVaoI6V1EvJOjuOyLRY9Qa+tByl4Y18IIfu3KTpxdISHZiMkCpzAM1Uq
wvsWDX8gNQldoe7zhsi8r2v8i2RNccJGzmnWNqAA4DrYEGkMLmqaTImZT0W6Y8cKGUzmjxrUfSXo
g1thvi4ujoHqsz3304/t1kc2SNt6p+sL+MiPn8Mswk6cAcogFgDhdZPIpavQz12ciPbH5sG/+0IZ
1MJdON8brZ05I236Fc4omxDoOhrOP36S/5Osp5cOagr8IP/4lVeNYaltZQQYkRD+GgetUkzQ4grh
tDqgZ6L02tcCJGybuVKiDsuGnWgVT6LLvuvy3A5xx8LfKmry/2+SECKLe2w7jBHyxEQ95Zm/zZFf
mRqOHBNCfXwRJtjz5ztMdYpXDZ2VmdaIyDw5CJAP+ct1n8DEk4I9qrFWBsK5z6UIEX0wa7gVSAPO
QHWNBiKdCcoe8N+aYzdiThq9jdQDoFwvH6D9qO8xJy4F4vqqqk72Z+VHbMJjL4z4EJxHm3Qb1Rbl
hHhTAyGmr1v7SWKPMxAj2qYwN3DzSMf9Kk+RsdG6h2oCpMaki/eGWI66WVgJiwigCgZtndkp3qsH
NZOx/EXic4P/kdmGo473QvzWNA5aVlOBcUsI94gA9ZMvfZn7sE0C4QXmE7YJpOenPd306dsBAOkZ
jOBC8SfzjyASqlk1IkYpkraZg4Hy0FBP4GNWW84M+NGPG9gaCxzqMXb+cqcfCjLJY2lOzW0Wbne3
L6CMEA2Wm/b51X8NIf6oHTIMc5qTQ5s8MG6vBEatvUDkPO8pqYXXD2/p28/SbSKYrqhXartkdrP5
l3LFhJnueAovM66ZPB2PpHa6iMr+pFkiER6mVsIFTkd6ClcGXuN45gsUKR9uhmB1nwDnGyNYElMH
OHCBrlt4l3bW2Q3bw+aJcLI69hYJOa4MIf1M3sw6wax4GDF77K02BGSQMViDo/S/yPos0nfiTKMa
Vx2n0N+57ypqAb11EaqqTRN8t/1zxngxl4VDhy+jYz3/Z/DasUBcSaZgiVzVH1LJgYe7paD2Nabi
NsCyYGJnTlIff0471sEdAwsLcm7OvecqyFEk+u70os18liSzvBmB+hE0Qh3tVj12pllD1jWzM5na
vPwggQc6upTv7x7Okx9DC+vWWgCOI0WsJLaCDzFXDURuwjFkFxwH8odM5cgtGGKQC5I9yeyo7X3m
LD+3F8appgfUZ1hs2Yl1ouzIQiEGfW5Z1O7l5f0AF/YsVPf/oNA/bHHP4Har5Qqbt/ZcivLoq2wn
cxILeZPfBiPTkM2kBlZLLnyNwsrG+kjaIkXcewGKd4q7Q4uvJg8tJfYuCJBxGkbxYOZ1LkzTPzTO
l6b/jQ4szduWnoS/FcI9FhRX5kdbWeRPDW94VzKs0+m/xqnFSOnvV+buZo5nT+FgB3l7u/f7KJhc
v0Eln6Kt5i9xLAGJIcS/VPPkOJIoxYlDtbYWcxo7zZGFyiubeTyBCk/ia9wHxc+31nuWGy4yscQM
DIPLxOfMRqA3MBrUHOMiSdPLBt9jbnm//XO7mNYENLGz2LeFp8dwxvpT1Qe5TrTZh+eULCPPyAAF
c8DaY1PyxaqnSq3iKXBHsai3CECU3euSuTh57BF2WmobT+tSwUcWpgJLZYzyc+lmACI3fp+yvLN5
nO4wNJ6U7L43n14INn0NzA/rNxOfE9IO8BQZm/c3iMUgaM+uzlDEX0Jy0ArVIlS/19LYhW2hiykj
khHSbnJKJiOrERx9MYt9n/W5C43OTDNtiPKFktm7dvV3vSdfxbXn9bKYXEmRUhaWAzWJR1vWeKel
3681UwlIODakGGnELUPiVRaYKwmDlApMwlTs8zPpQ8ZDRu41tdj4+dIIAFClOvOKisg+n+NkFA1y
jr+BVj6bkMZlLIXIueb3WOy3+8wnkpnRit0xBHOukMdYcxNPKrwl4CQpulEvcNOJifhGUr+0mDz5
897hE8G9QZKOtQcLSQ3lDrg51+AabxT5Uzh/P8x2+Qf1zQCiLjAMicrs/BJHu43jY1BCcRQ+po6+
nVFtr418lsTiHzkEYgIIZkK5MFZ2dnZc6FGEL8n31AjgaP+M3cw3WT0WDDnhIIwRdJnA0E0qlJaU
wySx4aOsrRgJxitRA9ZQtQ5ps6DcxhexNpY3cGznRuNpY9yfzd2xVPraTv3VC1V032i2JSZVtn7F
ifP9ylVkZ50VZkX5cGvwLM6naCFi6tH6Lg5HQuPpNFvRr3zF9Vz5n3hgHoPJLe1CLL49G6UW8IdL
i+wT3IAU5QhrKHdRas0gJd29WPnvfW/pCtSVuY9I8iW/Ffv5EAEVcfrWlrlq++WfBGkG1asDwMez
Tpxnvcr82ThzguPPTd+0wXv42N/CDHfihUX2zPM1zIIAKc/fXUR8hlSR1Un4ZcBOgGimGFoZ/fbU
OjwgO9Rl9e7tPGKiZTigTCM18Vob/C1fMx+m6fOLUvIEMGZq7jA1zuj88wo91Knkoc1cPg1/58tT
TGnMcz+OVgIO5ATANC3FBWp9P8R22QLlM3sdAb3ItzFR3XvqOEZQPgNdnmpYQ81uFIci2ON922oY
IZuB54lh1R2NuAa/NpbuYR5IHhlrq10mwD/SHI8l2WhCxNYBJgX2U5h+uRmU6SrBqIeYJawWU8Jo
XO2smw4WRt7TSsBChQDGaHbh5qubfcxWkU3y3HV95qLMlqJX8KRm2K4HYhkGqDJ3cqdpQgOiemJB
QyzY+N3YE4NT4mMGEIgB+TdwVRQELLMow8Q/KWHLrRwAERZoTB0z4aBCG14ilMcQ4VND2MIYueXC
CEAgZx1nud8Sn5EGwdK5sqKWOQW/YS4x2LIEN62q9pt5iPwKZsEmYjRYnMWhKuWhLJEH9WGMhIi6
F+3Iox3rxOztTjOYFbqQp7qhcYCJH3Dw+8KKAnvLebCB1EWa6oyXK8xksxX2CSfI2bqSDGWg5INC
P/ghgcFVpuSW5cXfHoDAdltQI5WhWsy9+U+kV/L6eCS4etHSA72VZ/YGbR1RSEVwf7izElsMKg/D
bFMRZHfyCxS+/gh9HNOTB0O0ceNaF6iuxIW8MeKK8UQ02HLRH7zPEaI5PVSO5A/i2jUo+HXZNpO/
Cu8D4/1o0v6r4RJ67VJ7Kz/zCCHnwIPu95KLC4MuZ5yk5B0xbYwMRdOyqKokWFYQAWToTdt0KGOx
NlVP8Ynat74skixUZXRmCtVuOWW8th8gJwb5FeQ4eGvNyI3svoZnLlpk81h1xZuNk8MUbHBIOQ97
AzK0vsQK5UJM21W/ktDXiDJfyzbWiHqY3wAKjoPm76Xt1sGypcR6RAZ0Qlmf2DDfgViPvShoP/qs
TYz1B1pawa5V3axpKb1xX8QwN6LAcHB2FzTbhh93uSr0s/nx4PJnujheaL6gWb/dIhm5RdEKN7Dk
y5P9KXXO0Nf8jZEkEld0pV1veuCjdLJuPdjvu6dFJFb9UbKKJNK3Z4EYCKc8A+c6rfmYhU24csxe
r2XqsyWTRnX/VYU74LAuCkxVpIjW1NS/KZNDLJ6RwkYtbFPvQaoSPHMPlca4XjcK9GOi0XwKuw3r
1T8XDi5yDs994cf6vCKaLpYhbcnyTm3MbCQas4EY7FNvIla1r1QNs59Leo1/KwcYEr/zx6AnGnvZ
eb1NaUTfhYn+fh3BhFoB60SpqJzLcFGlc10xi9LNbxZkSDHjP2oI8w1xxgMlntEfOjUXKdc3hjho
jYHJqTYova/OK6P4d9O2PPnBjQ0hnq+jktNNQOcFndYn3jOYYtnoU5LSXht5RUGsge8qPgsvRXVo
iOeXNM1WEaknYVtSKY4wjWlLLwWn6OT5pOnPvroOOIq3sMKUu1OrIXWJ5sOv5nZ42yksMYBId87j
JqFeaZTTN7zraIHfwg2ev8QmmWeC8nrQAjiYjIlg3S/BXTQ/l9tGt4ndhgfPoc48BquTPIbuAIqq
j3MvJ16vp9vPXjrvblNcwh7dbLg8W+JbAcl0UzWF16etL3nOegVksrbXbiWounA2ikZbpiLknTPW
2wuKRgVeI7g43OimPMychIBBqQsVhzLkGOw1G0S4bK0nYyt0IHVO8PcYEA2L+HwKVo/EfvLF+aE2
izWoNk8E1V1Jin38jGp/YLWny9WVCnEqKlient5hlSOA/si7lDGUl3KLFvZMi5ryCqZKBvvmnfPI
wO4hHydPWyeb4uDRz2UnxulLVhE5JS37X21IhdTILyjeE4YgQOmlczqkVIsYP2rnRri+yr6JMW0A
AjxBKpozshPl/oQRhumaecHRwB1r3S40wBpjsbu/VTl8tEfRfsUlTCjzmLuq9bGrLYXvQHAXYSl6
IpAg82THIySt6xvGHYZH/yEMW6NM0Sa6jbOtOzfqLkxO7OlBZUVVVIQP/0lRK0fhbsC8yeMX66g9
7WYeEc5C9/qo+thZ3xqYshrGs/4/5l8/0PCWRNLOr2Rz0DM9uwmwQPzSTEuUKKbESFMbyGn3LSsk
+t0kjHVBm3SpvqesgsNCHxZAynEdknYj6JdUA73+XurSBDtqBlUEOTGXBAJ9PjyWwuW4gWCWpBw6
ZVG9DPTDxL+DPXkz0jasUx6n0gvK/3bZcoB7MQyydfP2ZdwqWa07qZ9wefwRuLBsYljEUfglbmpp
/LvSQBGuC6sli4um5x7bMUU1b4PPL9bpPDLTQ4BGzEwpQSSp9AcbXq4A84GM9O7UXjBwU0qG6XYK
c66CqqPSPf1JHsczVlHySD7DuLEjRk7mawsZt5x5xulJ6wce+WLaAtNz47yP/D9gi3ajpd2AzzaD
ZNcRKi2THQBV29Qz7KHAlu3Stg5d2807N3o7fyFqKKHKpdhEU+oPtByzGDCzJ/jV0urXJ7diKPUi
r57yCXLKt8ILD45D47lJNYQZwoG1GJaabNlPF6gm6vwoKrWoSuipVKn17Ud/WT/L/pNIKeu1dW8L
BRdmfOlELuzxXrHgaXNtag1YoKbD8jSLJw6nxM6sqc8QMabUTGq3TWikEEJhdgDjdfkCH3kM1ls9
JW629laoICV8Apsz6GXROABI0PnI3pD/+/z7DuFCd/FxxN7nOSEfTcdQFeZ4f9F5V2sOG5XiV6fm
MWSAKP+oFTap0w+kJjZyaxYPW7/PlIv9DJK56YJYnPrxJItKFtJ75xYRpjcAaw8MlK+3NcxEmwbj
Os4zf1KfelsfXDdj92ZevRfxMltNcFeFYWBXGGtZdwPGDNNH7BJgEpQ7Kq3HyqOq882Lw6l1t6a/
UlYAM869mkbolk3AE4f/9pLZLZv+uAfqYjVp8fBzy5rfsJ+Ea6CtsJVjXjbaKRSDXXH0zuLWy4e+
E1a5uC11C3xokjZ3xrc00INXUy0ohL5ZDukwq1Ltzw0Fl6EzBM7KokYwXzNJR1UfUWsEmpD8FkOd
HEDTJDHtggBGoGMy2MYX+LRC4IslThnQXIzSiAnPCpMEt+nKen4IxYHXPcY/asl0YNyZoVV+UrFM
pNQ6YRSFM4FJRYJsGR9PN1V06HDmALkzY7m9ZVHQxVt9kkqv7vr5xiOXb9AyFaw8OHpPVSHp1Uwu
ACJGly7IJn2kgh+iflgr4IbCL0FzgowMxmIY0+DNYF0ySRgoY9N19XrJZukEV9Z5gwdo8YX0Q0oH
4ZPWATOORW5GLjlA6jCl9VesOHArxUSIoQonBcpkX8a+gtDAynuLRSVgQS7Yl/lhLRfOFT5c7c+G
XXbMKRS2WLMVR0OPorvnUhpEaZkiG0Te4+sf85Y/OZBp0A2qjTbnhD2U+huhFeijMNcV/dcT7qpo
5iW/cKi9u/o7AOlk0Np620sl0bYOUvdytStz00tFRftvlAOa99wUDcpks1zwFVVHlbuD+L0f2VIf
9zIvoq1B79r+y58C50kuUxwIlZhN9haE8Y77ey4m3UoOtMflccfmN7KRJwAmJWWCj15GWnK9JKZ7
j6pWNM9ErD5CSwXQ7d9Cb8srT+DIMckIaVkord2ubsw1+v1Dzjh2a+YlwXYxV2c5GXWvQ+Hmu2gE
LeLKHQ5UWencqE2g180REVcfkaarveZw9df9Fz4OjGGGecKhFZ++PBkI21xrGfUl18b7lP9eVS2d
kEm+GuOGjWZGZCd6nF3pBpFp5kyuKJU+Q4XbKZ2jxzwrlgcA8gLdpeFdZfY0RNblyHDmYBJomVx3
D2U4WJ0P4dqNHR0xWtNPrex3Aq/ujo53OZD4yHmDmMX98nnAy8LgRIbLT8a09tiMAH7fcHHh246M
zqlWY/dCAPb0+BYc+2CS5q4uAknxED1KbTjUtVD7oJGGmmNlnkp+gVVwJKMRXY2pFQ2QYsuw4I3J
tJ41ucDTOSed06/OXHwXvbIVzTa463CMy27W0hfKd4KDPphoa34+ea6cO8MP9dNHIILZMY4V3sFE
QR2VPUPy7OgNKCXpAKH4SXv+NhV42dsCGFu5d0lmlitKO0o25GeU3tFZ0+5P3bsIT6DeRaTGyL/3
c5DgSuxZDBLKSlL1zbLJK8fQ0sjcPHUPtgUZTkUCnz8Fe928hxApT7vS3FwXTXSSuk2IyVGF8IF3
JtUvT9DPAodcjhdvDiFVTeWua66EHFOcUKPqpvU6L4XFB5aLQueay6eqi4DEw3TmBCBxwu15hemp
DLAru3r1GW5dPkLLKDjaKUZRGu/oKvyYsLw51jokvacGtAvzeq0ceKuv0LLEVfPxPYmj+DbJk8ad
+GNxF07mbXllHhukPomkSdGoHqHI+sjYeD2teD9WaP57g18A5ROTG1CWIuHDJ/z0sS3Vnlo+yivf
GmHtkrlhMi5uxL10UPaQkJ4pfiRHMCHF4glF5biARwelWBEO5QHpjY/z1fxxT5U7n2uwnGGrYzHH
eIO8hfmfHXX30DnpnkrUwCihxqUkKB097Puxh8aDAS4dRmOQ3GQT1C1MnHp/ueK6DjIYJ4dtkITq
1cqcDKSGYO8ihUJ6MLQnykcKytr994DHkGVL/fSEEISZBnAK4/ZR7RxKIJ79ysk7lCA+IxVD0VEF
Lm8X2mBA4voPeqaqN6WvVAcZ8PywDtGK3o0tsRBCuiiP0IA+5ZXzb9zRA9TyWN7YW7PdKym21iLT
bw2pHnun6IGtByXnXbca1jukrcLcN3IwPwhosXtjsV1MVsvbqHImKmqVS7BVKtLxLPmzVN+cbNiX
N4KBe2aJjkBdcfjwkBrtVVYv0ORjXs5JbgTAsWnzh/p6iAnEfFf+1PzP5WbDSdyPFxs11x8PUMus
FNLjqr441/XsI7B5MRZgX/fuDuGX3UCtBVWHu3x9GmFg4EaomNq+vlUp1ttzvC82mww7j/6p9/tE
LJeuOh2ofYnMRgFbmliQtdXFvIEASnw5X8R8y+B/u6riLR85zNGqK7U074UDIVycQSLRV/qq8y3d
lY/rqLjGDzAyMisPKck7zKztSoOZgz3a4LUe0KUdvrkEAIHvvPgGHZDnTfIQKK5ZTo2Is5ceNCty
dvykw1lgTE6MoqaECcFrMxNQeYBQvAtKSLE+26z/C2Br9vMeOXenpSm96a0TopDF0LulS95SlnBq
Yw76gHv1XdFuHrmzu8Bxjv++2qz6d03AqCnWqHxLBQcjLREemktfbxbiY0kniG5wKWO7WYIdfEW9
RCA8IlF3a4OFS+cxIksvTik4FNdKjYKPg9V+/C2lmrzptF3mmHWQ9InXc7fKHzNFd/P4h1J9gl6i
y7KV8WBfsaBaI3/wgXFFtFKuZoQ7xI60GGlH0yAKCaAm+s9jhSvHZZHnK+MqaewcdkfC4itPmpzj
gjumCobRxs+pw8lYvgnF8ETx9RpTK1Nj0VVHHCOFd11YiqSGz9eS1zly6k6kzJY2KfNhzInnrvtZ
nz4e+mRrG0uYtJCX62mc+iNnVaCSbk6HZfc1K3Fj8RXyJ+s8p5FqJwIGP0E1MFIs8Yzv1wPm7Gkr
/ffjioyHIPxDndti2fOaJRtJfjNJ4A6gWMrJ1MKBLJCkhLKZiy2LrR0j0XTPT/c0gS88QDLCsXJu
Jcbw+4vBZeijQWAblqjYQ+vrUhtUOczXbQz6GfkiQrU16R/Ldsq15Cg8IOItqu8ZoTyd7xmUhwjy
8bd0OWiW8XUw4/kElthg3o0qqicuVFnaBI0dnF8dlDsldibsaf/G4RLwd4Lyc+z06MF2/dKatOyo
529YxNx2+HOhPzm6iIr+Si4OoM28n3Yf20YWgpHmCGipusiPjdEx0BJUmUETuHDqTxJbfwcQ/P1S
Q6gIAjl45ZuE0NbUBlZeqyjxTBV7X1Z2RdprUQV+cdZOOFaM7ezbH0XYskTc0xqgBZRhuxJ8Lz1u
Iz1Z1r7iOZGpUSOY3t+JUHfc1EU3O7mf695wGSfmTq5FELPzRpsBDKb7IC6jtprCjHXaQF/S+fO/
33EIE5Y3OwrixLBDpftG0Yvdm2wV6aUD3btq6mXxBuE2RsGACeUvTTEWvjB/zWrVmW8RcTHty0FU
G2UYiV3ii5Wvgq1hYoImyWmnk/w8ycmH1gCSD/aBklGZyqRv55jQWI9D7KQW7dpJdBYJWbZS7nn0
qTyCOrUyRlX3J1VYzEdKDfDN6EGe/4cBqBvh3dMCmDE7/VYp+upnK+UUeXM3sV8KXQAmBIsmcCtw
xzB4aEkwekqC0hR5/1Hti8SwW4sKSOp2USxeTS8l5v4RVAV+UW+7NKcmPRgQYnNmBt5FGE31oadX
Ojk2H4uNPsb8VmnsTBD8wxfrvXVTATDcyg8G4Y4RU8Zk4sS0IfDWPT5AsfYLvlLEAQhWjZvQT05s
yMX+kBkq+bHdN/9O5bV/gLRbU3+rRJEbGp0kNwtvl/7lzSb6u957VYaV1zDk5hSYsKoUduBnVRBk
tM7b73LqXltC2oxTI9VTpDOhTCHsD8MjLME84cLqIXLK8chpD4hvXegRSmsgwY/9QnnJoUJhzSIx
ra8Lt138BFTFxwzWwTXWZcasRjiDnBu6te0tXgUGbRM/Nvez3bhcvtDUqAQqfvfgELZsupz6I+nW
XNYUH9SbXoa9HSNDekr/FlNpwoOQgiGykc/TKJmiYY1w9u4S49kIlp0kYlDLrG9g1ekNjijlYde8
py3GIQ4kkhPGJ5LSKcLMTlzLdTRBh81QI1nv3jBdiSEjse/0qbb2YDp0nl9UGg6g3Nzco8JxDe/G
wss5rOPEwfGl8ydAQbsV5hU9gO4m06zN7zGXFm/EIvxSO55Jk4i3DUei+8owUrFZ5aJC/7BGrP6+
OHTc7qqNZrGYWnh4EVygaf2g49qDP0dNF0GRRjehWFWoV1qVF3Alhib7Yp1wID3g2jXhPzNxT5jN
+52HrE5Dv5/52OuPAbziyG0CmBLN7QSncgq1zZdASlLisHbr7lx+KbBbVkHl/rEZDFW26NE8HMGU
GabTtf0dWZNIa2RxzRJzuKZCZO9Ch4rt9W35Jq/dUH7yhzNksPcr+Uup+cYb+o7IpWEvqzDdfm5h
TD7FVofLTp/Kp23FJfuic6WUxQSIqiilX0EPyB7GfXablmdDzatiIoJa8Fh9N+xd0ZN3BzH13sxQ
XRnVnvNYeWPVg2Vx78/bKvClvewXaG6k/MPnlaPvsQa+Gm7p+PE4+SO+KhV+lOLBBVyau1A/Yh1m
5HlyMyWZ5gsKtjWXmiOgL9xGtrdJkGynYvqrZh7L/pbh6E56uaGIkrV1stqUh9xqEN/k9So4gJih
T3TS5nJfH29dQ+buTkOehE4WInXqh6A2VEBkMmWLSEU6Zbc5YtCgi6bA9KgFwplowk4oc0bfcedq
WvMCtlMebaOy0jueGfZZOBa5ZIWtwWBuSFDCTiwv0X4/ZzHywGp6qILsztyEMkQ2o2JhHd9MWkIS
lKLzVwo9UR3IOoWSAVB5RRze80ZDVEfkMgwyuAuYr7r7b3HObFbEwynPuOkWzCL4PIFBfuBy4lnD
8GjuhK13fiGKaAWQB8nnB2+0n+iHE56YLp4I5MDz3n31Epcd2/rK7GchgcUWIGSj15T4WGHgcQmw
VhWQ3Wk+grenXch3uZjIWJGK9Jir3mrPjWTxcisd7cKHpm56TqCeJA8xX2FrxN0ZXAtjNAeepxkJ
a7n9GW7gHqLZcwp6HWz2RxwZLxdqdOh5jkUERXZ6YXyFrZ+MI4Ja7/rZCM8ILSip+ocwzYaOSGW+
yu5o7Slo2PHTH1+nYCJhBTCXoshWCcqh8R0T7UkHdOdm3Q5hkhX6+vEFzpOFxsyFAG/Ejg/6HbaY
do3IBcw6kfdCSLjMv0Gzi4R6oU54/Fkub7xl2Lk3GDjtfljL1KXDWdTJNj9zsJrVFAPjaMncLmMB
ZoR5a4EOQSwcWXxElNN3ecMwteO2aAgNki7Aw/neAic5R+gXDGAifMaqnNqCdGBk/ZHRO1eefIlV
lcCGSqM08jJsbzTWwdWFhzz0aAG6pHVRi9IhagWQsHesb+KDHmoZj7lhAaQ+7cccGZTU4HUQjrXK
PvRNIFSJGOWOKT4BPIQlQN4k7El5lhe9ktHq480aLAuJmUb7RjEezFy9zl8KUrHjIhVVIvDJYtIn
YruU/WTxqodIapXE3vKkDtG5M/D77QnAzzOlzPpqVzxeJIIrANXYY4ufhW2tyG5b1V7lrPRSkPFM
EjXDSBskcC+vrSy9dmDb+z8hFSo43PPY7cd7e3CsMe0FKqyeCOjrhp2+hLnNhQdC+3/NdVqHQ6SF
Id5pyTnI3AS1upmMXDP4lrPqlXgN8yRkVw5G73ufMQRs/FjkKQGIxOP03vqduZY2eeljUdDe0W8T
IyOZEiX4202pu61u4hz6ipcuwZgfFZXEsbcBO4QxI1G4IuMg3cZCSE2NUc4Sv/KhpCgzuJTvzM9B
D7Bh8Uq8YZ7iUzrXMq2rH4lJqLSx/awnXvGM2xdA8+TMMtzpzpvWaD5TSAfEtohYgTKbNvgy8+Eu
Dv2+aytGj1eVUxeWwrYBw6pHDSRgMPWcxJkSQkNa8lObaipj6Adm9zPZoCrP7Us3LzGM645cWZYi
QbYqfH/sUknwDHvM64EByelnzGG7VGztgGgjtPI07yDhzn35PP4xaK8ZI7yTwUkPiWdzcEXJyj06
bUHli95xyRG2GENqxqOuUWGGyk9KlxEkzzE52xG9rl1meow/1Tldsw57WHsY+pDRwNsltZaJQufo
1l+lWBlXH8NzTu6jbttPYvO9sITQDvRl6jDuIeQU0+A/xXpE7UD9q97n2HyvlITrqCP1CD0w9do0
+apisTVwSmj8QNYKhYiPNRckv6/Bz7VozQTxH6Wk+pETmt0XLvAYNlKk07Ms4qp3E3SgnOWpot00
vQAhvVGWD0qt3YNPH9iLX67NR+Wg4NXp8JgPnBMJkEyYwrNTIhcj2bWquSGNcIisCd/UZXteXx3W
W8ZUNVfXKsZC6iE/s62TC39GyvDpxH5rwauuTLCgrRC4bDX/7JWThWYqKXMlEF725ziOEP4GF6Bb
3vF4wAn0gERwqZlryTwpiiD+zXwlsmv8IHA8S19EJrfdTVDWZpEaDavcza/MDOwp7ZxqseoBsvTM
eghgugwll6jzzzv7yvrlbw7Kwce35SWa/+cv4rzO70Vkoo6Mo75W2k8eChGEPZYDXDDrPRI4xEAx
KQHsJj0+JVj9VzvqJ8x5qHaSQDnPWCai+HUpMnSXEtI1KBimnvDuoz14i9GferQw9alrRuQvMunp
iYsg4xeMv3jtIJk5NCbSXBXZRq44W119eNKfDqU2TYl5cEJLJAueGrREMxAmrKEX6Nb09OmEsPVk
OQeUGDTKNlIU7rWYqsBZ3oEFSD2b/JsOZ/zr1yGjPXbZx4re3sXwqQQZNiwl3QarGA/WMN53VNdV
UmrY1pJuGmBRP606BUVjpiVsNVJ/Y0ILrZzk0Cwrl4aYzok8VEHR3KXL1AJioOBtQuBdCfAIH2m5
Rv7yeLP7CPcwfC78YF/b7J0WvtTFGbvDtP/N62z56QW43++7XhmrtXg4goPBW0tOtBuryVV8n0A6
LxcYwDJnIfrXoeqDYpbP+RJE6M0aeQJWzp2mLJ8s3KkdcqEpxtdj00trDRi8dRjZ8iyBZyTZzaOq
JDYRUIMtam6Zt3nVppJlFan202mO340h+jcV4A2mMp/xcDnHcw2AP1Y0+otEKV721hDEFYFxaFVB
fditoviOpdR5nPBDcyxfgw2uHLqh2vNzGuG7IYTip6VDUsS+PJPYncYFtgwg5/U3i73yYzSLQL0I
6TzBVdsoSOvJOKI6qRt4ak17dgkRxOl7/zbHlY2aQJpREXdimWEt6Kdm23iOuM3jCM+OS4eZKobA
iUZ++3tOrMcUudl5bbRPbFrG9q4g7i0kyIsdaaFVfdOCW9pyBS9hf2H8TjRZ4eD304SuJrTcNv15
w1IgA5U8hcWhTHCt1sEEJmeRLWumHq+c3HRDDtVa8gqtrJYpIsakYy1syncG45ofLhB0Zhvg+Kxu
PbEYaCiJF4lkcuDPIAWT4VmJOU9bqkoL7oPTU0lXO3swfwwL/Ssx9Wh42REpBrBCVG5RvVolZjD3
tXimjjQil3c7Rp8u2PlNebwoXpVCMk1IoqmlZpkMGcgvmJE48IXDix9t1IzAFi9E9utvn5Glal3U
Di9RxiQsLEg5bs0BVwOM9cASFfiN6v+64dVUZEf4noqBOwBiG5vrf4rlR7mvGSbPj4rYNSN5/v3o
Xjd2gc3/jnb60IEHICpmHGujVHacCJnPDfmjJujem+qEOnsb1KsrvA83PzhwYUlTr1zIejuxeYYt
+DOSH1oytfnRB5raVa1KFfy7TYQGVL8zmMMeDwsFuxdbaDPRLIMtfJcFtPEABys6e+pqjrSPzK8X
swYx5LFpeoqPIiWF0J7UKZypqR1gKbnIyXHuetYBssYEpZtg+HcUNmtnUEsSqbw2xDTOkwkXhXs3
8HiIp1uDFfPhwTcnCpmDAry8llDNPfLrAWmQaGyTVW7pb09p+3fbYP9zkMBSHbUicrIoLEFDc+YD
4c5aVnQWf++jpdWCrgpMv5d78jEHB2ONFxUX1MBu5Ew3IzBK9/ko+rcn90VFBZ91BGStPUMyQGTQ
r6SFTgVIZTfgBSJUeU6Y8AxvISHg+/aYtKRZbYgWcWusb79RtlHjIOFIjQJU6f5+qzSI5tFpMV63
zVWeOXZXZ1eiFz9z+CDc+MNVIoXSLkt/UgRw7gekoDm5ExqJT4rm/zQ/haFo6ub47SnHWvnxncdk
WfCUP2QDkh3m17HAGjWjtWSJOF/smDl2O3G1V22OPwVLivUM6DAjb35MQiS+bPbUBxDJc/2Ir6zq
kz59YLWa1NLovRS+gWBvC0Up/7R7nvrTOgp4wnel94YVjZXB77Ydc9Ddv7BAl6l0LayfV6DmMPqC
roAdeqSSPM5iVxG+xvOEEoQ0d/bL6xFQhtFHg6sgYPezYiTNDWy/obW5cTCxLKvKZtSoIjhWsgkb
HeeFnH9QlHH2d86i5gjGd7trncAQgfF3/VH6+NbmK62/ECDPEXXpDoSltmAFkikfteaqYPbM8SF4
HoRRSCFPeKW5QPcHL0etVAXuyPBY/n1eujf8whvCx2JbzScTbbprGVq9pl7/TksSbKJ97Wg7KoN8
c7vDBwk/Djjjs9LxVySSix1Nh3LajupWFmJMrS6Wy+xr4Zk+T8CJZG8fjxITqx0Eb45cfOVl2Vci
skNRQ149AiOPzGa82fXo4GAsqJ7fMvoMeStrtEJarzGabwVtjHMUqzz/rdplbKRX3DxisRkShsg7
qJ41nb9ekFrj6v6hTTAU+lydXoh9niejTm4t6wQ0t603PLvT3VPKkB/PVl58yqYAewGLG/U2Oe2Q
FwRX6LGzEOBtFi2YWwiSYhixG0+OJnDnTlcJxSDQ/GxB+0e6kLAsATx1ONSC0MJyrENpvIgqki7C
ORK06gxBG2hC/B+Tu5Vpajgrmb84p4Clon/TeuesnutApGfZs9X5+9VnMAGppFD6bHK3O8IrnO4/
UV4Mk1acRhUz5DzORMfcueT2YFb65AG2IKpNBl6Rrkf8zPswVQCvd+eA3XhhQg7eT0iFL8wLSx6w
ABHXq57pFX83ja3OhSYf8C3Qlsk08NJQl08CdGItrXGiXLf6y1+NAisab7La2shL/kGbAFuNUopP
0jVsAvK8NZnDpWl3S9q158Ue6jwa+esptoXyCrFc2i4qnUDXm86cpXf2syi0ewOrTgR2m9Ym7Nwd
6bqkIyLAoMXPgMkKlM7mSQNKQk7U76r0T/zaNUOw6GayNhYikejQsfLnF/53FlO0p44q+rqII9ty
hTRfMZnFEfBs1nnwITlFYs8qIQHRa5Xt+XHbYu5/HIGfL0W8VutAeLmKQTQ85uUjf5ERUrMCsULz
PBffPZZrrBEyStul6ry5bGYgdz/PwW4p2ldXFyKS4iQ9A9hSYHf+LBWTkWFm3MzRv1Fw7abKFK0q
ERVQT1chISNA7O7sAe9e+fRPngk/W/N/9K6WRwMIkDi6eNARWflGM/QhhBysxRt83WHGrKtjFAbH
8wyXO01pCo3hitpnhKGZuQgdxt3/wuVvcMzYxeoHkXs40BVy3a7MT4gLrSiTmZ56z5nDHd0r72RV
6cPz6j8tAJEUOmaj/7UWGPauIpjgfilaIaPa1rVZS00WVAlj7NX7GEkcJjwhftgXEFCVRFAxwb0W
hfF44Lp+rEf46vEnFQTZHwJeUlTI2PTwCzX5kRreAUtxSw4JBrERmnF6l80Y4i+nOQ3OxgKz1yQ7
eQLgy81SRjVp1wZOTD4N2HEbH8RGj0rjJ8JVGtqoNjzYpFWepssT1dotaX/EaHNm4aYm2rDSoUar
etxKoXM8xbawei8dexkz0ag05U9RbP1QhnHDXK50OAF8EUCzkETRf+4y3NyjgGSLy6jHTtwJ4mx6
DmK/WzVsWzrD1QMup7C1UL5aoBc1R+8GN/zBDx1wmjb160GWTatIYfAnbuhceJtR/Tz1z2reba6t
f7Nr8Sn/VTEHo0uoENXs0YRkM/ju9qqsTZp7rVztxwGD2GFG7ds8hZM7vcsaGP3SLB6BRslFbK7S
YMLAQqIr73bZp/axVqsSSPVvAzli6DUFqQeI+xNaHcQrFaEmhfM5I99woqGDru04/ptXyb9EGXvX
kr2ElGWeYP5Hjfs8JrZIWf4MboHCeegiRCcdjx4jrmJSC9ed7pZoN97JkT1xqtQ1IcUN2gCHcdT2
gYdXkLbeJ/8Am0Rb11bzqyfjy1QzvQjLlx931ujSCeQZgZ7wTEbz3StkddeNfdVO1ajwh7uEraHG
0DgsPSNLHSzB+L0S37chCEew33I1jKt3hZUklUOoG5PG0135z0LgxCAJ6VccNTQea66YBeTkodor
ST14hF1GylLCmSE+bva5w/2+cuOkMix5Jxyg5z+XmH2MHgHIVUKoIqdwf0Ld0vgg8M/dZkLC2Sva
IOr6lVPvAz9c6xGVX/oLHq1QTJ7kq8ahTnCz2H++7dZ8T0Q7uJt9mpjv3o3WQYiSQrqoqrQG93qd
Kqk+HAgxYF0xBGbaJO/f+GbOinOMtGFoabvCE52Ogde7ph2FNGcxZH9vnOtYbkWLXtIbS2wavjLa
jXmYUdB/ZonvoNNHti38EhctjhraZpZyydiwD0GPY7JT3f8QItXmx2+FfxYbOkIEl9rLqNYBiUty
k2xBuurFqxo6FQggBVF2JlpmN0qq4+GBIfB6NGtuA4CrZRwOVhMmJ5T1Zwql4yUYqtAjgdUULOwa
as59u5MnvPQxUgCFhmPTbJVGBLTYrARwAaySgmdXvY6YStOGXTCNdXTXbRwD7SvlYLLCYWBzmyAX
eDUACnczrzI5TkeCyRaUROflUyKwhZ2vsbmgmsIrU0c9K0tA+9xhyyq83OdvO985A1npzuns6CJZ
ND3n9uY+jwRXfVuBSn8ANigC7htWkZJzpJvPUtylxi8byexRbSzPqtRv8AbmSMiNQcxpY1M/ryVP
vIagSJROSNTjRQB2xMqxRmULK0wN+DE70+n/If+JOiLH4IhWE803PoUc3vETZoef/dluSmj4DKYW
IhEkwOuxCrjRccOC32TF3WEWdM6bqRxZCIU3EdhSC1+aG7/K8DynONPNxq1jhTMu93JZwTYlm8us
iZaeLvynsbDD25wNUG18jk9Q1uh9axecfm4Cs8yL+HKFehTPrckDxbScIv8lb2d9eW0RRual45i5
FHW1ayUu8Cblz8c8TG6520LyAdJGLuSZ32/jaYZ1PC3ajyUu/VWTGklVp+hLgBJu3m3rgQkWJoa1
Vf+T2WbQjl+RoQXBctU5bSVu/o69QUaaVkPhaBqmvUJ5RYNTN2CLF03daa7uLohCjYtOGAsIGSz9
zURKvgDSBr7szWrEWpdRJZ8BBG9eIiLEuFpviBpojg+lQx/7qAmZrcceSMH+ezbX5DH8txFY7Fwq
210RJAAiwVxfnZS4Q6P/Aih1dZYrPDiJI1DhDD0Qah7jsAFleUI/PNYFEe8n+OfmntEG8uEOnhX/
HgzIRY3CIgGMuuPlIttY8jVd5O1Qe7iHxAPTM0w2qiLCnYluzqZRjozB2MzWPBOjyhG+dk/187PI
evIokylFQ80WrMnr5xQGM9lNhtS8Qkn6Jt786zEMWRQ3OfoW24ndFdOH0E4yW+MR6zdY10mkW5Ss
731yO+fxWBk+XS0nfzxrAne9JZ1Cg3gT4LOELWxaiUO3e05sktUX1SPr890m5Li1GjFXCX4v2TRV
whd3qEsZFzAqxoZhuYa3twG2aJ9keCNvg6bKlLbVIpWQv3ioFfvoOdqeDjJkzwbUWzr+iC0TDU3r
IvM0UlP+ays2BJYSHbEKIFiz6SRKGitSyqOa1sEvq6B1AeofHwWzHOR/O0C/vLvR+Rn3G/ahN85v
RcjtKBmfCem50/sUj3gXpxnmUp+YVdNJ0jZMQZK5eHFOgopbU6vXRNCsSgT42bwU0UpOwDVJEOrC
dHKwZltCck7opl72uZ9GqRF2zwO+RgrExiqe8kJJ3v+1wjtU0q1oQKMUYnoOlkyGpNXK992XkZVm
dLt1oPDQ9AE/l+VDxA5kwsFM2AxuEJxzDIE+1FxpEuT9SWscDtft4yuTuhJUz5VoIx6/Ufl6t2b9
Yc0/omqOIsv981brIl96iZ1gZipkWAqCqYA4f3gHAt5EOoaT2sIFvPL+DlOTXl4jwu3cTUddMSlX
hnOCDnPYoAv8BgL592A7X55ydQrNKfhGSirah/yE5/zcCJq3ZQ0pAgo98G86dreYEwZiYkYhiiSC
0lcemMCIkln/yJ6boINpdupZ5AeIE3HqU8r6t49IbGSNUZj0TEtq0KR/eOCAFClizKu9zAT8uxg3
27OVRLT4tFFx9QzArnH/9Bqfb4PjDEj5+LMIJfar6mm0C0kxBS9JoBj5rec/mQDOrfL20bhWSu+Y
UVALvs/F3ZmMuapgAqm1kHculbfM1Ji/1fpsMdh5X/VaigKqemlVAa59t/kJoIjkKM19/ZEfV+WT
+CcABl0TGi8RsIFUpHMeBPpR9gdwQt1UXafhT1Tfk1lETBNrR2LzPJwH3Pu7HAXfOf4FDu/jeQsj
MHknX4PhJU24AuBy7yP8mE+5g2UGuWGQC0F9kR1JZsf49NWNdxNr7y163ZMKW4P13ytbBMGC+kiS
DeP1rttBidyVdSJYMKFQpPsEGF3nolBLINvOygPdAGTS3DvUDmxjgvw0xOzSkEMNRlgi4DfasUhQ
rfQARRkiysx2BhvPEpdMkWfGj4qZhhg5baAUXoerwq/JPvy6PmRhK9c0qnmCNJg1VM25W1VJetqi
gPzfcuvB0KE/NnkCQ0vxEYSmZ2B8OEHYgJGnrrEKRRmhgAKJEGCusNsHXuDEsEvI8M9IqkoXpeRO
+sxNTGHDF6gENpbZsa0ok0EiVTI4P1eQllWzG3DSawIP2VgRO7iuXwrFqtXOCgzGYpJL5k7XJN1B
7uXaqo+BkR7Qg/VBf4+PscOM0GWn5ENnnuJfXbw/2174oTIQrfA+ikpDWDSceQCD9/+vvvk0775z
OtVkVLmXG/DPIs4bkW3sz8+J3gnAnaBqMF10C1MB8JbbNGNMVOf9LFMFq6SGdIZbpdW0twI3rxsM
dFLmXYh0nqmoll0beWVKKGPVyzb+k5o3f9ZMscUZl/4BOWoj8LqUdskJ8tRofe/fZxIW68dHrSl2
a+1WI5jnCZqhygMtSbunSolbK60U/tii6mNXsI2MRCg5CRcOHoUl9CBBe+22KtKXdTYkhvlzBMmH
Rmps4hd4v3iwIewcSNPa5zernLepklBn3jDFEvfkdxHtuDLCuebNs9YJUA96ALKSZFqx9IPdPaoc
GeDAV4JeojuHrHQIs+C+ktImFNOiqsv1/aZkAYT3xgCNW/NfHAt97/fMU/RTZJ/Fzr6afUS55+xV
bQHvK7t7rJ5Rbq26zU3P7QdZFVB0N8aC3/a3Gh3yeSqhsQqsPvQzC866NJcEWygzi7UF99W3kwcQ
O/5E4xnkb4wTsJlxmVzixSV3g0WK3ik3HZNScVvVAWrdyAuoMNYJweTWuIUkkXDwkiaEtEUHboGu
hmtqIme08UK7N8j1driIyi/+T4wRCS6s4Pg9wU6RHkG2rFIMIqtvTVLLwc7hDlqD1W0zm5WNhuYg
s5PwinqkSjdYoZbTCkqHmd1x4BJ7yXHg+rjOQMU8RSfND5+YHZFauZ0DEKk0FE4E4Zd1KggHO7PT
CrrfDQizBw4uVWXGQPMS5BLnryl2Q9CG5aVeVcozBVPw8SUeOmwpLxPzDc3mJl8AO4t1XgI/O8AP
qgl4EOz/ysly81Mqcy17vX7bcLb6TMjFODlQeJWzwgpfEXfeZXSoNMukWuwsXVdQfzdi2HXpBEyZ
3/cHeFaVj9PBBBxL3UuLUXRcNpf83ia8FBiuphdHZfWEXNyxeyT7RB5YwRwGyy5nPlnQhrn1EZEf
lCbwI2/5i8Gf8NLBMp2W0hEgNcXj9K+4nXJ//G1PtS7z06bk/BMjAUyRuR+pN5xxie8ODfvBnerk
2YAJCXEGDF5EEgwU3BRBogcnX2LAG7dKLG7/ZJAUzkQZZduS1DQhEKSJ+dqKtYE+ZuskyNXoLIMH
v/PnlsB0tB2/Gdi86At1KKutn+M5rE0DYSjLh40AK7QE+lBccRQaJjqTx9ikh9T2ikoHFTb2Czhl
1Yx8v8DE7agem938vdlA5/Esw/epJ/0aSsCyJD/nWluTC/aNUPZvmDLevjWfvEZzhM05IkF4E85m
icHkfRVTNQKcMyqR1/G+EH5c3DGPHzBZraGS0Jqsa8O5N67A2VAzcGnZ1OAXMSalvvCv6weAZZHe
YuldwBuYC07swNJ6G9yfLSKEIFQpOAPcOilcTc3ejF5CzfhybZpjOMjnOiiErAQRxYHjhKBo+IXP
dYQnX4BZu4P4LoMBzowQVOaAa4t8sGSLd1pAQaC6vkx2bYshku//gdF4B6ZlH2m6QqLzC3UvYh/h
8vGzvgLobeFHOMvIk2Oqu9Ms7ifEHmjcOhu5ivsUh0BEywN2kGFpShQwhqVDZXuP53fvWpEH3i98
0WvDWcpWoGtX75G5eBRqYehCbonUD9yWyxC0J8EYkNtf7IeUraStnAZ2GZC27GM4Z3CUz1QpYkiN
uF4gpS9oF7W6vqw98I7wKq1y0sJMDWx3OhZBYlJyjNkhsuUhK7uLhkSuFs8kBtp0optwKyERm4ib
1FEVe+jQzs09/JkW5Nij0fhpECKCU5djTlPdj3+AzfJ+TmtBOHuaq6xQIooRBMDUBooZTpMCiIVA
sfJVCh0ZY5zmHIUsoMvlng7XxpyLb2UBsWnAsPrV1De/Qls+PIigjrc+v9zGskCVRU4SjDGU1WdZ
b4BHmMUEutftVdBXEveRklzNsg5c+buNFP1yThoIZkop+QM71f06Mg/iTkKmZmJVL8lVL6qu8oni
/APxe/WmfYRK9WDwL5GAS5/MonVejGZGcHWOwKHhqzk0yOF8xFxuqg/6eU1isgTghyHtONT1kj7x
6WZsCQwnJXV12vhr3EfjKs1tAP2/NYHbkiG+xPJAlueyfWcooom3PBUFhfCO9TB3T2I5RBbLtlLL
mDWT3XL+Yr/53FC2cmXhg7K3r2EekPoci9eFfEOTP8DaoH5doM1I0ImxqPWblWMuUYPuF1FIkNy6
N7hy6B8myUfibHaF+PTEDQzKbaVBHNwFwgabeeiLR7ZALoK60qHCQOBBaNgfwM/FpAvasU/fNvrL
CAP37FmfhMHW3uYqA0XZTM/MG94no4D+mYmeLBzZ4PlD3PT24cVYxJS2bG+S2z7txWA0WqGu/Uvg
eCKR9P0Eo0oQGsJ+VvABIoXLeDVGS1foFxiDsuB+KISnzVZ46VqwaIug06GcTn6InV0TfX4ThdjI
6KjvoBCxOI80xaCkd4/jKKYTuxhqUYvsC2Hcj4t/aZR1KUxhroiWOFWZs/O60zrWtIQG7d6ToeYb
1vdE6MEItgHq5aVKvmpMKGIdw88FnNvz0SPnP86YgCcvW01pqcDrfQ/Sf37TW8Trp/3b8UDZmjhJ
yGjgaoGNbjHz8jZyc6i/Zty818vGeaRrrwKsURLf/LRUpsOzzUEfhQQimu9BbhK05pmtOLMY3+SI
j+wMRXEbXmDnlG6MvawhFHqxQ9XG1BZGacpb4E65QMu69yOjnkzTN5iHEoFu8NXC+gLfdtp/p/SI
4sL6Yc9snzZuUgOg0seeAuOzQqkU0nRsq6HRHQlhFcEClf5bO9SkdYBncpYaZ2t+N6h/hL+5j/I/
PQnqXSdvLHo8qsE5//helqp9x31/STl+gLLS+cXR1NcAQa8uEU3Ybxa1tc9p8cb0ME0ynKZz1vyJ
Z5OIKQa54iuA8DNGylK/DMByiN8f5XXuJCMaoPCOpcNgtZMm62ZEICbgahZts/gZddcXGrvpKibR
+MzQEz3Oogw2Mjm/xoTJkgWRdfzvqS4nrKIwNZbzhZxzEnMymToWG3uAhxzXG3znBb0kqDMQHQ+s
+xzqFDecWugAY+0Zhr+a9wjl2tziwaybK+qDEAmu4ojwNioQFdhYmPN4gHRs9Sg17s/yA0rLr/0o
npa956DQn9G4/fxsJ+6zWbdDDm5bowKCkb6h3rs39tN8i9Rq5YOjtsf7j3sRcsQXsWQdaoCjekgp
iuIClEyI7i6ueuBu8CY+llpc0+ppu8p2QU40Ne4JQ9y0Kw3oabZEj5KqMa/3G9UHzlvXkTLbfmN5
Mf/FgilDN8jHVTCu5kXhp64pG1omS/t4HHHQhKZvQuKKs8Z2ocMFYG6PV5ZyL9In3NdQCb5eG+7Q
hBnYOu7ZGNKDLeEIsHGqPsfKRuuwDpcpAqTuRMAuGAQQc9sV71A6vSOMLu0/K9GyiIYhDrElYXiy
QbOR8wV6oiXL2ZPm5Xi8yE+vookVQnukUCgKjmwkbr+PMGlCLTSjDsaFciTSx1/wW+PzUskRZ34r
z4jAsC64rZFH8ibVyQm0AdVVqvmTWxK3HfkNh9L9Pv+YOtowB6IMssVwhVsf4Pui5q+db7oEGN1X
qgaCrmjIhwl5YrCz/e96mq9OKpzo1Wy6HgpKFdbLSzEE8Cl83nPRvt3EOJUIx88xEqVJqKPuZaQz
zDfovb+FPBh06Ml0lxt22fXpK8iaKKb88NS4ajhIi4y3NGzS4Debhx6MBpLcUFusr2vKd9SZOH9E
q5lQ1GVBg5zgOuAKF8JDEhSO9Z9ckn53UpTAnUaK9VxO979fso3DhbFn/jLSIJcfPx0T01ngp7sr
TBvvAiO7Fz5ogrqMiYMHaFar4g7w7A+9PJrT5IrsQzvGR/FH0ORDimr+bf59pTH2jlcACOekxJa4
mBAe/ops3qxXgSyodR5nLdwX2lYNiWiFxJMT1d2m4RzurAinBYa+HHniG/Ni7EOjcQBRGM1GFEZf
B+SmTh366MGhlT0NTZLMPcFD3luMnlGwDVTPaOabp+d0+CQXIJzmgXMPlMriOdKQGYJabMHMJRm8
V6oVLfRPz5O/0c8wXPHY5rvvUCYmMu0w5UenmQAMF3364g+0drd+PAhzbqSd+Rb4t8vYwifQ5Axb
sqCN9Rt89/Otfcf5krVBdYhO4xbttZhI//hOM+wSZcEwdJnQ0a0a8uDVQy2BSdnXYaAvVqxKFkak
mkcVaAo4QQVtOBBMJ0KYpzkaibeXTqyQ4zVR+ziwbVqaQdYMDBjQOO/W6BQiJflLafP6y5XYiwMM
jJgoeKxnswiU8/FA/I2Mno7d6CunutIJ1vp1qBRaJMj/l3f53mqx+fw1a4uP8bOCrZ6ZNCS7U8qi
gwl45f2cbwkp/J9+x5rZbnEWc+jtBK7eLKxbIDScGijqsybNdmvbBCKCHEkuaoE7DPnz5eA7AoUo
2eho8EaHbsD9Bdf8OJng8XIVMvqz/77TrKNNqulSWo13EweRjnhbk5D9t0PdYuKkOYcpc/HLPvQz
tORgHEExTcPJ9zUqhNctyBSukb3cpdMGULZO3PgVaFoO7ZF+aDeSHfe6l6wiXa6Jb0Vm0M6oxjhE
gRWWQeNt/6Tr+dLQGFB5xwsQjogcjh5LYyhGdR3spGfUqPvvekkcqV1rGWh51hO0J4kQdcYAfcgn
sJLVDy2vy7SblfbUSRqjpuuApLynHEVFkqmZWF4EtIqDBQ5wFRDJa++BmIkt6fKGuHw6TRIVl1v0
2DlrwY15b9zAMaQuTrPuLV8xHzwphEljy08Fm+enmBmVsd2NcRSoMpmMW6fzsPwonUPKEMZkBXlv
6EU6DZyLtUukZhHbFy1fiQO/kUgMCjpqLMQx7S9AggKGMCTva86ASBH4sHj8F70vYX2+6uKDuUk/
3ysfw+wgj+zDLUeXIXQit4bq59wD3E1v7JW7TrB+RZkSKB2pUfq20+javXaidSVhyTgP9um1erRj
PMRzyJ8UyoTHNVD3TDWNBwXst9YDq3ZP6TrUiUTfUuxr1e7CW9IvaUPkaYefAFVYhSYJBSowCVs9
OuLzWPl9p1K5V9t9NF7XTwUP8O4n7kof4Pi1yudc770ZVMAbjLoA3RIUbHeg/90aO40pbr53WoMf
X/vLDnD20ZhEpxd/plkQ2Awpp5stzPVD5BPmEuLXTIfHVgUvcVSabtBZivGdh2xhp6xDN7K6Zbuu
5lxr4Uh633SZ88NSkkZD2bAFSvFEDCWjVGrU9/F+lBEkjzZFGvwMmDzfmIApBMfipqwQmHTmypRb
Utk/fClRUB3cNbd4Wehd0YD9I05bLhAD4JKAaBzdOvmA+UV9IKI4IOJk4Cpq1YEsWiinKLPybKdD
SBY+q/lXBHLscz1q+oBgE6nQwJpayOHoTjLnlPyLkV4Cv402wjNtvuXu6Y0FpAovyu8wwKgXC8Hl
pvzDj7Fma2woPZJlKW1+HOlCQ0svk3HXj1MU2vvPuCxuChOTd865uQQGQgmSt9OTtSU+ajdNgpkF
CBN2F3+AP2VsRyLj7cmKtxX8qCKHeOOsbprkSECgzg7w9c8JhHqHZ+biCMKxBdEltbJX2YI7pKpQ
eWfHr9PXSnef7FTmJJ32AxIKzBEu5dSpn3sbuUbG5znJM5rvSNSTO12tRVX7rZaiuaixcotisUtK
JN7q3YM+Z2cqsM3CvL+piLrE4t3d+wC5RiKPBY7AOPgNcXJvBrgWCHLwxDny8hrvJsFTRFpvtljp
dArb8sHZhwUn3SO3lVyLJQ5DtFhfB8NPnCbLHtpnA163FyOJ+6svY/UEHMxcSURWSFBLUTmL2GsU
eJK8GNcdU+1Wyln3uYBQKPc2BUWcIo5S8+6H8aBHdhRzSt284HBQ6Rb9S1a0SkKwPS1yY8AvPBjU
/7iaedWSShSi7VSd4t9ArJGTAE4vYnNcFR1p2aH0QPlgtIDuJD1LxsEa2m8cePwjXXCdKLhkf6Z7
1WONdpotT+Otk4uNL2HigrsC4nHJpsJ2NkTzM6mzh7O14pII+bMLNx8IGx3SkPtLJo3nZBQjTkCO
jYSACbV7oYTDGwBLzMHKjp0eb/yO3vhmQJJxPNbROSuSaITHHTgwAGAuC/TQvPKXSTMpd/S3KhX9
WCVaPuYOaw4FNBHkCegn3dznNdEwUzy8M4mMwQXZpMgmoAxDY4p4/NnDIDLjXnOfIrNQZdEqAsnP
rf3HPCAehArEpvfEw0FFFulL1ZEKlGuajtGCwtN/ZkI87XBKw2bX9ODURjrcIvYBsrelHLYuDCYp
UQ2bKr4ecJPM2QUjH9Pji9mFzgMWoGE7eaaCIO566EqaRAGNXZiWRPJI9dINNu3Lg6wOtoQ3/WNT
URc9k55ovQwoCrwg5JLooed+gGwBeLfJitqhIo06yeIEol0h5Azkhh+7mSQLTcWLvvUO6Rn04JNh
l13krLe4uZTU2icWDjx3Mwztza1NliXiYxa4i+y0/+VY/YXRuPfCPL2cE3tSJMoVW6BKtDd1ahRy
hVgb5vBVS4+FOZonb1DluUhJ8qgwkuLo6Hdx4/Tnyp2YHZAfwIf6mldBYrg8X4iXVx9egjCqi9Hx
ftl1enD9tTCVvTcTfZsuSAwJy1jtqVPeca4SqBV6pQrZaa97rLtIWNLgawD0FSaHdYNvkcsKjpUe
v6haDaGDLRTnJP5OtSvu3IUtmUZmfO+hlbqsmaWa4Em6ijyzF3Iq1DtypJrwSqRiLCchWx6YnBca
YkZqzUjNiDxz41Hblm8BIkULHSs5zy0+RVaCweXyLGe6s+HAmDrOVmqFdENI7K9Th8o28UkpQfu1
ednpkUTs58rk7AXp56nzdAZbKjcBjJKJbj5vAh8hnSOFtBGkz+TDfZIYEi3/MZKTfHWOrDgHMlah
66MZo+tMnf9FmkW8OU3Bw4HwfUs6QlBowAfPIkccvyftN7etLQ9TUhLYnAnOVSXCEdYG3CWfzPt3
zHe+j9yLvddz6e68sr5XKrZOTrTpVrw9GPFe9YJXx4KZCJzE95RhJ92WwMHpp5awZrwKVVLzmK07
GN07FkIjUeMqMALM4PFHnZwdVGouqrdPWwRgdXQ/+K64RGOMvhe5EhanDpy4QHciqLdTTHUNnYZk
//NaqOHBajhZ9/Nlf3B8coQygzMb5Ppw0UwLGszOkASavAsHCP97a6q6aEYjeTBKYXKA7y/7/YEt
OalnXLj0XxBZ6VmuWlWrFl5n8AIZDfkwAZDWMQ56cJJEJ0f4lnrlKCEndR1TU1PimL9Rv6ErRL/5
GWyakpLXcPi9CDhTgdHlNTMOzO79UMWkGT4slp9Kdc2Qt5V/gRz8f3lERB7cARXK6XGZ90B+eTeb
ZF0bwDWvtNjWhqrVVoGEq+tHzF0DeybgmraJFR+pu6wsW8wJffe8poYJ8JFLOcKHCltd8b7MhNyW
eAlT/ZlTx2BQAqUMvxyCq5AIYLxQzNJL0aL569SyEE4QLgINclxjmbK7p0Rsh7domT5ouVsb/xUD
FvJSPklft4K0ZqVZZDqVk8SBox5DdzPqlTCdFCSCiTzo7VVyBfqAdj+YNXOTVljwZL9R6dxWLfT0
1xdaG9Wz/qIhE5BwxRCgFoVjAsvgXmHdZa2Q1W75AOs1VtkYzvXxG5xXv/TCfhc/jckUhWoC3fNv
E5PA68lr57+oqZRGocdm92HNi9mqVBgHCVlq6w4Fg9BegLOwWcwlyYEZicbTVZNmIaV1zJjC4Uua
i8bYZMbfE5ymQM7vjMpnk7jDf2GkED5HtxeWyTE1l8p8NYfjEGhoUGe7q8feXRmiuowlxnrrVtSI
xcUa3+EZAU4w4XlSxm2IRNAn6pVYDP5EBYWmjudRxRYPpT8g31Mooj0XFTc0X7/oHAKLquIAHbfx
i72SRqrnsRKYRRCSMNx+gwql8NldvFiort/Qb9P6IeFjrr3Juz0FqezaG756Cvhgpt/bFuiD8dVF
OArAzTZ7Xs4PYQhFT9Bdtl/cOHq2U4egXMPSyN/2HcNZY1VfMTtONDY3lTTxm5MAcJyxNde7x+fX
33sQVKwpAz6DQLWcpyX3yo3WWvWSy3rpgQu2giDKfPSyV39+Mr9X5cg/SM0Yfhdz59Yi/niV61tc
OK62gacI40WweFJSbUOiIn1qJily7ZLvYVFtQlXr9EJiQEzDIetVB9cq5sinWHGWT40LjYHMOAzR
n/vH2hHwcdRKbUSVcmIoDMplOEPQ3ShKM0FNDo8nUkWAo+UaSO2CVZMwWL2nUIFzrgsK/Sp8KwcI
gDnwgSOd8lBLXVqsQSEjNpO/8a6E9nCNVbXOn7DupfWwmevjKsdgE+V2uI5kVxt8C7+UiPw/h7io
7dDJzziSO2QFozlm51l9wrHqukew4HxtegmuMjQgCt3V9rzfNKl20Hsc7SDIMnfOFC6QjPwdKx7v
BwinDEG9ytuhZUNnATDjGPu1MXs0xnU288peCMkvFaOrKJsI+BZKLoLKWJalK8JpTZW6khCZCrpB
eKgUwtSFEKLs8Rz/d+5sfqocyfGzSiv0WWVqJ1rp4fXx8bWQbGqUC6Pkj/Pfkby8pG5TSWAhNug7
+wBT3L84uFWNKD4K8ztTlEL8PYErJ0UnNsEPjY4Gp/CBGPag9mQFu8lFog3UYjAU4G7Hjq2caD21
QebOHkIlXiXtJTfGbmsq6CAryK9dSO0KdAABD3bd+RI/71w0Ty492ijXdSchvr5gJROYVOHgyVlz
BQ5KsBF188ftwvdjuISDmgsmwU6IHx6+8gorS2jJyyAQUX6x2r8eAVUEUt6Pus9RM8EU7mYTH5Ym
DXpgtsM0/ZMoHBEKyTMzp1UKlX2Rgpj+H8qiBbmEtGK/GZDH/mpdWq0Fi+nzIbHzC1u71xgZfPv7
qXXQ1R77qb8rSu2FIsnt0KpwySOBu6Qa2lADJKxyZZUoGD2A0EI0WtZPJZHO5F9NJ5IlpAgAe4Qz
d0YkbzqO0nRor6qNkayther6tFoSneuXQm9nWigfmdVC9xrF3fW31sloDO8mNmIcmG8EiW2T9WQF
jvBkhWApE18SFtwkDHgb6gjdCkshFySBGM+qM8SjecsD78j/2UCsNZk1YiEZduc0XtQo5l8oe8rA
saDzxfa26O0alHUUSnaPbI6U5myj9BgWbdXGurWKzLZjId5S41Z5T90GOrLdPju/slR+jaLeooV7
5whsMifrXCMEErZ5c3zCWWXbRsoYVXFBdie9ivlSm8DIM27yE7eZpruWubIXQjsGOHFfH1IMOqN3
CRfOtodBdCCYT0Qn1Ehl3yOhBaATAAVnmEf+EHdS0onwYPKpkayZfPtAb/wpr9vJTOexZdHz2trc
LgEMkDtpaz7Pm5rAPqvJ+tfEmfeO59pv23fac0bpaENQEChQoV+CLqnb/lKcTPYN+1+qZlj9lEUv
h8jigOgdkYjqkngmtxB750EjbC+yejI5mli476/vsjtJukScvA1qehWiXVtxPEtEq+KFLa4Zi2NA
OrpuzfRXcrGIlLjM84TueLnTuygIifJ87P+Iu3yybpGFDaHxBPQvQiZwvpd/rmXLInvBVl/cyOs9
T5O/mw6WQHUCo2imIj2M7uFep68n8Sez9HasAgxEi57qe2kWjKOGe9SeuoVkNoKNEdoFCtpx1Pye
aL4/8WXv/VDSJFLGG7y4cR356Luu5/1vJArDkcA8/kJyvdmF6pnZTeKimCxdCuEM6LJsdFUllUKJ
9OJ01zueEPZ6/rInC+rmA9hSH88sMSM5xXLvZjz0qydIOzSFBQesXxbZH+tM4rqzEtj8BHwd29Qy
EkZuOUd+jKp+3j4ZMCgBNJ9DH/fYPRXRa0wei9+h8MWtLmnNEOho+WkNVsHOKlN/Cy5CMY8VoBqo
cOZQhlE64M1O81vy0lIzxapvJ5VFa/Cx4Oc4GXO74EYGIpQK/+vZIqBJj8gIHBY2hYY5jpXTzJXr
WRuQMRn57xAPaLOdlwvFqlPVLewu+8VE/bvmhHdV7yhShkL5LwAL1Swm1yRtx8FaGs1umqKkVlLk
ahfw0EUAzaIgZCHc2Af+mPqZ3bdo9d6u4ds6DaiB3oW7aOLOgBwXv6wU3fZhtQO+acizrnvrTiY/
xcXy2Glh+TuXJe1Eh8QCDqvJPKtg0I3eGk3nLfYNqZ97we4EsWcMbWRfLxHg0yOytITJA/EC1KQo
tzUPSVlYdN/belpLs49zQmi9JXfcbfW8/BH/uTe2cZJ7U7SlpaMiApdJxmANB/jFvWHxLd5q7L48
Qi6RJDT1VhwkrvSFNE5h9fdJSq3JO9MCI6ZDvaZOJVkYw6QTrSWvdaUneX1OpacLnbyZpGjZH8Id
/6riyJ3S3d9YpcKS7Wt+bj3Fuuhq7SaPxM2ez41NhBtSvICtdUXXlCADCEwFoZez7adjxAruWjyz
VPHKyv8hjzKdNMYr38sXJI3BnyxQai+7L2eoAEUcqiwbsiVPDZkN3Qy+fxuuuhReNtHE1ZxgH6rR
f+63KCWTlVF4cfXTkjS9A82qMUuD3+iFakUanoYAnvdEcT1buYrW32iVHjoxB67WXj2lZMTxirch
Ida8QlKbuxw1ETkQbsglIIw76JRSaFTAPqnOG9hRTswbFx79u7gUI5d/uv9TXbWIQHVdibj5EgPr
GJIdOohT4zL5KDyN9ePMhlaq8Q6zdIukMsi/iw4WwJ+X6GCvoJYDkUZT6lDUz1WbHsLBaNRm6lX7
GeCL6Ol1KYf7jZ2NnaXo6BDFJeE1gdyM8LxeKjSoTLt0BePZwF2XmcKrvN/v3yOcZgKoX4qgNVmQ
Hvap1bDFLNInWi2oZshZdOqFJkqzkYaaStnr55K3wmY018NiIDKOAS9HgsE4LQNihgI4eSBWVMWz
2rlVnCF0dYyn9Q5ZI5boyF42sZfJ8kzH6vMa7BA/YdyF/IT12+LaDXjcMVSYDuid9zQiT+DZ7Tlz
8q92H0kVjtm5nbr0DNsyaylDPTMQq2GG1scnplTwrr4oo8SyEoljz2GGMQGJCS/4FZBFhm2O5MnJ
D20OxGpr6H//+dpYsFKvOzM+nKPGr484rkeblq+OK+mMyxa9ltj0xAwXL7iZrV7LftEKplD5L+1t
xevCooJbK9a4FP6GAe3udG5LFqmgtgBO2JgsSo6we/V+NML3+p1iGZRb0ktbFCbvbQh3GId0bsDI
k7RIihnY1kLmP5MIG6bocponBLLmMTReMgb2ka5y/CW6ZOEfgoMVRTATvhLXKEVj8Av9Atk/SPox
rfAZganuYWuHE3ZK/8syXjU2E2bvpZOUC0VIBO1wF3phJOfIQd3+F98UJXDMzriwE7XAS6mJUdEQ
6s+DH3GotX32aok+n0HsS1bM89rgU/vCyuN7sdc1tNPbIkL6Inrz9wdBiKpqhwGBabQ/gnnPRgsc
Rauw92WS52W/ftSFw0duML0ApdonwyyncczYhifaCKQUXqJXFclwf/QjvbVYybnNdSRM5p3/ySo1
3gTp6AZNQMOplWay1+fMBIU0er6KCcaYxz92d6SJfY2JdSlNFKKoX+v7PcW9HyvxjPfRpsMRgrFm
junn7nbbPairrEkB9b+Tz/oKKV2fBaB9BAwshAeD8eyfbfTOfiG5K0K3rAXYrazehfTO1uH5yz9B
yYHTp0FCzW0Lx72YTADMGM1I3RLkSO9UGommbx3Ko2CAVkPFpRuicbl3K3T1zx+vui4hrQbF7bfz
ODV0fQhAoN1NnaOMKdGTh6hvPj5+9qpjpXp1DV/M85Nm+srR5DA9gx3w76iYyHnA+t1mChfPIyUE
HJwbsvTDKbXi3hlSxbIxwAAKSjPXAwdkNlF0C39x8zDXOiW1F4f2/djTUqWbTYifMje63ubzXo5Z
GH8YRxJxPB5Og1FCINzVWn5rAqhDkOXLH91zQv8fG8tx6ptxEkpUI61Uw+SIoW0Yg2y+FmP2cOyR
yJGQ1vGlWFn7AaKUIk/lgljY4oOP3+zMD3X8M6+X/7AW+Q4AYwzx0rY9xpGZ8pATmh330MdgRM66
tqHCDIK5dRGdb9+janMVzxtmHbB2g6i/Nus6nqqxs2aoS3F0385g0qh/iE/HjWCkWS3FQXsinPyL
SpN/bQcHDxtE2CSjGWjNiw5XzkfpDFCkght0NA6qkqIp/6jJcRjy9lOHyR03IjtlffNppEqOYiMN
ep1JtW5eWWH1jJtJhAhPk/EOdC8DMNKEO2YhXD1v4yvU0fBO4Fv4gElljcBn0Fxdy7MY5ECtCW62
ZnFNPXBfLLylBYgXhUuGMg5aLmkZwCLMo2d9QMHjaJbiV6eLtkttXduisYtsuusC7FE7wyoymmPC
7KMstrF/p4bd70Vc8wYhJAGTeFbWK+hnD+ldenDv58e3O1UlUIJrqbp/az8nLMCksm9v6scY2V+z
KyXSRdk57KgXOGvWr3WyPA3x3ro5l3Ol1KNDtmomi4wse5WWXYrdjuyuktHJS+SJL9scaROPanBo
9HgBN5rYxVlMO35YpQ6l0sCg81v1YnePZ2ACATqK0Y8cvMMX1+zfR7/+977AZyiCMGBzcp4bzdd3
W8RBAK3VwQm6YABr71c8pF5Haird+gDOrMovJdl+QIf7Y3lhOM4FNCL7KvktNMz5m/ivzWVbmwvA
ZYQxEPWshbV/w+fvAqnMy1ATfjRcsC/PxRN/TRwpbxUnAUbgzFMBu8uytXr7PyNFGF7fSipcy9VL
3xXAuVC7DlCMr5i+JlJk0h1+m05kYNAKPzhLp5JAOurTTgdxSZMVImeOjWy4VNnJaqLzLI2wH0r8
6VL/5ZF95AOHoLqkXMQLR9LvjelW0/XZ3rUoQOPrLzPoSeN+PecESrlwDB6XNYKEhNiVWwUe59wd
6H9XXFfTeaQ0JpeKP0GmNp4nJSSmWJHfNggI3FRuII40gBPeEdwyl+RhAGNwDjgfPhGFPArbEqXN
RNItNn4VS9aaKxB4Tn8i6C75lGVgy9yRCXww/iMuue7xGsswWKARxOJa6GNdsK2/aMQ+du+p+Zi0
gTqHfPh2q+sBd/m9xB+c/ByV7jR/AZAAipzVhCWcVQ4oU8yvSoeBaVliuKtaCz8nHKoJD7uNJBof
VONT60p0o+ChaEM1easuAmjE3gcltceG1xq6P/LHzccG5wcrEuQM6l+YJBMSLPoBWcxsz4qdPGCt
fqouKLQs6gp63yxB138TukZ9wUVOHG5my3s914kVyo4RTkzZA9JQfHrSSkJ7XK2vnItzZJYBt2Z0
qZ1Ju0lGrSTRJQ51X0Yf7yfWpQG6K9fbp63c8fSMNKhTD5y3du0W4eYg8E+eTByo1lVg5jxPZQfD
mhyKfWbc9RN/pOUG8qsOLCMW/8xvcye6X9w0zl3CIZObCn/HGomofswQL3dhUKq+kNC6ZpyFtVdN
7945Bf8t9P2cdHSnnP/zsEKSonv2dAVQ7AbMAkzNxqWBPVEjO+c4zADubefeP50Z4f8KyIftCWUL
JJHOWvBk+XnxJ5WFuk/DCZjiFL8WXOkdMNk+UqWX+MrNLbgwkUmEjqKr05y+OfqV9CbhR51H3poB
eT/IWRkWwlLMh0TOZMhLteyhgK9ChvPtADFeipwU0rS2OY8FrgX/uqg14LYg6kDJCy5AcSzkE7la
l8sQvMMYcw42nJHKQHCgAhE4R8vFD3t/Il6r3zt47WQEeYH4jgYuXE0oFtyjyr3YCIOjbd7Gblh7
vvIjBdnuOvXESMYpgDm9DeTxfMhJBllfsbH4hFTnABiSyReUpjllVIQrbzZd56qKcCdFC7lwTtj5
R17i4s4u+xYL9ZS8CFfx3LTRu/7EOmCcJF5feCWt9QsULrBkx5G2OkYJo+jf4wrGBCv0gQVSzCur
Q7G8fr1L0fSRwzs84vPy0OObBQFNkKEZ4qVSvsmCGN/ZKpAHI+arO4VxQSDQxSjW4ZCy0x/jSEyy
dJMdl95S5qHByZfBhJTvg4ViS5reOLy16lkdYbLXHFnx3MhrX92uYs5+XhOsqTDLen2VTnghczzQ
uwimBRD0Pn+X3XMM9yhQPXrpk5DkCdPYi/icB8aU8iwr3mRr6Qct/7xieYIp0ifc0Q17LUKLRIqe
xP9jtak87whoiBte/ytYVFBeKMBzj8QLbc2FACj0f5c+STvuNG7Yt8cDtgMRXPXhPpJ+/A4Lawwo
TvIOhlscdqAVX2jEdUUgOOL4cPGVgyX306VLoLX1LNhGmDZecrdBqc9IgOALpVbUyG5zeIbwVT9t
GLQCDdYh7PhH37BrifBRX+LX7cXzK2FAj1GnYgXVselXA8yoWJXiWpDbALnXZg6dt1K7nzMJz7Pc
sd0UhiH9ulk+zDe3fHv+GD7Uh3lA1PKkOpvBdHIAbJfyzrtvidKiCOyljvBw5WdjSBes7Kiko/3J
YyffPwx1sdqjAFZI6NdNA+eupTmI36VVYfZjjAwMxuf7CkXXdjJgm5dvB8mzWT5xme57VXfqvISp
VATHgz47pCqHOFrhzmcVoLPmXhnosJb1y/CClJN2cHPt+3Q8eDWLYD/FsiYc/EfWVXspA63RY+Vh
M5jfBiTefbGV3BCF/S4k5xs3UmtYy+Yip45+wrIAaSbKeYWrkn2BsNiC6ZF9yOVZca+nBr9qF+Ex
n0nOs5svENDApe1Cbvm2YDAQ7sZQzYONQlXOBjBEUiFYm4bg7nZwq0Ws3qtdbm9cysPMbALHHWRW
no81DAjb6iEmYQf0cwwZ1uH+3q7yQ21zU3pvcG5lG6NEBXdATQsLWw5teVKafUf1frd34F5bny8M
DqU4HK3caBdPZymq7zTLcFNRN4h34I2w7XgYcve/+E+3N+S4WeuKYM5RyDBpIEyzVakitxriunho
KuyVw3utjyP5J/m1H/ZULLcsnmOhyQ1/dllQLsbmfjIG3t8za/CTeeqsFtjKRmQIinCkBUm4UmEF
nHu0EDOVOLh2vtCrAiH9zrQW6ODJ2vYrk+LgaI7YwM3EfZLusYkOM1qArKZBb977YpYWPG00BHem
DTEeVvkUbggPZMyMGJO1Qdzg5Ff8TTxRuYBB+6gbsdER4gc7LQTVXmSU2QuBYlgZu/YwIdcSsFwX
ninal30h4FlFWWLJZWfJiWeFi8mUxyZua15HqctCwdoORO9KNTa4xRedtbtyQ5iLTpnxhaqlfF0H
TgeTVEoCGdgWwZBhiVMcSxYkjscYj/TPfTVj0TZs16OLm+JGvmLxF4b2PmYmh+/Ry0ep53Z8dpxd
X3tYicriS9u4DBdheb5TSegaKwNUOzNaCYdChF7XyoYsTDiaWVZFmIU/NEtpshoSd9JCioE0R76g
55w1jpgvLugsgblG8twLObOrWlvTehNZhw2ofbxBUE48Z5PK0X/ZayQR5JsF/F1ObC5yxxvebM4K
bfuvKrrdm70rUIRaaESfWU3HUMzVjYlnuK6SJvYkVnFU/kjMNVQVwJ7wQKgdCRApanfj6BQ4YJr5
l/PV9rZpZYL9xuVicJ/kHDzQj1cbSJcHzXLk6NFKCMskSmJ/f6lYkDHknjiSyclmndAF4KIX2O51
ByA5fujDwI2fUAbaji32C2lbd7xLv6MSoi4zVmWJuKyzyNfslxpqlQkKPUFq8nS/ZwvJiMp5re9J
7frDBzQSaCq0uOt7fKFBWr8NViyHZLbhDnzcpJzayGN+8MXPCLFkN/u/r5xqN60sR2PlrRRRG4Kp
ZL0Z6rgrE73xtU8e2L+HTLOrerHShSZ7wFuq3U78/ct3XgzTMyJEpcKoiP2CRP4uuuN9ihbij/ih
s1YVTk2VjuYbnFS5NdpdQBG1FQGL5p15kKkHp2LEU5r3pWniORwmwsAZXkHrg7U8ZJ08Wg0e3iGb
4PGqNijwCp+mwraPy/SQi8tCoVkpNKIFiBkDiBWOqd/qZWNLF2H/ODI5szio7VIKPI5YI45h9Vcu
pANwgRp6+PYdfoFcFoRuglecMb4Tv+fVdAqup7zOs9XqQ5lxGszZkFEnpxhUUrWahHh+d/0NzlkT
K9Hptcr4Z0TyJucOUB5v9MAHolvGb9Q4mgwKKQvzMK6svRkMJ+6xVp3JgJ4kqD3XNYpmy8jHAuBq
3VGoulDrpKXW1A6exawdNTispEVn3IuSI8t/Ocx1oXH/Y1T7QoFzXY0KazAr/XuIgGIAU5vgRNb/
Vi/Tk9TOizcFZ5EE9rWHWwUXpDVpJDVXNRRz0vRQr4NbhoZwpJwhWN3LtrAIM629lPkhbuOqOt0J
S6saAy9Txob02++COpfnlGmFQ48Cg5NpuL0YUSLwfrMOZAqqUH+jvYfNisKbxgWHJMkFNSixAjti
nb8ZEuhXaGRCVkW7LM6dDURGHgpY7ZnXWuxP/0KsCkCpjbG1kZoHLF6Ucg/5LFHsGSqeANrfUMXK
rVG7v3236lT10XLBfNt0yU+9qDxN6wQ+6ByWNmrgFMbgSy/0FMkKZIDDAxQMa1bsj3w0xL9yOsRU
EcXmAZC2PYKq9DHntvVw6NOruZxc8iKij2OMtJtUfEfqSubpls3UzUFPEfl8Pq/iqbN8vnHdpb/W
XfmOZwcP7V4hPAoFt3RPVR1Ef8lyrumyiZMOqnBAXnIbgEUl2RsaZuW0dk4nEVu1/F45yMesP1bU
wQ+Sjtmm0o099np7auaVvyiDIAJZ7kwciyhoHYDAHZfkRIRJcdApfINw2ruqm0K6pP9FEvnIUTIV
Zjp99YZxFfcdwAYKzuEBywLbisGDvtyeCfvJ636zD59BYwhjizc5al3qrh5x1zVjYMQpg2JVb65p
iZlvP74BMw4IFLNGTMMzk9te1gEjQ2xjX6x532Fb1W5qCN7lWPARok1je8YU86ImgbUNiqs5gTLf
qq68B5vyBz+2fef08G4ZsMeqgf7Ku06mxK9JS59tFUY1VIn0RThC0pFKht8r+10N4Ds4y9q7jQb9
HEU0B6sQNhXht9oJpRlSOCRDfBUctmJAXWXZnBVhN7HfKr+PT+UeLIlAySJ5Ly1SFereqiR9248Y
tffOUHqONrkbU81dcppd/+i1QTlAPW5rbXL8uErUjpvghWrmiOb/hMReondJQ1zYY8iVZc60+Bsy
3qta7zl3zkxoBpsc11MvwC4uZD9EcXvSVQgHgKilbq52GbCkVzSCDuFMrP2NqhjlMUXY2904YOdz
fJATHjJOHhy2HqtqzsyGsYrQ5wutoxfhG2zf1wRMonVhLD+ZApv9wHN00v+cKFQ3jjxw0IAbv4Wt
tAofmbbIsuuI/5AngY/Bgi+F+jpDjGupMgPrjk39BafJzlYLYvWw2XKxrLE5oYihko2ztgeoE1GT
KEHzrAMt6RJ1zI2d7W28kvxf0XWQTch+fzwQtUUEGtKmpE2YJWjPPqy8v8QwBaezCBmp3z6+YInR
LUAY9JMM7KgOxh9tyPs1ozKRen7R/Yyo1xCc5MqYZH1KVVIK8coVEYeF6obIixCU/jLOwpqmmYlU
dbxlw70bRBoOEJexOp7PC60mzUs6PzzKUVI//VSIDrKNm+6+HwP2l23dCCQ2UeadxWqdYLPM9Oa3
8N+h9crEfT5C+XXcbLSvXry7o3UrpJP8Q+YvxalnJFNhkQoPIpUO4POggaggS6BdrGUrFgegDOlz
ZozfdX5txxitIjIumI2a0hV7WN2FyfGI/XfpssgRMofYW1kLvOJzTyfssYuDwN0GO8mEH1xedXe2
NGOVPvpog88Z9MrNdTeWSPtUcjtWBrLXnWRw0pN2CU+E31Uc5Yyi9HiFqe9h5muDEwsJByxfUH3z
Q3g+50sU7kGwd22HfnyrYawmbS4PogVVX6PC59gMgW3GS4alNVvCFi+DUfSWA2MqxB06LAMwd8TG
RHuoUc/xW0/2tmdvZW+7HKZkcZ2yFwCKEGx03xqG4MlYMv3kWe8Y0oaF+u4XCHlVfDFTdudxEYZD
SboegPAY2pUYapKFxfkyYQwQUVVfQoGPcJHV8IrwCi+nk68JSr3FjdxkFzlchCpCJVL9KAkSdyAw
Sm6rvJwBEJaCSjua7zZuEUgEztdemF+qjgaBsB879RgC4ivAIcaE6YnDES1irSbSZD5QUpeyLVUX
S4uZV+DkweLN+X1/L1jYsGqBOVnNbwWACft5JYa8VbqzkXFa4kHGY1LvV1gRqko5aEOfDc97NuoO
Mggq/rpqt0jHD2DeZ/cfIuB/MepSlunwgLUGi/GbP8GWNPzvweUA9jHbnjKQh2Hl+AUpFPMZRPu1
zDqbfcS4bIsY0w02EJvpFa81nH8EPHHNsdBbR2/tiVkXVlBbGa5zDZ6ypaLH0YAKpt01qlnHTSWT
SPDNka1jLY6GcCt6d/uoxzgojAesiI/Ww3jNvTdAml/nlaQkWiYiOKR+hePub9p1ak05lKe7J8X3
nqTpV2/i/OS0ox61qacg4PbPJlmCm8pJ94U/n4JToSt3hn/vse3PSb7eF72U455O912kqdvQKUWP
H5qtLuhR4LDqNIQbCMhAedFXHY+U7N/+v/K69+16xjjuU7yvJcNhpRGvDX6V7/sbgLdjZdV6Uz8R
Nzt30gn/kbubB2T4eur+2HC4w1lmugmXvbHtwntKxqaKumBpO+4wdNtPbWRfWPfz5q2BOxQOkVq/
5jlT3XvJEZIbGNbbegxiKGUofJaPDVD810BsB3Gwjv+azYi2zMzs8siIp5DQGc8e5gQWvGpLQBvI
el2MN2zuQFnxq4CdhI18ZNDN13R4ML70n0DD6/5ESOVNdA7rf1ralFzzaNNuiCoOIej0o2NOpa84
oSDc9gT+JHHVOg3y0x0vRDrqgxzzbDrH9OC92xgbtbV+iLnxWnqy1lY7UpYvr7vVg0cbTklZ7b8l
SYAQN2BKQ8Ut6SqIritsQBdaA5l9LNtcfSKUG/D3Arxwm/XmoTi0kzbiL1JBVtkV2s8nKx89VYEA
qtqMVPHaHuby32bydclarWO29+UX5Y3Xq7T4890QQ/4TegBL4y3IOmeaEjDUCgFRBkIvip5utAMF
ogKV3i7OvVZljryFVnpTiP/AWrZK4gQTfmBIrBEPOniB1oIISdfpYDpataVlXGiSNjXcC2EksJkz
rn1lEW9U+51ji27LgXtbzVN+4AGxyQlEdFymX9yyXFvRweW0ny0WCbJ3h20aoVopxYvAByXm/p4R
tmaREGhlYCCq2cCB1RiOgY7CuyVfD50nHL3wQ5grfPTDuERQHt1fgqZvtkGIrMIw2Mc9F7oPzhSZ
vrdSuKBhmN6t+qlh+KMl4Q46N7i2j5BtWx3KPZ2w1IavrsA+YzvqLFmqWXgP2KMvBkHU41DFk4k+
NshADwSqS1IIS0nXAUoRF3sNzG6V41FRY8uGoLN6hVNRYbUvkeE4pUJB1WJ0HxT/WRlRVHjKpRUx
+xtPByHl9q2c4KT5cTJpM1Cpdb/p821iDE9DkNs3IxNfLalVRywMW1y8gI5hfV/khCxZMFSIMT2z
afRbkCOq9U0evpmnUEtiLBk3OXh3LoZw4eJHNCTtmcUTpkyuQQYeqEoIOWhQVmm8yjhTBx++H3cT
qFo7AGNeBQNnnzBmDfCSTNM/ANVPMuxQ9BAD4vxdV/3ohJjGRb/c/Li3pbIgIUy4x4ua0+GyHRjJ
N+NiAbNcI3sdSZfG+6/IqFCPSo1EdnqzV6E+mWaPMDba1I0P7t0oLspPDmoBSc0RjLlWZZd5Ea6H
s8piXJVortIY872bI6Moj3dZZegBsnMLgMGFyeP/eX8zksHAuG5DbnP92aD60te7HChjPWaEW+6U
7qpXYaNsKfJfdPaNqbUf0c4HVgJxnSGlGYtByPqfKOFmxR9+c0v4C4mHCLvubVLUlGmVK3eDRSC0
WYtE3Pmv4X4TCqZLpBgLvY9OmjggGJdftI3yunPHrn+fFOPnzFkWhTXyb+jQGYbGdWSvoPgRfYt8
jkWNMgAAsO4sTv27coeSlis9vlAyx/vwufMpeEzUorj6VUpV2KgoppHAneyqHe4oraE+UqXyf4zW
P5ii6rWDVhNR7p6pKSqAqorl6YLUBPHERwBNJ6v+ifV6aLkFM0pFpaZGTqWXIL2RY+B77OMs+MEq
duzTFeDh+6uTG/ET6WDi2YBTkQlZthaq5frvy2eTtLpMqI9+zEP+xRosvu88tAHu4bjtW9QQNW+4
uIIW8k6ABQjNq5vCw+RxB8wpU4u7WQupuIKdYhprzSl1JS0K7m4FJSlTEzbLJpDHek197bSztpmU
Tr8+w0/3bmnEqTGDuQA5s7V+AZUCiGQeOCMk1KbKXX3HzpAcewNlvn8O8J0Ti/4VPRp19K2O3GI4
gAOo5A2ut3V12iHSHf6g6jnxM1n2Ai7zap6dg4ElMcu2Da6YvGLrhG+oS8ZX+UJvUPKrq52coWCY
YET/7b1m10pByAxBvuhVJHpFyHmES/YucaRaCAnSGB2X2Ifc9yIWgeWU2Qkn9vF6frAyzf3aPcyw
DerBq3JpmGU2HEyMk0Aa8PWQrMy25pjMC0Ol4CVPRzd6Gd+99zA+lXT1um6IDJZwXSeuW/uWKGP8
sPG3F8hJqUtFRCgi0NeaSm9VXQ2K+bkie+WO4Vn3lCBADAWK5wjFRhRb1POfP08oM+BiHT2eIpFz
Dsf3xfQOG4msGpvXbO6tjqNwAB8MgSZTchptXb7gd0nbJfCDXs9f+Mf8x7+Qw92xpzxtfuLv7/oZ
X4mP5nAR5OdjJ/Q0g1msaUi/84C2FlKJHzhpPa+JBp2GSVJUPCjhaafdarsHLLH6b9iJTGyAvk6F
+5O63cutgKRcTSjNMVHkgeyyGabI3SqlpfJ9L4xcv+dCgjV8g/r39+WxLz5vGmUJp17R5UEkZumE
pRhekPjn92kDce9DU1ptLMs+n88l0jM00d4mvat5Ru0hShO5AGn3oHQTMPg6RSmqF3o4rByZPWo3
s+y8j6utHe2gStoaSr4JWvkmrUzXDI/+NAW6ljRmOORsu3bdqEVhcRvDOJWsTiohKSKyKiJD5npN
0YA8e9VWjMMP15W91WFNDIOx0XyUSQXsR2IDGwlqhE5cdKxgSQLDivxZzTTgkzp9gDCEpog38yjv
VGUQ+UzWPticBj2DrYVW/hXVPqAPf4sZb8L0++Gyvi8yE+Bq5C8XAZJE1tzO3xzTEGOqlvpBwNjm
w89vMB2WrSYfvgOZA5tDykQm2iucRHyAXprRnHXKQtx7h0RkgcYYNbJq0ffpY0t59PPG696wp4Zd
QoNRAKk6KvrC4EPATGINzO39fLiDBlLmq6j/ingtf7ebpkvRC/VQI6neW92+fm9lx9xxppAOa8qK
ueV//0QdJ8N3NJ9586f20Z77Cmm6hKl2TvP6EjM1BSbCTuwTvpieOiQfYfP9M6gwvOo3pa/0A9pY
bhP79weKhhSRpEblbVXMHUo0J2deHtBUMwuFgqhSHNxyoWHre64m2C10qhqanrIu6R93wSY2J5/W
9FlAsvG1PAYcAzCILhLuRyceIyMxf1WrMTZf4i2E9jedDoBrVhHns+ckA8lGvdstyVTWwFqjECY0
UnfnARv4+7ESDLuV03WuOTRpb10EtALU83TE1mGNFzAMPxVeMVAZ4M5s0G0/gonb+2JNhoC/80Ny
K6s/JImmJcmgKcKx/y6p91/0AIKNv3YQgeadigFKq71eHG7tL+LleYwh8hHnh9STvhLPST6A1jW8
C2MWqDCj5XBuf7tZxfyi4ut00sN5CdJ87q1/U4Vzvk1KcwnZD7Ka4Dm4okXAzWA/dIlij8ck/dkw
dCWWAJro9qFVfF6S2hAbu+k1144OcTXB2CGIr3dFFdFVMD00xvTwmhPOcX9BYjOQLgR6yg/zEGIC
eMIKXYkt/kuUxJikmSBOHKIB6q8Zcou3apmDLvBxAmGkw4KyKYNSHVhEsXSQdhgRtI0RqX7YoleS
Z+mAmmbWdVet9K3p4Z/HjZO3PX+yGR6qZXhA3jD8BedLNiWtQKXv8A5kQ5cdEie9SGSFdunZ8tvY
0J9UHa3DR5YTFNJNONScsz+kBCnzC25FETo5BYVBjIx4V/DpnfmtopxIdCyNC+kRv5G6FiNEU6Od
T5lsAInx/o/+9jUWggB/sdlQ53cArD6NTEr++2ZXoQw30/tgdAajt3cixWjous1LQ+BjvSaRH8RE
hdpqhGXxQlgdI4zXMcMjnGIptI4qB2MLfsoRT9wwDdEwZtWgURxInuRkEYGM4QWYNUzcfoixqu3T
GqXuEwR8eDmLqcdsbLMGnY8dZfuc37Mjun63mENpayWhzNbnwhUXintOuYZnt3Fw/VfdyDfE2NOT
k9qr8FxsmkBPq4qAtrGJIrbiMy8xiw/aDh9jpK5BcGoms8iwmE81RipluU2qVyT1pj7gD6tUe3+C
ts9HyPuFnqV+UR3+Y/gmcnC7Unqu8avl89fch7po3j223qA9ryqsKOwM7zFhATFehTEO3Y9BcAZa
mk1bVS7kGERVF1Pkme3X8iHK7YuAooM8fMGK+oejKjSEwYPyt0eBRZKLdUIenMd0JyuZidVVD/IM
qf8adqS7jQMQw/IVQLbc4h6Rf94JKHqkJzZ8T49pXMHwpuys6wxMLQ6eN2ml4KeszNsP+HJ357Lw
JEf9H/Ku+9OQdUzf48v+R8H+bkkuNlPYyfmNrUFCwFsfRGoD/CXlgR2R9NxtQf7kaMxd0fRHtVg0
tmh97f/PufiEgVqE6UlJDvkiV+WisikPViYKnM01o+KDsvFLm6CE+BthkNmSxTjnZVlqGX6OaAxv
Kmv20Q3xxmM3f0W5sOApCWiLHV87W4Fye5819C9PhlKZFX2hSC/t0mco973a1XZcBoaP+OhSWuDW
9GZiccZeW3M2IigqL13DkhrY/wQusqejL/6Sk2nRKAbMjaqdUp+nEp5R8f+r1kdB8yClz9uNgyJw
q5SLFMJ+b41PhG+uaL1Q72YygCkIq8RBSFofgCysN5oAdm5ThPwsZzsHKYTQFX3VUnXBGl2iceRW
e1qF75DyFSXDIcAhgf7eyNaSY4VuSK3F0m41KwMk/fjXDfH9bBq0bsHwyQP+Geg0AtI4Utv6p6Nc
UU6cjXM2IPQq9KuUKWit9SB1VxRnI9WPFhQvLHt6hUox15i2g6uyZ/NowCGhvhzUwwTlzVu0X5pk
9k8QmBuY32PQzV7yoYuzXJ2eEV4ZjhmHDN7LfkG4PtY9wEO5+mQs0SVU7I+mqYXyxPu5myY4fCe2
xBD+SBBTM80+L3Xu4UNFv6YA/felb7/cFnXBxl2eqT2b9EJ5JRd38gMLNRgljwtGztb6uivOmg4N
smDDVGfrRYX9A+hwDDhEQnxPraC9hhDBtZwQKHccTAi0EUneIK+NGZc0N/KXIkVJMJxPpRWKjCkU
94V6tHbnezTPwszFkU9oL1OHHuFVltOOK6qh/lV/jW68RYluCG8u5CsZuM1U7WPXaIvHutVZ79ip
Q8CTkcVed5VQQpLL7yQkQHZSh67oQHeySK07eZiIgRqUgg903up0g5UKvW9WaRzo3RwVR6fXBKLR
qJhPsVWuNj/NPPYl06FtjI7kEsSzhkOw6rEHuLJQmpRFdlKLh1laPpaXeuLxhduR0yyN+b6sBRhL
lzzLOZja2CfsRih+q7s3RqnoSmwKHTucgJL+fcJfetxlb8SpkHOCNtebNSNAR3k6vjr1FKh1Lb0j
3+8Gip5Zeq+BfAqLNHtuJ8v3tHsutPLU7V897b/SAUyAHgTwmQt8zJ5RCMfe/f+ov/KBIEfhpjRU
acF7prVbgl8+2fW9ClcgZYrioH0xWyFGSKTjbttqsFT9kNf9gsoDYr8pVImN8u0QTJXMnD02PX43
sDezPJ5WS9MRFRCa1rQ6jI5HWr6/MH2dN7bjW7smfT0sPklXzFpV7hQAKOYl1gnd8o17eyBLa3Rw
psvceCYg52VYCqwNYtIciZzaj/adYidmCi+jPd9NyY6b/Yg0WhIQZpZ3byHnUwHon+AtDcPwNuHk
8KLZI8U56HkInUAV59hht6rst4xV50NqKqcu55l6dWYysLswZkqUgLimp4RAlEJuoDgcanKJGlyN
/AKYDGBLjbNgvCy21KvwYGEqUeji+HOBrkaAxHLhTKRqZtf1etaNCm3zEN2oS0pQCa9C8jdkHFBn
0Tn84nm6ZiIbOJ1F5jZ31wFl/lCUcW0aGoYOm45FwZMvL7dnfDCaFfPvfMsjoq1P7d9dBy53XKyJ
nrTqTfdHUzZOyWtkFZpIf3zOmRlVQyVPHmaPw4Yc3viTSuA2X45jZgxCUb2VIRqofkLpnIfIpDNs
4z4jHfF68RPhX+WewfePda8SKWBsCy6OFpRsDveLTvxqGLmcsUTktrh3ZQFWe64HKeJGtrcW8mQN
wy9dDbsTzQpecuo3AojNkTl6rWkPtU8SpiLs6Eaq4Rv1oAmbJfZ8ML7G7LJsf9hAkH9UbDpKKuR3
aZqsTv90GYiUxUxMyuBEeIgSoMsyJd+jjVi8+Ij4EFZuNYRQcVy6JHM5OXCPOhtg4kBlWjDsjarG
0vLIEzy+a29GdPuDLeNxzRULMeeR+iwNd0yNipFg1N/2yZC+5C74vwno7zDhM0MD4YiZcm59QnJQ
YBm5pzFlxCNPCkjtbI0Rj7eSuKMtlFDeQ7fzqzoXCFe8mltYjIkTxk6uYsqXGEGHFzwEf2nwhHPd
A3sjLMTMY7JSlQ9yanwEL6S+5UKtXs0GXAkNVAlWHj3JWpbDiSNkefx39mUOa5iaF2NQJ7bG4eyK
75fK8lPnLwGuvrVEguCDFGPfqyMqU2TwNsK7LLMWBOO670Uw826yD2cBdvddVklzuZHZRQ3P1RBD
q34t51Mweq8I95I2sg13vqNYAVYbeN1svOljs4LoK+eKMVNbFpEFKWDLA/7Ai3hfByH8Q3D5waxz
F57IdS8k5qVNzez45yyC2tejzY1OscuxcKEPMnBBKlQg9EYsdt88u6+alIaWRa3nbC3RytmQEk0P
roma/adW/8j9d5bQLORlH+S+QTxQfRdfPr7sUu2EvYeBsr7ytQkFC3ai4t4NNutqXwcNM4yQRwBc
/l6Xvkw6TMCYREvgcchF2lQtPz5M5RyzJrvQePmvmJjNgvokn/DF/8kvFLPRK3XLw12Q2qjyeo7D
TpSfFaqSQPlmnowe41XgoJ/oIjRfBdYWBYRV9C7aOK4MXwmVacIGAbSygqijWkzYkgTHyfcRvM4v
AzB5icDw5R1HzcyT+66nU/QkgnhQgxqNFmuKvtfzMpFDi2/FadEiSxnlgfQPg65DRoPQnMeXapeO
piCJkZXq+PB54YXACiRHJCGQA44MOpsygcbxv2A2SjpDMekm37uwsKkauz13Wfz/2Oiwj9GS1i7J
5MsjAKAEvbfqRF7RXt1bmRrWLSkb6cp0VkueGG6eu3ZGVTCtwTn/aTK/BF/Jb6wxIcbu+xnB6xCR
LAgbe+Zy/TzGbapkgiPXJmN2HQwmX//864i90kchLChmDc7xqamzRGXaREwROSu7mwV8PvKx4ZNW
06dgthmRtELKWe5OG1ogqO7B9yoSrCyRJ2/UJ0JKc+UWiJ0C6HTNN4MAjOXsx6mzc0rnP4srXEIi
69EzyqX669a0ZV603s37mu6KoSe6V4/ddGRRNFSaXSVtAzW+rVq9sMd00OK/QNGnkUSrBBZa06nD
5Unl0Ld0VJpXAVjmUlMqidx/RP3ce5CnRpMxOeM5oIRYtiHwmjzxf/eCpG+OD4aJUWshLmdL/ht8
nBeAQwUpSDMZBZPICH2Sp56r0S3cZSoRcL/6hFVd+Elm4Cf6jULi7nyg46kvkl0WARmYhI2fuDdj
6JFmMUAKsMYeDDCaZqJ2aRNW7fK5PsENiRvHPO4skmx9VOs1lu335wDxl4+A38EgQ1ELeODPNn7+
IguIaDOdv51xi6LG8DF1pAHlXkJRxdlB8NQOXgf3y8W66ExfE+mUUnJGG60tvly6hIscV9BAxLPI
cwZHxM6qGjX7zxr0io17itvRjtaVtEZpsitKgTWpRaTvp+uugsqSme5nX9Trh2EV9fTCxHqP+s8p
nCshh4HXf1pDiVpBs+pxPzZissGizwkAnMDdwOOTX1CxJf+NrbHxYwfrvsiSm3jX3Xs/fmRGR1J5
ZHc5K9rcH2la9/6B1UWN9P3wfEeMu1399+HCNhe4OJ6ZlL8+OKEal3AQ4ig2D4AMvKbz4MOSxH3v
GiCtH/9EFPYEA8Mm+Iq38tRqYP91miNLJBF9t4ZzaR0VC7JfYkA4UaWRA0/5KWvboIZvujxuNVII
R9aZeD32pPYWNhR2M/KU6TLdi/5vIQ4s7qLs/K/ruYUZWmt7DUI5L1DZa2kw98ZlHtlU0GbIgtMG
/N5aLZ3jIfzmP7VEPm/xrKEKzVs7Mo2JcSarFAsP0x33T4YY30t3LmVj+v6c5zaM5C/i8y+jAXI/
OV9NCXvMrbsdw+K5ZCKZC8wpHlxAyUSbMAjLJxjO8euCyOtxNihU5m6ZmjQWS4k/kRsFTKoazKnS
W12PwQvT7rnUoCZuFQ3ZA0XUfWqkZ9pqMqZp271sNDNJiaBBihWyzkViqY0ZpBb6aeenbffnb+zy
MHBmjfKjfKM9JZabnOCoRqjOZSpU8bT4WN7QgPTtWIIQF0fudyiuyjHn8F1I6lrpm0NEffp/qFZq
5tiJjGJstJXsJvTTh5IRiMnFn2Ftfrw/WfeOpkAHk2sDeerkSIeG7STTnt3zQ9LxiNN4pEOZ4Xx7
+ZOxvu3ULPRH964QnVcVoebrvUku1isOenAxN5RxjlRCHG4cAy/l4tNN83JdXGUYFdniMxwshLkA
eKBO2eo4fNILq0qNDZy00tGFIjFGTLHHNVkdptkoiQ39zTtqZPcWGw4SnwLCDAvzS/CV6UwSNodx
p2d+Z+LReSnCuyWbMSwjwmW/kJ+hOYeDmts1odto78YMnn8DtjR5rzcdQ1SelbL6bYs9xbSxGPJs
dl2dPHVIE58Z3sthCia1hhaZaQe3JPUYB2KPwTunFzFRDpRkzvybnTpgklkcXnuUBb1Rx6f1TQvb
9FqtkOhinH9+3j3zsJ5KtiLaOG55V7fmQVsrSHME+PWmBB9GRBaTQtfsD/c5GdxACw3nGkvIh7WB
YXNkBppj4nCT1ZPWvcoy90mCnGAaTgoYAGiqWk3hbjR5eN5LCAInv7GS9jS6gATPdOqEKSl4fHbo
1+WyMx+XIT/pK0Ykdyfa/r5AOwj/sB3HzUgHumz5FCuUMjUgBOjLSq22aCPEDoYLPrn7Mi9FtQjX
JwvdwOfk4nZ8qLA3e+4iYAduDmJj2RF19L0pg3oISsipl8Q8mnxmDntqKnIAcU7nWY3IGojqXJ1L
LIvwEnc0ya6ytfSqHWWXH3Z6IRhrXNlQ42oketPzkkQ6MFn1Evc3sxLNV9nCODtBbCsn6L+6niSr
ZM2LvI63LTD2ej7cAOsc/pxMM56yBxy4VUdbrAGVevruCzI3xicjPQr9J1brx5hKssbH8ZvVRc7j
mgOH+IswBJ3Oe9ERNN48C9lEXTcW3JHxoAD1Hn1NE5jpUZOqOmLlcH/6pjPEQypfukFUdKNrWYEZ
hcvQaZgojFU64MdTrC9LHK8q11woQhvRwRu++95mWmo42VEQhJSNsMF+pMot8M/mQ75Pbm7/klpN
VWOfPLtY6Xt99fn7B05eqU/A9fTI37HuLtdep2cswbc2zFek2Em98ExWXXebp+drUIBDlQVWQXrU
OY3/liQdnrltcYdd7hUpDtJXAF1C0XmskT4/hwpBgnJxHRPaaYHSwPuNyedpO4uEPsG20QGTiCiE
FK8idkIMa/nRs7WusPpfhk5zMbm8aFocWd5LL0pId/GRrTZTRCmn6nYZhNlNOp0yDb57a9kXvjtp
JWXGcnNZxz52pGfJCALcXeeMy/NUoEjeqRYQp9Ho+iPh9ZAAGuW+4IK+Ltzw2cKvtfU2hFSxhwO6
mVv44S2zrHNOLPbiv1rUsS3qCJY8qam/4dQlVgGrrp3F41Q8u7qkLd+hkIme9NIUrnHiglfn7c8t
pevq6SZXrNWcmv3HlQtea8KRUPtd3+M3o5gHbspfDQAVCAVdCvrDaADFKVXirMOMairWCUKiyLcS
LUUFEI8G2SxmiwkAuLEsj6CgSmChDpZNblvgOA8cc3IVSfUdOQOqAxNP+f1Ccqmp6sNKF9jWZWjv
umubFgv8PMoRcf5XxFLYEm2rkZcaSlEhNkJrn4zdnlJZQIhe231yJgQ79HK4A/CHQAX5nmL/HY2v
z5qahl0S0Y1I+rGWtDDbqY8OBQK2mV0jKOE6aRcgZBiamdG6kIHnw1HV2Jm3Liu4f5iciATIElVZ
ZVYhh2O2l9Jz8bU3u6JpNmbfJomdtHy7KWPfCA8GCIEHnPz2dWplaSmWd4YZKAWwOQR0waMNDDIx
tOnr06diV04k5zOqnw+jW9bvp0MjxD+/EAxsB4m1yEpebij9VaJYSptHXyDucaOK7JLpKXwvnNJy
OLDdcCv9gB9hY8XzeCL10Ww4Wv8VJdScrsWrxOBVyfJZuj5gDTuJSySL3DIS7H31EFXDtKeBxK4F
OIrqJS+DH9Bq/pJrg4KfhswyfCpcVxD21XiW0B/uNfMa1OTWCazUBWhjEH7Ekzov71/I5/irn+16
sNiTPjZaEugvFFOF9ZVHYD6NE0cuq4HNLai1zaADxxaqelYmVyzQya2B+f/+wkKIDSdPiQpgtmA0
zkJnihulhRNNZh5dZHQcJF2WRcWnUCVbSulXlAwDDbWetBd+LBaNyHcNBImXCuLzj2t0rFau9+QD
FkupZQUN2N2V4BPcQZK8/Ed0RPfuh9eFQYRBf1G3+or2CrkrsA6pOvqj78BdYF1ijoqcXK/qDmhS
enWaKR3qwaJK4juVY0geSIpO42h+mMYjvso7eRbtt6UwShTzVrg2r7CPNz2kjzP3Bif9b/7QrTCM
StLZ+7nFc3UTJR6jhxx2mOO0AScFSNqKppzxAKNiqRz4x9x209vBUNbbqwwD113Lq891gzK1T5kg
Zjx5d2r/O7J4IAmDVLMJ01DuYJ7+8U3uHlNEy++L0gGv6qSSTkjWh3pM6N4HgFBG4Ehpuff4Yj/y
85HkJh7bqMmP2JFzuAjTUh1AR8d61XDR3o0gGhWRIQRPxSt+atQe+nLk3ILNIvOzUxQ+6U5/qinn
DPyNxQBWbQoFNq9qXACvLnCiG/dWoHqYMMDEUzI6pdOpiwDc3JxmatLf7p1emk6Ik2oaXmqL1KFN
75A+TKAlzuamb3B1uAcyiGnZ0zsS6ACwxLirKKMbcOCGngxI1ao7Dbdw+wadLOUqWrtRHc4rgTcZ
kYsWdI2jTS4XHSb5gUfW+eA/+nxnrBqf/t5GABkR/LdYEtw42TQAve2sCeX944eyef1E/8Z/aehv
DBgrIZmanEJJwKRcunOtiDMibVP9t989FawP6AJXKeQdW2nT/KKCmGSu4VDB+Nq6kdVmvbAZU/UU
2IZhDjLSYRKXXej3Q1Fz7dZrOk0XtR5ae8XWtYu37+7rsGZ/FnJT15lhzMs4EFP08KhcGkcJki1/
UpHlSr80Gk+MTA8QEkRKSKib/hwR/+9Voi85y7kNro8iep0FaMp9WPwsw1KcqXBEKWBltUhMZCez
koaBa4qbTcJkAU1N0xftTf08nvqrRwgLtPh44hSiEUjqVdWal9MIcR1YWiyAGMAsLkAiB6H+uCok
T2L5H76c+kt3vCz+TZ61wWFqiQ/6uS8XjOo+mRMsLUEKhCotWshKzhRpKbAs4hgkcxR2LTw+ij1d
vs23Z5xNXANJ1NF2dGgHWqHBeyl1OhJjr37acyN0452pG7aldkVgETMX0NBEF60ugU45UrubegZ9
4q5/pGZvVw8+gUkN/DmWhdQn2qviA7xAcAI2Uy8JjBzUvJWuDSwEXr0GK7H3L9HV8W39yVaSVv/x
t0LL4scl50Sd0qx7ubReBwvuQcyWZQ8wz6o8YuDZpNxVY78ae8J7DLykR0PnJfUHzDc4tvc5e8EV
ozXfK3ZJSA/rnYjx9R3Tb027sOVf7izaGc4FghwVxb/fBY/s0uJu6YBS3vJbFoC9ziUkyFRJl5IF
T5igg/ugxUME+yIryXO59+ZTMHbebWf1D0EsRWED2IDdMAW41GG2H+yJj/e0HELmWiZMv+veydGK
wbQ9zxYgMN2PTXG10GD2y6okY+rfp9liuKMkH0QBU/2OdylNTkLT2XOGRzG/xehLsHJrNTkgykaD
Av2Q+5pUuv3K/ycfEx8BxGvXGEvNK31beY+3zCt1/+jG2OoQykcVeHNHqWCiB3qd8kWWAR5tH+nH
ijw1SuukyJTm71a2rUJXnElVuspwrA7UIL/7EtFOO7MmgIULATamIdAXKYsry+TAIBaA04P5odeU
D6Jl57lb0vUn40o408rCEABJkVMMooCktfi9R8AhW8+jKMXjiy8x7A30UfWqGb0UAepVjvr0ukG4
h56mQUO9rURXkIeGThbU2hOrSijPtKUZ6aW5/xcjGFo6JepR5T5dbyJZzgvEIJxJaCYhvp//9T6T
DzE7WZfpSIcwkHoK46eWw8nMpcwsHmtuc/EW3me0mBa62hOtRCEsWDdMJ+KgD5rPv2iKbQYwmcy6
La3IPAQeUu6lh8wIRRKnIcHeiB/P5BbZxyYp0DpoTNHBOiIYbdxvW6TtqcGgVidpNPdbik6orCgf
93t4YtBINjUn7txcYWGUeruwvC+gTiC49IDGbnWWVy4WFqwiQvsHG50nWtwOxrZA5lVqb/S+1W/7
o5YPcYTLre7rz6n4knRpv1wO/xzIAklO/iewyGqqzFmbR2g+LtWx0UjeKy2wYiMBfsJmlM0CDpdH
lTXtKgaN/7OsoMV5W2mxlkRSHUc0GxSThGr9WSvjAymobNqYFqikl2n/vwD9wD2ciOacDtmTxi7u
VJ0eZF1qR8h7DOOrWWZ2YpIAsgxUL7hMp/FXl5hM9tflqwfanw3rj2WyxJxtv7PLfwbSvxI8VfcM
GsLjs0DQUW+xd2yS2t7zotnRb+oHT3lHcoygeFjNCk5KDAaEqze72cDNI3ROge/tNFlfLnZmI213
DIjTZmRVxXsKM/kGoNEzM63SNEgt1YxSmvNdo8uc/P+wmxMprBr4GvWiZ4j2BKamdhqquqmtZfcv
3yP9Dhgvf/B7nznDIF3ihhVIAYPIuG8xTeCF4pZBTySzhuxwuB/akzJiPmeNQhPEu1nQCuMAC+Kz
WImHlEPbMz/9hM/pOFX++8CIVM60mPVJXAon+V+pMA1xpfh3c7NAzl7hMbKMd1aKzLJZJW5IwAUF
Xep25ixQg6JLJWiYorNPh21LCNH9lwVYmV8PK5cpcf20EbqhgMcYkJ6EMf5RUiJ7hCKwJChMu9Zd
piSrB8hmn2eLJe7CGGAC8GxJfiL2KZaLzwVF20o1ht8IcWS/lxCxHdq59ivkeqsLoqfjecr/rC6D
LsGWKNM4yIUAORWp8E3QkEawgHTP4+gM4rTUMjSJIizKCGZGW3/+yJc+5J8przFoz2FwHc44zGre
hxNbzsNtDUByknngoYBf2QXrGlFB52OoRgzgxR1YjRZiLfc3tNKFJ9JB8+c5I3tjBQ+bNJOnFYzP
DPiIZH3/PgCRtPpS90rbfaIWSDi37udx+6r8GL0GY0hqNW68RiuEMms1LuJbOJeZfYtBe9L9fciT
wnmQ64RH3zbWYVGrFxX83wL6P6T1WpNEP2THw7Rlzt/uQ1Qf2RlKUPnbhgnfskh10jx2lqaA51MH
d2ej2s9XURYkwss7XGJJzZGeM7p/mVKRkvSXcBEUePnnbGRuY19y1nsrOE5y6nEwPlwWN0A46y6v
JXPfTAFwX6iSXt8mhmhsB17DpHac9TkJzgLEfoQyVPrYk5L8xwH/SRBDFxcztWbc1XTxImtxF4D6
EymObTSPm5ucXHRucci9O5ZrkxMzGQY2l7dRfKUMLgiD0bGbvmM7lcW3ikJi5ZrVfdv6Iwd/Ihhr
q528Wvp1QHFbD77XJbxo8MkNHsFTVgrkAYPkZF87X5irAOMgcKo2Nen60Ww9Bs2GgL0H82HFCaqJ
WU0akeLuBHCEEYqI7voNmI7WEHsAra6GhHmAoN/fbVJR/U6fozdxslORhEedwDBspnEkXsDNecIc
HfEZMjUtLK1SKTEmdGCrne8vGv+nhmN6WDllyXDkS3QqSU2PDx57L+17T4RkNXNaEBVtY8QwIHVk
X9h3Mzjigc4BIafz866grjnVkWbmniezA7V7IW4xCVv+MjxtqMDrkppZ1aUXmQ/vLw1TjXJZIa+N
JaBCc0FTB2jT5fJiizAyxqoNYveWDm3RKbq1FSWipRO987bJ/xOnUBTmRotbVhmiOlI4w2VlvZ/X
vlXYGpxFcpkU2/mWKJyhfRReEqPQIVRJsmGmxTITjwCWQ6i6/1HA1KNVAwmD8eTOJBL83lLP/3JH
xnAgPtXWaByYmoFQ5vnzOqpTy8utpadZCIODQPd33tDLVxHSKhhCc2FybbFb/zdpubVzbitSCTnD
2Rs+Ck5/ShHRjbbl6o43yvR/4rOhgfRrUUtpSWoXLgDNgTEB6uyfgUY4/x56tqk3wxEoCbdEsTsI
aSZOtDQwFmZosumW0jddxfYXN3kJQDbF+RYzJp/MnbuKgEhH1f1GsFqtDBOhS73eMgGDwWsNy/EL
QLrOReH51bsSdfGosvCvOR6PmENTXSvHwS209h1Gz7n8omx8bUa84KBePKcImGgQDI79ucBGwH8N
H6O0xkpZTSTrJvArnEOR7ZeOwTq7EIEJ/Ee+vmj3s0g5+DWZW7erbvNT3COdDqzyacwVJ/IQIhds
h5AO6cBCxGa6z09GVC7kHoWTUw/GF/FzG9tDKv8vs1fMA/n0JPzH5LLhEhSzOY91I92uRgFqg/2V
ITC1WDU+yB1DjRIyCGsONzXc/4KLtj7419KmFSgV63OjhtT/b1dfX2F1LvVKK0zVBjrPcYrAV+UE
YV/OlH6a0lK5wx+UPruJTEd8k/lKBHkH7MFJ5o6Hh3JF/gbpP1NpkMLGpuIYE/bfHAbEdCuQ1mfs
TOI0BhAVMaG5lnwKoa2FN5g8dS3ygrVQ0GIaJNZaa8e93JiQF1mXgb1oSugbNZTu8gigFVq/E0u1
3zDq36dEp4LEi8iYtv5nKieVZ9ySEnZnluXH2INm52NsAC5UCRGUhFgoiUSU2sB55//RuTvcN3Id
8c+v6ZV8JX7eNsSaqwtpufV2Jl2+6Ffby2xp2tIerHfhmRAVER2C3IiPAwcMXUvuGiB7rQsYXnlE
7QeIS4A8KaxYFObdrPAJ4Rn9+lfcgOcnR1zLohJyNStNVzjsznrEeu6JAEr1rUJ9ymBIJgFpJVJY
NVWGlqWV34eWRkqx8m8Xv/Dg8vbRoMfose3oXpLZi5fjAKVZdm30oP/O+gy7FfZK9JL+nBFI3xpA
tHQADQMe9hKghv886ZHC8vrYpZmtydVKcffV2L47Oai6X4HVfVif8qtaUCfjb8fEaqjYo+nKG6bB
xtcD1dvX45W+r6pMj9h7NTfJiBkW4sXGTSMN13vHJCoqog+XS0c9Du7zEdY5fm2p9BrT0NTMm0ph
S1qAO3rfNXaTd09kYiLKqFMdmkEJAwdIxfYLWKU5En7lOvxX6AwgpxLRKpa8ni/DEvsnV6tWxleH
QrWiexT12cx36NI/oHOtgeCYDBxyxtovMBLmO1Us60GIdQOMPXHI8Qj/wzvvJQv2kSP6aVikEW+N
SklLltMu2iYKpdilB4/VxZzlMTFYSsjflfXGguE8p6QjODgbtWY52wAUKTuoAjw7O9DBNMwA3sAr
nGKPyhD3ZhdXQUelzspYpJnvt4Mv7dVyuT1Zx6FbYhZg3SyXuxPIFqs7KgDsRlFfksvRi/h3Mcz5
FnfIpA6rx+g0LWf7PPbSQuSObByw7PQKBpNgfQ0jZr9/eTSvysRVCoQA+Z8sGxNIRX5szLKzxyqa
045y9MFXFR2wPeEFwWO4m5HrX8p7JGzT8niMuigCvOGvpfebmAZFDDsna64jHYYjDZy6pCucVmDC
T33u5WbbSOwXXiEP38IxGJpXktKKihN0TgRg4/NiCih4sR4b+FGDx9oXTZD7K4f3/i2a4LNbi/9i
E35LZjravMumy89tcmk/2W60WiwD89r4qalkp3WR+dBNuQm+oKNeIZiRbnEuegtR768rl98aViwY
Na9tSIHMWr+TzyG6m3dsTC2SJ3NmYsioFaZRX6Gw8C9QW74WQK7dJEeoQxlSUjj8rpc4LmPfHyD+
3Tnizpg5fJPUokojYsz9VhYBz73JGzrxAXl+R9j4El53Uf4cS0x2SXtPIHWNPt3aj3eWFoZmfyg+
GkUf8ka2IJfx1ebhbE4kjVmaY1ei1xRLGmfHV8OPRNLkdoQNYKTR+eO1mm4znHxYd5Mw14ZClBLi
dEcgJKActGdx/APyNJ0cy8y9a43Awoy4XZGQNGoQzufsBzNScwa53wDMn3jJgv8cBCsowWh/w3bL
bsRX/ZsrfKMwCUBNcigJO5L03QwOHLFXZwjQsyenHujXof7ik0oRkf1UCCs/qdoouBaBNRQ5rFbp
xmucj6dMBTYL/p+mFMw9hBruanV4k0iNn7o1T4eIvXu2g8STj1o3UHXe2MxvzOjM4OghDbgVkxxU
1T94b596KTrW0k1XmmfB1BMJGAXcy/yVD2mlrJYhRa3If3sZt+zHvGybXbxfjX8nr7zNF2wFi1uT
mO3+ykLPwsjG3FluJ8t0u6QlNoyKONnvbIJ9HGIw9+hn75WMZIP3G2RlfsjBzpiDP7WPrX5fgqFt
kzShwvJMRsnGbBvPZr+ezVjmHwV0UMINZdjkgSJWLLSlOYf1400NlLdI+ku3r4YNDZ7+bfIToEwk
gt0Idxo1v/gk9MGXCut59PG7DqR45oo56rMzzonBwiRGWCUOSPtvrYgbDDDjvsuEvB4hLkmr+d2q
hgKlt++zTgdanbqpdYf8VcqEU8scR5mx6B2hhY2inDg3Xnjgk0YjUzoPNASXJ0Wi7UovZtPVhNOX
Nw1qQkdKxY2KCt68h2fQdMSuGdMse4nmTqckT1dQ7nfHZoSkLjUv/Zq5gCkw01wkU+fii8VfHpZ/
OGaFVaZukmVr6NayRtIQqymx2+fX4/srHjNjk02Ks3o2kw+XdycBMsHV8FuxluS1CKzP3YOHAWRI
8OmemorRTGj1uezKEANgYW8Uttv3YTPfKONEMADM4caOGSsir7tEh5HqWtEFpSI0ODcPPyB+d/zh
FKt14QfkvEsDwrs/UEsJ1wWod5Xt0ENp//Z5MH/ajN1TnISWge9VOlBbu31SMKv97w7ElyYyOtEX
T9nBGOc3vniZB7a71PiHzMjJ0EYusIKyViwJ6QCfltZGyPynXYV6hk4ajuPP2PnWlWK8/ETgpXpz
yLH5bAy2kvIKOF7iQZwS3qh09X8akcnyEoadq+o3ciFLGl8KM76ahY5nNdUsHNE5zqE5l3vq/xMb
jIcsHrF4smvmEJipQInokhjx5F5S/RMD5sJm1my1CM7ln0QX8p4TaoAqDv3ch3K7IQFsjGvRZGNu
RrEslKQM6uVt0bZwz4sxcelWRSBQUAmA9qZhgLLHmh20pT9MDCYmWaIafLlaCUNmeqLXmclpa0in
k8i+/FG5AJgINujTQKcG/0QBaGocrekgrhKqtV2FPIJreL1rr7oBGHbaiTlQPurCJqUrdjlPK31O
XKnOAJMo/4GA/rSrw+MAQ5O65WaC7/wCpDqbD8cAQ8TlJXBnWF/hkKlGgrIWnNYN3j+tXSahzh3K
3J9HK2CZf0UrtZWtPdxv029wa5A1GfKHaUgJGYQxhdTo5jP8z6lB+36KBL6LZSdYxErr8/to5GkZ
EmVQFXVezRPc8UL6fhDutrVbmBUXmeWwkpzdYRc2pWr/zwADL75+D/VFflQpIiTOcRMoOwnAdtFr
RSCMEzGtZf4JgeD1xY2IDzOico/IDq9/Ej0XvTy0PWwmiORswHE+p2iefVEs5Todr5U2wT8GlGyh
xNWItE0yNEAs6xvc+NeYljGZe+hhs+YBWzXEDGmU3wz/MODFPp4efOsBoZEmHlxlqyWapByOSMym
+p+3AcC6hfR+H5Un+jiAoAKpxazneaXrgUxTUSIwGP8m6a3WU7eFhVziDL/BUF6QnmM9rE30ETjO
nxhiyC4eQAnIlY+w0vSbY61+ftMHtYNSIsoZZ3shV135OkyEj6JGv5cbcDR655edGqnFdK8JWwMz
RNzp9+7Plg3wJ7UkK5F/s+bRpwZP0Jy1y1pAd7r65MP368nSHU6V4hazlTySPRbT8fivXgxCXpWb
HMONzuqrPgBgD7bU9HiGwN6HLTMQEUHs/vRYt69Ecp11+8pE2pdvpAsQrKu7p0X1bdKOCK7UPbDM
5yfTTiV0kcYyjvnGLbhDJDaYeSCWS5gycxuWeQZR+BgNKh64Nb2cALzc6uHdWfPdgzlOxkSSZJSb
di4H82ES8emKcQjrf0UWvasjDS7QgvF0J/RFz8vbOjlXXDPKyZDnY6xCHTbQxPNXsxklszJrivN8
7JKe47zF5trg8SVL6OufpF7nrfVlBUQ2q7ic6zJ4B7I43tJZ4VhfRLIqZnuydMmnF3NyAY71oZpi
QspK2KQS7gRZ+dyN4ve/NZr9PyHBc7VRrRykVZ/JeBH7NFRc1Ovj+pzd+rRdkRPRRV1fJAdr9W6R
S+m1TCvHEZQoiaTq/9QzLkIVRI+MH8/rTQDIMKxvamkm9KZxtW8Rt4GjRwhxrn0QM+LGTz7TNb2K
YAF14hKK4ajAzLeEIh9tpsidE70D8lIOIDzQN+CQTlkRj/k5j4dVhWi/PaodY1TK+IfK/jHTOmAq
SULRt2SwImEpfaE2RR8hbX4+2tDQk/5Jm9gDtXioAQIK19zFAQ2n3BaXcrMg7Z/zXAAO8rtBZ3h6
GFGlYW4Bj4EN5J2mEvFHO2B8qbFu+goE5EQosM8VQUDMXXGZUSmUKAEAk3JFv8Jeq5uVh2OXnTgC
SeruTri+6yj90emCiVgDkdenQ/0OCwOeWKVeXypHYKx41EBf6cy/XhAfD/qH65dQpw/KkPn3AGek
/4LoL8oIDJx0SVuLNurDQinDrzxCvedGKhgBpbK1dwwqjlnuzrMiQ3ksMmWWXrjjckaRCwsX/Ap6
jEg5Epswl9QHgnLIRr7UYfAjRsc3w72WdzV5b5rdtUqVCerLvVJnz9yZE0rn+1Ulag/nb0fkDN4W
tGyKHGTvkx3p9Zj+DTyoLwIMaLtNc8jg1pmdgmFAJLZeagTGBtSIViHHlZ48bQFYnT52RkN2k37/
zE8yXwc1zWpnHw/xe0M2kTh8W0VDVdoLbpUkB63yXQ5VsHJFC/t3QiPwgj7AD1LoNqXl3H/HRdMY
TnFMHEoYkb+cCFTo6yRuA2SQiSGkKDVpOFJ+ch9M/ERjiu5fJJmW97OyysEszSoX034khRRFcK08
TKuYYuGOOKnFN6WAvBncMgh3+8JL+u+jE5Ao68HTe8/p6wjT8VY3jRCvjNI4L911isulUFpaZPFA
1VmdqM++HnbvlL/h7cm+ecl54evzeCJQpFQiP7M8ChziqeZRc92uCvnzlWCAZBvXnvwOkdfLeYlI
3ylpKT7DnYNIhYtiEF2sK5D4POIf6IOhdkFDLKwOeZrRQu3Mz0A/zbZaku/Nww6O/hgDpCVcRabs
+BubOU3V+mksG9MNHFCQ0AFOO8Wk4QUPNZMgI5Htur6haTh7S4P3Mw2tMduPmGg1TN++nGkdQ/cB
4OMFJWE1k4Bkr5SipZc9T7334SV4v0wGK2ACF42O9WA4KkrtYXzS+G5czhLnhhZVtKN+Jz6dI1ny
Ak3rEG7xNjeWeSYTORoHaXrcvpxfgJAS8yZvQocXsh1lSRUXiHLLR8jdMkfEA/T9Juw/d/YNeNCA
cZUHL8jZSacXYZnyu3iBOS0iPYVUWV7PnapQzaqQuSURVV2+9vSTIO+wiqIwxUV1KvSia4FCiFDa
SvQmLbJhygz0uP0MT4v0MZAuHhcHUudmduy/V1aOpJAFIYot2YSzmdsyjge6KMaEh0LoQsqiUsOa
kS05JqvQ+itM7UkKvtUW6K6FIRrZ0+qNSUmBeMGJC3DT3xVQQ6kKMdKFQORUhX+P2hqFzGHJCYxr
c+m2hly1ja9Bqck+xuzEZzVIQWZa5anIEEcq/o3eUAHJH1G0eLO6tAWZ1sQybJzQlvcsgzyWWj7z
KIgaVUlmCpRuWqquyfYlAl+BxMKo5Ngza+pGcd8o+DBiDQXSeX04i+WPVNUdfNwBzvoNLExrVuC5
lO0Et4/fz1Kw1OExCed2IayKHrOoU08WrDOiJTL7Q5TSgyEk9ecHqNGTbE8uLMW1nUptb6p+CkFh
hXkwpCOrDnoxqOb0MIv6NywaVXpP+B90N+fEjQDw5aHQxwjjETa9twjskR2dgBxksQF4M4rELOZr
vmayRY4yl4ndtoX0LRAAfVn9bQa7kU2YEYtb3pEJfXgGwA0EhqGxI3mXrG4ugaYpBlbJwxoqomVn
tI3IETQEoUS/dyX3ehgqKUwuX+jz2SkozX0JVIEsyJj5dgUIzHR1BW4awqbbgksu8ULSy8f3tPPY
Sxym1w97kvQaIkCeiCRmzQoJiPxRH3+q+NPfDGwz4CSGZ+j0ohBsIlcopOnifroA2fYkBk2Xg7qc
rI2XVitFBLWwqkyX2sM/UfsNAcgncu4QdK++iaVKO+LItVg5T/XLx3/aK1T7SxQCsBZ/6FykA0NG
bw6iwGnlQJUrAIROEvnI3KxVn6LnUtU3LEF8p5YJjwOrSY6I/bh0e8A9VcCCi0NguOtF8KIxDk1/
D9q7cvaVbEiBByEoI/eXHaeM4sScLPz6UeLgRY2MxhWrIYsyH+uiMg4teVrcTwsR3bXYZfpfRW+o
M6BaW8h/IU3XHc0p/xoyWr7QgGMm8UaXLE6bQjCoW2cHBBtjk3dUvBHNX/eMc6Be6gnTorY6wov/
Or/c6MKjqj7ZFbc5VbYx6DStfhsQHQZqwfKgQTDy01g+/qNqp0dhFc6zr1DwcHYAsqwu7IyrHU9S
J2mPsvddVcVNgqumEjEWTKwE2Tx1y1djSDx0VTY0UNy1yEXUMI36iQnqD0rDeqXuSunlbhFMi8KA
ntm90r1rNjY2EeY0ZIj7m3FMTj/aUSAYiA+uDW36Ueotq9BhXFN+Uq7jbJI2H3qrIuw1FoXY11Po
YrNezRm4g+dNYtdxNu7Ppm45PBW9SbTUZUXFPH4d9wn4M6XMPs4XZeeXf4PC4E1vCdo/vpJTfcwZ
yzaga9HulvMn73nkodFDWbJl9V8UaFUEaB/PgONT+XZekDDkyRfPpJhofRBZapPVRAPTxl8zSUAm
mqDBBscB32Y82h+6qRZCz9qQfkiuNc8s0qFoAs4DdV7RdmGIZs7W+GUxfxMRGoRuGvF9hslaELBJ
JtmGaLo8b/U+wjyUWjemQSBmJdcDsC6zNDA5diL+Ut40S0zjEQsytp0SphmLFbVPh8t3K81MnxX0
0xNuN7CjkPOqS8+wyFDkrAJ0JxlDQruSP4XW2LYfwYYt/w/yCDRaZaVG+nhncASH3o+oXRcXTpd0
dqwhx4UzSIyg3FbVh6vF46OIPT6aWixWH5M7NUNBhBzIHU3/OGfUG0JU4Kyhh4a1ffBoO7aItbvM
9Z6E1lWlq+bkV8zamQ4PrBZOaENbUrOmKVln+iHUEkfq1H6Y7LAXgOuTMcC0hQYLCrE4AEynGmRW
WepLsJ7vHCGzxrB4DXNhvUFl6mZOwBex+5T7M0qf+fExtJtyF7HgwVmcoDQK+efXKYRDyv5fB8G/
N9K5fWfhNsqjPbK9Y4y2w9IGlwEibLGgBDmJ1DAqSG0ErMK4c0ALe1OXt5rHT3kZk/eJ2K+TCP8F
rhSMncUkmD5K4PlBzcozvA/p0LPRP6EuVsHRqRKMgDWF2vQdQMWLbV/SYz7ncqcQ4mPRAo/PkVF3
2DX1aQF+yPKtxBr4ty1e9cGUEik9QJrHX00b3RDblV6sRdlXMwd6aJSq3auYujpliuzl91u+Ug6g
vhDdjj59/0mt9vkFueW5XeuLIDPmYr1ftPZf5G6etln5pDx77OaAYeFSzjqotbo99e89VyEXyPkB
9oIeJlNfKd07BJV/q2E+j/ryq0z0suJAu41xohspkvkPlZbD8n1okbSSjr1ZXH9xU1kOvD8h/J9K
/E21ttuYYLNIj4TfUSWAw2XzZxP8j3XzBlfTFEjCa26YJhyH8Sx8dRfQ31Tz6FH52pidh7jHyti6
kJ2TMVo4Z2B0Hq0RvkDch8FmIel6uhb+uotSbWydVSIK1kNWdzyqvEN58vUis7F0iA4hd0TVLqoK
/rj35Tfsw2+c8TUBIK4p/rPe9kGNQr11i2TMFsXLHZZYn+YpXASjJzBUlH09d2qotZ0f2b2hWo1A
FP+OXCFp8IYdQbvxMO6cVTGTqvSGHSNC9d0E4vTZD1ZDYpiPddfJEXtq25NSm5NTBLNXM49fiZ7U
35FLyBVQNQ5A6Qto1rGduITYhRA/5urh4Qyk2d3hzoMJESM0nQUL+BSrYBgrPSGPaN9DSKTPfqvJ
2s1d6kAPLFqbMIeaOd4JkaA3ZOI9XgHRs4PA0oL5wzuhGSQgwPVfoDjJ4uCgdMXbWRmgeDEiBTvX
+UqCNKSV7ijIqqXz1ltOORTZJoJQB/0VUb/3JlXWx2nN/2NeIzYJA4fz+rumAGh59i9OAtYZXJc8
CYv/dCD3u/F708kInrQDA31iiLd0P/cCLy44WuwPvJOXSA4/V0uq4kAp5Se90/tkoNfYB75hMtOJ
oTx7fYse22ADPaNBt4KrWE3kGpp/5LBLP/2wlUNh0dCnZmV03WkyWz5Vn7qbAhe+HsnrXCNHlUEV
lRB6s34E3Mdn3KRFprN9+5N5P0CaSteeBBa1Rn+D7su20NNckLT3z2tO/CV9AiJNFkutkpDh9jyg
9xCHeStdK2G+mmBz6wa4pQWl6FockJ6aazOa/cFOVmcSRRW4fdKOw6PyD5g+1NdIYZOpDrQ0p10c
BsgCAEEOmV125Sop/wrCROlSDvWBJ7KvlzDPAI5s+xrRlwdJbMMhfdNxEgANSVa7kFjDpdRat/BX
v6s8+uTeFCbJHG85BOWrO9rZD3mD5TjpKu5oBqYPduDfmcVE5D3pBxtA6Kpt1YK5oAXgKBgrxbpK
P+8v+OolMq+1krly0f9LZGZ9PQdJmQtGDF3ajMIRT7qEjG42srgq9zswCnDdtVZrplZnlE67kfBj
5JEw3imxkrE7jU9bwgXuPxNeAR91Mg7MS/LfIwx36Ey8D6C+QDboWznojuqobrSh4wZaKjVOmQcQ
sMuLH3+IjHy8feouu115ohg2UrUO7Jmtu97b4ODdgLg9OyXa0PL9jVeq5PNRx7UExUyzkkp92Jmc
oqIyrLqM1lopKi6w2BYWTQfOVsify1NTvlvL10iz36mp/o23KsqssDVgFWnUBUOL7IIYl605h/oB
/Dtg8AYeHILE+e/ArH0eLnuRNJ//26aLSexdh49BLUFSBEYllQulCyNoIIidiZACb+rQ+b1BJl98
fu8kUJEXLAkLFnG2Noy+diWNk6dXeJDS5lf8PQoVydkYN3N4pcE0U2CuHkf80KziiLyuCebF9wJV
PoEsVDE+JaSo5kH7UQ1okh88PQzPpZMdO8Eg0RS7o52N1bvsW2fRENTpVJ0FVvLjH1TptnA+iFs2
r6EVJiAznx/uBCUkn/EiKwmADSvr7ar9I6m9dZK7WGtFEy9mn9mQZRptoyKZnm5niFtDVB9GKLCb
YlhObNRTxPmPdlvNxWabgSyxJxAebK/nfaj8uMl6Pr43oZfLPGaGYgvW+Oes3XgJiMWjtJqMBlcR
bQVekA9dCO0ltIabsa7Ksiv651cQZ3moPfDoMSSnFselhlAj93V/g7ccQyZ0zPVnmlKXrj42SBZx
6Ds0aWP8jU+IKuiFLPhWtOXOBlwtLqUn4iJbZRkgkcn0Bb4kRkj56A/ir9mP1ahE/YiQcSPJpbYN
FEz4MzSIyWISi/uRhtLdkz8+Ei+NXhmL36yd0j1X4Oke2MapQjj5fQcKLkHLu8BgPMDy996Uzl/P
ti6UD3mnmw9MhCGKf6UTvUTngUESB1n1TGt1rh8hj7+2FUP1996+ECilJMRq9l+hZxa3WRCGBtHB
ASs/4oNVeReOVbJSXMHAA7z6FyJiwfhUvK7ywO9zbVMvMEfXZywnf8KdrkRA18JNVc6tBucnMSi2
Q0Bo84cKks9ZuHDYAwZTPQSIp2C2OGcseuNyBrzhUIvV8nyoAnaiprZ1zTrTcdgT5bkN/sOUflkh
iMKKYfrUwFBUXx8Us06XzZWjmmppRH06j7oVmu6qms2VgZGqa6W2QQJ8RWbMRFUpgi9U0QHfH07U
XugRM7eQYtPf7+ugTX8HLhxY77Zre3k3K7PrfaXRPK0x5CjISDh6kinkFHbXmv1DVScSUiruHOgf
AKyj0tm1VqakSYRy/y27ytrriptJbnnS8/Y/fkpFu26p/aGv1XReqV7C0Z6qVYt5qjFJY6RsUq5m
RLrZDK7Ojr06nUnFZizceq5pQ6BCp8a018vMJM7hh4ulwbVCfsFmh+aoymgYnN+ghT/74W69qLlQ
Z+0Ig3qX+wxA74POJIjk/RnZazDu7t3AoyxXZD5afhxDJYjWWOZY4GOMmZdbNCuSFERBFBGEOHuI
oMywksmEWJ/Yr8eeaO7pMjIvt7EPXNcx5Vc+ZySRaVWXbdkpiUHxNVu7dDs8eYtMclq2wfoFnO54
KOphFWXmUdkXPRuFK/tpZ2IVcP2juRNrqgLBTJlepV+OVkpQoXjtwPyz2ulixIeFLxjvu6SNJfjI
kIE8WEZVarj7rUAEUbsErE+bfbOL/fZC7vfb0X6/wfp7Q3b+rOGvVafEX3e3P7iAii3pw3OYE881
uegxLl/5wHsvz6v3ptuaCfSJdVG/BURoomA42gH9UqCtQR6XcBNyei9ba9yoLin/ZZ7KjOI0VbWH
jevIt50pX6Q6BiwJmeFl/AkoBHkPUSDBJakIviqOHBfrBdiO63aKPl9pu+I/E36aJeAcmhth/aWt
Bw9ldVyZ72qjWMI9DKfdZU2UhLSQJC+5LFwvm8a/uaWcHZTGI7UtvyhW8XEALiQC3t2OuGWenmaQ
71SQn4zjUjNJSEKIP5B8nRiFCA8Z6HOiZq6HSyHkL2u/Tlz2VatcZn6lc5D3wqyRAdEui3OnD1ON
nK4rNRc/kX8TxLRfsJVkz0vMiqcecGAdUpdDhkJHiyiiGjIAxIRiE61GcLUqw2GFKvgHXKmjIl+7
Ixg2LAjasjB3lMLq4XcqDpSqdLuPUCizuINtOEM0NNYpRUpCJ2t0FGE6M2e1QrlJC4yyw0NGUIlZ
Pgy/kuv0aZQpWUX6JtjlBvLJ4ZeEH9v01134e73SyZPkckJgetBb4e4KJq473Jj132ratS5YHtwX
KlPsJddDqeO7JZkLqBUM+2ptyekpWtwSV70w0WrR1Uuo9kZTVe4GhsJnUegS5MTO9jrXuEvsd+k5
Kk6qaIpOth72POv79L7epKB1NovYBDriyWMt8KzEZxo/zxikfkwliJYUlJOSpt9AmHoyE1s6bvYH
l2+h/m9xzMr/FLuRjIqj3zkZwkvBBCxblEVDcKCQMgbih0n5yBUJ/5jJuajiv41f9XtBtBqNBCbI
g1eZXRUIaicG3qBPQArUlCKlOPylDis6G+cdL4FyNQWC1Lyb6JUExzHP+N52w36HMV3oXBGCsf5o
a7iVzPrZr0+zSjf6hJ/vzd6fI2wFQ01hN+pdA9ZSWTjhtp1+QOCZ+f9HLgQ2f9fSbCOoOenfokLB
7NKa0d6Rs8xn29UiJtZE+V90oWon9p+BTKpdrmiW8rEqxCJqeJ0jQSnjAmx0zFbdIkDPfmvLXUDe
15PpoJ2OFRTRS+ZCchRL9JszMS9s84vREEI64DAn5OFfZTOCv46mEXmGimv8szThJfdHqFm9KiV5
NGkoYkfwCTtK5BQpyq1L9VtTCDzVkVP3LKUIcpAYIST1aHaONVxltNZ8b5Y2orWqX7v2VEJafFzR
H/oU0XLvIwN1LyUyxgrMbHOZ4sD8UxU97Lk62SJjoNGaiE+0VsfQZR0PWU8NMH0qS0L7GORlfcH1
lzsuZybC1FvfjCiXIPS6/G+RZOHdLRc6OE+OG4AjCsH5p1YIghhtZKmDLQtdfRwPq8tqjfsVWioc
sNCFBPW0Ry8xY3NUNfATO4tLF2Znn9wbnaQxputx+A40V28yMq+wRuFvIP4L9V0IzpbfLWqjBf5K
ksMZnOCIGZnjK6aA9xiLqlZjW65ySQVoHzrA6rH92n41OvBjApzO/DnPd8P3nW1j+Bjoz4EqGifD
FouGwvCybierbsm1QzbKe5HAjoI6F8Jq7cXVESzBo7v6yZ0GO8KRMXF7DiHH9VsvZIrhr37GOrSN
J/vckZMOj6T21SHKXaC+76J8ac2K4GW+pmIrLCgcuAwPHvVAYc3nkJvjzD9cf4a315GoFmNbk1kB
5UjXrhLt1Lk0nywnD1ztmFKvpl54+3dR9k8S6oohfDY5fBos/hWyu33J8WvQe/Hv4mMA3XTmN4P/
Sx13lzFmRkRzm5NHMwUcwR5hardSNhcWMkTjqXeXwTpu2jWuk3Xn0thZ0xnzET148AHjoJ3h+nzU
8pszQ+L4ptcxPUA2SpL+wYmMl6+nUQV4enTmCT3U0Sd9AT7ch+efuulSHuwYbQo1rSol2b56Kn9l
adY4jX+cWMzkzvLmyiSfQ7Fg3MCvE6mDJ8RJ6hfX/WWAlpnbpGhFBidc4Up67Y1Ov0SFpImM+jM1
mcxWbjmbopq4kPkDCOHMFl/mK3NIV91T1fy/e3aESCjyaVw6tVjLLz+BGzm4E4rq2YWCCYtQiQNF
PsKx8m2O0APas1KnI+wxZzYM/784OxwO1OCRwIEMZnwTr9B0OFazcJCJICHrYnVu7KNdaHcpcPv4
BTWM3cGOWteXGSOeRxGwFJZEvFzLDsVoGxd9PWmft3XfF6yVXd1wShIlHDK1LfQl/gXcprSshBMI
IS7OVuO3MQg0kQVx/nOo32DhZAL5llXCkdJ3VFfX+Mrb+yzZbjC/BjztLpgRvJf4/jXRYwC+aUmt
NtJhfKfsj38/R/Qdww4pxJN1D8Q+0ckR4aSQwp06UiTHPMj6OCXacp89Esw5H++xxG724Eh/hi6L
OcZGiVtA5cQaeyNrQRkqMf7oB2iWm4bqjNQCM1uoA2eV6OtTm6NEtQKo3AiGZMIekdfh+xCII3LE
vyLLXXgNyvbwQ3X0+KSgo5FoFcIOpJrC+KdmAMQlXYTeWjGg7Yv5MsWMW+i9/3hJwEdbbAPKpCuu
eVATQWsR7Nn/lX4u3zSgj+ZOIOHkpSFEtCsi88FcApQscV4+0m4yc575d2Kq1ZncMMyz9HlvfGQa
FfD8yZVFRKEQjTiZgKr+CsfaU3Ai+HhthsFhgMEM36xrUzL3cDkM1LpvET1j28FQ+tgQbkRZ8wL0
JbWuT6f89581ffSAu0W8HQEhATU7jSSNOPNQAC75j0FnWwKA1pQn3V0GCg9xC5YsUGI+VCiY/p7S
5OQ8LmkGP5bGnc1BB7gW7SQhWNgpwXGYYj5GBwW37qdT5g8wFSOfHMh1oZSzkrYp/GE85DpoFT9a
fd8PX5fa+9uQ8l2ZghN77FKxJsEe9zY39d8gOdiy5XiLgmZrcF6Ot+V6jjmZZgQ/Wk+18hOIyG9i
W++WWdP1YOxeIaIDwlrNO8vB1yzZJlA6+6fcnULHGLhcPYpMRm4DIj6QUEnHAmvpZqC3H78uoQP0
vTjzqYI53CvL2KaUpgyCXPRMHXr1DGv4aP8drNRGArYLOYdn5OO1Urum2zdagE4xjFcvG1jAexTX
bc1M8Rj50ZI5ezcTSanrzBB3mlCRWYI2eOuG+9T/Cq3eDVQ8x29GUkeqgIyjhIc/Vo26och+3ZuB
qJ+t6VhNTZilxtzGwWRFN+ezdPuHcqDSDNp72kkr9hvravbs1oz9zpUXLFsa89kDB9NraSNVXGPw
Tz2Xb9JwC9OVpqRDxAzQBX+USJdfzrKWOfrZwxdSYlugyLF0PVVm0j/pRu3RC/Qh3C89eYXeU6gR
WBOfTGovQJ52Q0jbxj5qSp0yluT/vKyuaWAMV9NsUz92wYbQlKZAIZB0ssQZd1SNkCSQkQe/2enA
DdXav9aYKyiH22w52VCQPaWJtf6T/5u/68w5tLzVkX4LurEKAjfParQevp4vUtltcE1ze9jUSZMQ
qN2gbgulWsUS/5WA+Tdn6UJtK3xZA2eowOQpT2tokjBv4noxSL1WAB4GTOUGpKUBhAgbCGNIkb2m
9ffxVv+vXDiikIliR1+sG8H0y20i7DPPdxoUdRZlYZloBIeOxCYLD/kjfVbN4JFG6+Rbh2rfBYTp
NaQ1MriuTqJckKSJiJAwAm3RVRhEBCQ00oHRhfubGIiXzMRs6wk0MFnOOcEo5k66MzZvCLfUcI+H
yURv0tU150zEfDP0iHeHv6B3wCSNDQ0aihKAiI+XofayUGh9gPQ/Pd/9mknjqBn3LZLAuscnj7mk
CvODqcitaAifFl5hOvsb2S5MiaDH6Zi9DQGLDU8a8LFnWMBomtW18IUm6zehP4NGh9MpIKDL9MwO
yUYWX2Cw36sNFB+Gm5FqQ1Re+3U5lcYLX1wCUbd8d8zaBsAko5dppRQXt+5UUZX8+0SSDiU1Y+5a
m+erLNU/aXYb1iLzCMxqXgSjg8u6OAokcnL4HWOrB4+4BYXfSbjH+GobPxoeh67irqJMB5GlOZUR
xmWh7LyOyRWgoAb7L7gyCLJ4uPgPLF/Qn01esAzYIADD10E0Qh2a4i1B+HFJi5Nyg2LoQjTdDM3m
nrmknFl8EHoQUPt7bc5tc4uzz4q6LupjSzz2i8WIYtfKT+lgMp9UiHXu1kiWZhRyi9yYNwuFc0Yk
dnwiOdaOYF9ZtjZUSQyZY3y3qVmvAsZJBYStxBRHsZYVsIjo/DPnqDUUsqx3F0xzLzwijHZBDVUt
FUuWlTM589ncW8z/O1uHpDEH/Q91YU0oAwlsLCNLmi7pcXQpPyCvN8KBCzXdnmdVYfn320F4m2Gk
FM7wsSF1gOqBYCXrG5vJKayR7y1ELV2/oX3ylZle4aq2XhUDOZEd2ksEgk3IxIjNM6XR56n3G+FV
0RBAggKW5/NmFrypiqwFeEW9rUi0k7NK5pRPLOO/s6KNoFV4E3wrPMsVZai4ncO24j7tLvvfb7K0
jvB/u7ezKbhhOKDZg173/G8gVylB7/ycrq19/G82itl7YH9iGBygHrL/jXcU+RU3G5oAs4t/6/O1
xkR8aw/T7MCaVNKvyzHCbZEF2QXj5DZS6B96Mb6+Ht8cJKgYmR2/oq9PyaOEiXvkvAuFuHoQjSyX
17pLHlnfphiXHDRQWsQaGCYiPEcBMrVPKUlnVfOEobwYxmlWyINE6OZ9n/hVPkgJ09YAaQAqow2r
5ZnkUYfkDmVRbFRuJFDl0sUFDdDRRdGbu2nOVB3ejVKTmRHxJvMIhPITOFNA2kphQQB1a6m4hGiX
gu0EuoNAf+Y274OJDqy1qEGmBIAAt4swuOFK9LkFAqr60v2r3DVg4Z5hJxeuf+M0wNbfudEPwJfQ
jF5DRm5KFp78gaUyUK2i+Da+Rywzm/T+oCz1O7QRsg0jY1CH/rSFM2H9x1xmJD1kr08OuLdm5bU1
RSdJ/3w1KRfvAH06yJ33QFRM4TgmaIDheryYjTzY5iFaiml5mPuMy2u2O63MXgJTECeAtHNdY4un
ekUETy/hceUN3aqgpROm788lAbtiCA1o2fsX+TXffBldqYRZx3/yt2+tn+IlClLmLCD3hN9jifEV
xW4rg9ZNz5srK7e+s0GffxeTzNRZx0fVh2GkXP90zePPIscGClSa2Fr01rt7Ol7kJVN8g7BJjHUZ
edGEtC4HvDm0AKqcCPI4L9yIr4FwmLPklYZCl1o+Gvx+1lyADJ6tZyCSVWgDCCYBroMrZzDEx3lB
LpCCtYsWB64iguQmxAtsYUeXVcevcu8Cc+s7FJ+yGFUbeYnF+Rrlew9MLSvhs2TG5oM28NDRcYHX
EwMOfdwamyJOIkF5GInqsQV5O/YyKnssjCFP9PfrGBxsMvJCzotvC45VBeVq/vtCso6d/OhBVK/V
V+S2MbRPXefQzlwyuZFMHmvHOffSJsRwEjU3TjviLvUSxfGw+FjsQunSXyJu1Sj4jbqd+e4Uq0YY
grY8nXCKrwVHt1CQKD/aEjvkumdWlyN2MPLN6r6k13aLdtqiH3IJLCVSNi4peNe3zOq5l94/20ev
djdTtrWZbQP9cOAqREszIDKX0Jd2A/ZzBOr/ZKVmhwc11bo8o9YrOy5KEkfJ2HYnKML2q2ZqWi9C
tiRcvPw31JLyN/TJhWrfAYn8Cp3/kTPxWSAVdzqmaLsPmj1wJZpvopnqHws2GAFpLtib5Hfu7ETq
P+OIbsI7FyBdA/Z9yFYS6g32nr4BmC6dRy2Y1eh/omT+6wIV5q++xbEpV/qFucxmRyhGFLfKYMcz
dOEIGLofTGjrWl6bP3jem3rlUV//QFVHOaLr+ttxwefZqxpizfCkeIFyC4f+mp+ZznpsHS4FRIC7
Jo0Uvex2Iw+3SdQ2AXk5RVcX+JYXbqNGXSWacg3GjOO/TQTublUlcpfd9eDKbnzuunF89fJU43KC
R95Ds7Kbt/8b1LCuKtjGRE4Y1K5kr1gEg/btzxT39x+UV4TFjuRgSNp12ICYTEBJECAStJuyEVcq
6/Xzpq3jzf5m86/8JDewmMEl5NrZz+aaAosvMT9vuKFaLJnfa+9jma3/lbdYyqw0x8GfOH/HPMFY
zBSAUzfyu5I/znz/V1SzoNYHYvPT7tria8vQbMyyDZEmQ213PpEpNMShsTIDm+j8is3S+Rlrg+BE
4kaJbX1jdVmC5WiZ0KbhR9l2UNBXYTNeB5GCyTxOTrvDbdANL0JtOl99j6a03uN9UgTkYwSKnpzP
DrtvUHm7OtN5LMT6p+cfZCeR5C0bXh6A9AVtk4j4DgTv8lv4uOCrQ3v8qaAnJlpofEQ9v6HzxmYw
KES0dx1uKciH0utlyX6KNdSvksKAZHtf9Zvkc25sqyidgRluCeRaTzTqvrO68d/Y6h9EPZB8Taot
/0j2jvtT2K75c6Qo3h8+Esz2fYAmHeUBAjRSoWa8OVZSwJWBMEzV34+nkj+GO83gTqdEIB5J6TvE
DFfFgbQ8aoP5+T4436v1NEi2JGG9DwUmZCPCW2pTBr8shNQSh/nXxvWYbtpWwS+Ahs9064FyITn1
xKYK6zPfKBvcXMg8mCsLD16y1yyQX+o808gFDj7H0t3U6mfs2+m8o6sr75RVi1BQV2nbmfTRo7Dm
fpu7Eboi8raaFks5mA3ZVQUvphUGSTeq2fvcKG+WysoUD2CeBHF6XohDT5rKXqcm8O5ysxT2hcrO
IGeBkhdosTh/H5zrG8Aee2KWSR1xe+NdFIJSlhZBXgn0BhtQ93SutsVo0ZYd5JVWXw7k9FdyQUHi
wouKao4B6HSMgRZh7RdGniZuT0sFbavt38Ee7EFuhjaXgF07cEh1WC3ZitZC2ClXp6T3SV9hdktG
gH6qGaMIiA/2KqS5L/Z24fFnxilmzz5elUUUdb9UJilw1ovaBtKZVN0KxZSR4MsqIrz5kMRR6u/Z
OxhwQlKIk8TsIHq4sojr9jmn76MTwDx2pCNKsew5NuyhfR4bV91dZDRGpaBNnkhfcPbxZF937P3P
z0GKE5VM68ysFCo/difjW029qFATqzRKsmRcyPI0b3iuBzxghFbNBdHRciBH1pQWtvZHt+j8JTI8
sWwZC0B+Wv5U0rbU9cj03pHZPZUDBbs8aejh20bm5Wo8IJ6gCzmXzj7dYAHYoAvHkWFY+w30Jbb8
w3HnflslRSDByMNPyOUewPXd1AsFLXktY5Agm3Fo73QKsHVIAQEdxq82Zwy2/JgJ2ovrunQNxI3L
7sOxke8eq/oxT3mgKg1npwDmw4D2CeSMNIVWxLb+ftGGDA8Gpn6G5SggV8yX3EYPPFFT4ShmCme2
CC0IYFe1TcFYiX9ccysKobucF4LxQGmBUwJ5/Gub7dATmzHpIBvwchpF6MVD9AX91Eh+b8H6dplB
4Sb9uAuzEx2BH7rfn9rpNOSVXGmcTmPQ+i4IRxcwCzP8ghiQuV9qU2BAt1mD8TVSYWjVukfwiIRV
c8tYI8TfuqaIlK9TqydQ7juKhHlb4XeUu4KxYQmzfCJqgPAf5hgcHt6cJAi/LT45ucUUat2LZeKa
knMK6YMEhC3f68hHatXyISr/9jOCLEfEodey/pYOZT0w04Ld+mVy68MD7uyzbKbUClG4e1Qayw45
7vtLXNM0o0TLWBndW8k+ibNrz6/RQef1AL2N0hWPz0q8yZ5tejVweFENxKXob2ymrHrlCsmNw24F
iRUFdv1Kb0M82F3sGEMdv69RGGm0v9Y1plJXhDykBOWHM9CCc9qLNHftiViv8JyqB8IX9YRADH29
DrDgPQPpBWo082hwdzDXw6M7lIreM8DjwGVmtMfOpXtZTCd0aTnSEKx8BpHjk/ccLFLlcBhX34dF
J7UTVk5CGO2ZMS779KKB/plzOKPFCFtgQAoIB8nO2h7IXRdRuH1JoGvw/C53ysEMezKHa+ycN2uJ
NF1duCLbZUawBZGdPjvU0UK51NKLwMn45b+eKBFLNQPZi4tj0jJr+k0+Lv5/u6Dl0d3qfn2UFE5G
F3fA/Mp4bAIx7b/vo5A6/CbXBnpGTJ0E+8i/sXlMYxCbK3r8j20mQRXveCLO9CUpue45gAtE+kK9
KceZkhvR+NJLC2UUYqnsxcHv1HP6enE7tE3s+6i9MF1o2Y+hp/QItAXMJ0EFWont5787h3vDNZW6
met8sw6mbeFa9BvH+x00WpAha3kzFEEwZMYWbhmz7qsgAyuSoHr+wUublRQ5UxNUPh29vMe4L8EK
gqHfeyer8sDUajVgZ3Dzezulgor7bQAVnsqigO+OnQWnyQZTxXBGThPTKljIC8Fuhb8fkvJOdtyq
oQW/4sVU/J6lq/GKj6aNE7JFquXUhwUOEbBr6yf0EELBJ5nAdEh1BpF2r3jTTFpox2KVhJcTqCpW
FD+p9l8S9JCbeLk42u1+P0EvXt6+JIzYkB04TvcFd1yrkaHGsAGlEQxHGST/MOjp1wrFar89TonI
AucO1qKHCh4tLQao2U4mAQGwjUeHYlRmhRUwvCrr5yBZfxW3h4DvMGWHYAUqcRM/gHVIZTjh3OqR
eyeDc5ZllLjD4t4hW9j7MxvazjpA5bA/ViDQVR+9C4TUY9I+m6x9KT1tlPS7540SgfH1Xovt0tjY
/xMVj8CLNrvAZNUKssk9hhvZJJbm79lWEW5tw4YGCSHM2IWh13/tu7I7xogr2NsAD31TUf05xqVx
HWZ28V4u2ubM6fI7UlFh8wuZmFq9lN4tU9sXOCLS5vPSSwXJFQKHuL38XcyjB6Dk5Rlj30kh+Ank
WfRyu7tsqsHm5o/1DnfJWqL9XMX4N77otP6v7bHpeaM0AYbcdIthrBLvS1XxM/1LL2Hb6aEvkfHU
hUi20CAwT9rWuF10fICg9MSFHOzaTCLWl0oEixsk40fxn0XB7yDPzog1tLefvF5x0BKA6HMj1apj
lD8D5xZOiWhL7zQ/R60PIKfk5PkrTjS+2E4ZSITnf3Rao8e7WYiJfylj+fMINFlhrDDvzda/Uywx
uAKl06URFf9zpzMwr+pp5hDRoSeep1W7NW2NHIGyawId9lr++Nn+QIu0bBcRxsO1me5ZEsLQ6SnV
xf5YjauDgSwG8lfaXksdADchKoWR/rlOXkTc0Fl2cdm228SqDi/DziPh/jdcRk6QHo6wMlBCiaZC
cSPungKfNomYqfDs3vl3C9cKqAZ294md/h30la+8ZTTJm2H3wPgOZZomEPvtOLevH7Dukbkaz4nw
NxXbnRciKF8E3WVu3rp825Q2fdbSl++Zt5A0c+hFgXQ0Y54LZ6TM2MrLmKh1OaSDeG/gpurjTwrs
hV04t7DeMeOod7ySIZRXBgJf7tns2Z/VsQm6sPuekmKntkcsjAIipdcT+C3bcQrbi5YGqabOpNvM
NLJFN3CnGsbfb7LlvZL5IJZJnRcV4lMcJBvl57LuWOgcoNwnfwYN9ujvwQR/wCxDOekykbHyXuhl
h/a74E6Vu1pI98WZ/X/TxTNjtrYZ5z2tgDsoQeulT3bx1U3xoPIuzwiJMbGtod+aQPhWXDGedR7N
nKiUnOd/q+YiinyQgnGCvOW55Fuyiwdqd3D2WmYDStzu0IIG+X9dsxEudtgFeepsVZfNDIRTiHc9
MYaXS6O+ly10aOe+LE/QiJGTWAxY5yCgEO1ZAxTtZYEAoDLuZTwNOf4EnZqU4FVio6bftTmdv37q
OMLHA6h82gauYtRqqYI9srLoZiF6KLiF35fkPjLjLoguw/ww0Cu8FsZGT/a8lzfS7fSgDzfIdVyh
jnh1r5gTgptzN+Ukopqe47CYs4+hikIRrHdLnIKyoULpH3PRjO/+pm0zcGNw8+4GS6ELSdaoe/IX
7Baxi5J/WvafbWx/K2beIqG5rhmxMts3ZqiCoc11tasraMbbKkTL8/+bGT2m5e5NuDJ/vcz8XxiX
4i5T4QpZAsDQLSe13H8kEzzlCuiTPI/nOeaO6qT/P1bt2avvYtnqR31TuNkGU5HKwZ03NyZKlDrX
dHvcbedddOjTPxEf7f1rNaMXK8KuwahV5iOrDO3RHSnJAcF1NAJIE9sMYFlyaw0pATLZrwDei26q
ZqMT6kDTnvGFitO1/R9XGHhfNnRZXPG8Yzm3/VXNNudQx7JpER6ZXLOjq0w5TNw9spXyzbcr8zcw
3nC/EqL+Y+Eow1sBmyAS25ljNHeLCacD+piKbtHpT4ZLPSF3LrwunyPx5B61Zt4FEjxvH1+j2Oup
SGS4fkLg7Pmp7pQfEYrTejMySbNUqLmnk8mdlZ5AuTOJJNCdzq4kfeAnaDT+D9639FPKOEXkQSye
q2Jwq9D4bv7YvlRqvd2mA/bS8hxpoLuuu0S3t77VObGDb5TQG5MXPG7zE7d3+CpX41mawdmYTNO7
tXl22Fdw0HLPtPpMO4xc65jJQN80zjcRr6llhkEbsbn4UTXhGFgJvrp2Gd/ZuBqPO9mA3KWXRQGI
UcPAVeWCOadr4xdnztjbDzmQ1g7UBZp3glH6Y9peUsKOCmcx4aCRL+qJ3E7hnIjKy9ROkrVHaMRb
PZQHnJf8lBtgDsAJcbD2cxAYKl+Lj8AZwSXBXS2UrbH4q/cggKlG1xAFl1fssQ2ulxvyDYAP8ZJr
JSw0KvXzAUTd3jQElprE9pi7e8fdQE/+EGQanfoKyyf45TwLUbjHe0GeB+M7zrsIPy+0GgKt07qP
7EZPZFaqyUbdB+WfVsauBTc+6MBbBwcFooUiCz8QjI4bQjb1qhoShvEAYSHGBSWZdT/mR2KICKqi
25sSEvYA+yf0UKiSTdc6Ov9Qk3EJPO7dLyKar/rSCDqduT0s1mPJ/KGWICNtS0kfDgqut+UljfOT
cti/+/SjNagdTsf0bF8AzZjHNzi19NNwiFz6V0ytnHbtpX0/yMbe8tXEq2OvJwVdrS6ap5XTBZFA
zcBJmkregBfBrMYzNPwOmcaMpZbLIBiD6PI/MTO7vfXjKxeQIDdV+kKdzIrtLGTbTu2qfQNIjbEW
FUGDAMa+QzVBwFnxjUioytIJG2HPkAI5aOBmziEcJMWGTAqkwBs4RoXTvTnGs1/56x1mwGtyGjmP
wra2hRsXyGX2mE5qLCL6BOubs8++1xkMTq5fGNDyXVsBCa5Wob9BwOCaFKsG3rk8Hvpktr+FIiLR
7won6sDHCg8coc5HNMuXofSpGACTGpEYPStO0qN1cIpINC2ffY6bt904jCiL2Xo0ySrUyy+4bHPP
jar6WzRfX/M41c691ttgjDZtdrFnaN5j4ufiOoN0cipgr3UDgsWueUPM+YBP4qqdFLzqyl5qC4oW
vnn2vD9EE38SnGwR10YWqYzvuXikuOauPBoxySuFyba2bkvyn669q9dD7hQlA570c/0FObPypHxn
H2NuOogr2A5HDAyb6PokC7oLZcRvBGOUTIz8fne5/3SpV+GL1Zch2X6AGru1sOWMtMhcvVn6aMqV
kV9DQpr1fBXgOYxzGLRqgbag1/W5gZZlXpLHwYgL0FyRbEU1S5RxKl79lBg27DPxGRE4qtQjOr3D
bAHxdUTYYE0ZkHTTYotMMzTSOUwa1ockegrmagqV3ypG5joCCCZx5+PKuoJByTeWZ0p28lcnNdPm
OS5ymYRaCYSmT2lUUyQy6BD/vOMw6ivDLCZMXoFHyuRoG4cd2UK+Yo9Rnf4K0zJSbIQ2i/mS8Tn1
QqUZBVdBwbXaB9kHG22UfRkYdM8+h2VZT69cOD+68+CxWPFl/uTHG8VwV2voK9OEHStLfeZ9WTV0
CFBg2QBF+GYBiSUZxXcHjFwnFKwjXNULPEOhI1I/fV12bDu3LC/Jg6FIro4urZY/oY3PZxiqeZBw
0/gGk3XHxRFLq7TfD3TOxxyIgziKXl3uIyItdBAO757Jz1GxYucHU2YizsGaPdLssaMr2EqtnHWG
LiBekkvtDH2n+tBAL2ofqQcP23TC9M1bpz+Kb9yx/1S8tPg9+CAhxXb9SsmkWdCVI54mWupyL4wy
YMJHTR4zBSDEmvpaEbKLoCAf8NKZH1Wj3Zjh+RS2qqPKu1sh9B+YfhYhQaAVeLDqrLEr0lCT5qp0
QsGqVQRqeHLp+7mIZyVMPxQGY9hwkUqlFrysEFRVD0EEG40Bv/MQysGx6C7UBHR9GYat5hG+of1W
QdA5kDon8Kgc2j/M+H2yBZD1Pl2OwCQOojf7pMTNAItwwN/CCKQsEJj7AiCJRTS9f+i/YysxgC2+
p5s+H5ZPnuCf35oKxu5a7NGG421h+Ie9dzG+Nw2OQOi6dSWaLtXFoNhlsP34Fnbz6XnCymFojd6s
C+ONVxdTsPOlf/AU1AxOvBILX2wnAbX4dQ1iSsYdUSgIbBgk7CPqrSNiI/T8KNohrTOVApbllfbv
wksgTqN/9GrCTRjglgh1yDm2R+zwD9Yb8PdBWOJHdSX4P1L9xBk4ZDwWbfMpiwqS2j4ABJVrZ3sz
L6GyhnH6aNuMS/H8FPUERbXLvn8NwWsFGMAAKbKYel6/wzdqoDLa67V59sNULBg1X9JTz/AyvJSZ
L7fcKalq3zR7HkgXVesPGI1xNQYh+OQf8jYAhPIP8NwOrCxGbQLAcUiVEDCcOHTuEfXsMJulsAqp
GrZ0XswcFkGMPHECsSSt4xy6rAKTi3RgcA1d3M3GADZJT1wMcSGTHa2cpair5iZkqMBmEL2lc/2+
p8lohjoT32PkhGIaGiM4d0xqsLeXCBLNytzUMxi8oHWK2W+2FI1S/EJ66FgVJkNjKJYytA4NG8RE
l0j12UuE2Xdz8w88qT2Oc8mIn5aaZjd8f5J48C5QEv56ojKhM9IOdb/IalRC41Xyj5uqZcPHgTwS
mxowEe54jQ4hdbbzSrZT3QeEWnhTuY+RVRdOgHluRccb2t3L5U6orzsddKpyl6zyylxnL5+QBIi/
7qzB9XNGHiTdDYZ0ousfFIv2C9zuMg//g6RIaUIwURKrZ/cIvW1H+qt2Hbl5OCLKRygDDmbCiIe4
x3Jw6jwvEvcfkGOypiyWfeZiE4JaZqlvCmuG+x55BpU39vwgEYioS8jdYSRoPWRmf/L28p/RWqbQ
kOo4oDXwLidwcrh5lwewc2gPUsxMMVVcOzsmXxXKT9ByP+0OHDDcJgIKrQhpYSfw+006VKhUZzmM
d80C5SOH5HJ0k+t6/zHmxFNIYQNcp/65BA9x8cVXhyiTeE9sMDUjtVZgnErWbCqeZvIkTL84/fDo
QlbCasxGT5NX5n4LrKd8C/Md0LZRuKQcK3CFm1t7pDhIsKBidjVlXvd3tMPk+rktfWmWm1mp/uk4
4IYJnzsDyCmhz+dq4t0RyHg8CIT268gGYLjZXQif+KEqocqQAUGzJC2jmV+Q91PaaBXr+R9kYjhN
MfgZKclal+NTfzfZ+VtiQ0Ha+MoO+HInw57b5esJq/oKbj0oR47WRnaaYaKDnRfKJ77U4QZl6jnI
yY8SAzC3iOcrz8Gw0gulEuFoIvn/DZYEE6hUykygRNRuZQCJcxdp/MmN5YxnNqnMwS+NHOmE0sXu
8fbXcVfH31Z0FiO1SKo2dQJm+7xkO4/JgGYPQrzER8A43/+0yKVsquuoZdOeLToLWeE2aPmer8Fl
caS4y/NWlRC9y13FKikiUgXHAt4gpwnJuoVQDEpVlIT9mHSf+3esLrrproPb6BPC0zmfttDD/Wmy
4qaioe1ZdIay78qyswssy7cPxA5581enPqC3nP8hpzA5+RM3TgyOPjhbisf50tDjygQU0pJohNZL
4sDCSjVpm8NnnSQx3CtVcqVzI4VCFhl0jQrL7S9bpN5lyL4Lfii8BvOzlczRCFhc3v8nnuM3CdR+
rHR3lCHJqUhAo4c2H1UdCUeN1wcjGlppjTNqju9nPSm9DdSizR/zUwrzpp5+EROLrJ0Vts1BAQIM
X2w4T4Ak9VRUrmfdbtupuJ7cjnRNnAC1Rfw/xyb6sGYkHYKrg9cEHJM/DVlnCTLEYfQV53MGjlqR
sQzCZDFzhmovQSulO6k9DvyMpA0BIjHqvf7rROBJdGnrEXhtblkkZrITdMw/RWkkI4G16FBkSMAM
9RCmrOSL4W5o1b3xv1CzxSced+6HsIRLN+DlJbb3oXjyJoZHJGg406lbMs3E+1efGEue1x+2xIDu
Iv+Es1r06mzs8wNfNVTSBZ5K6SQgqYqofw/W1nKdH/Ge/QggeupHsoYAGtvuzW1BDcqJipitOEVh
71X914zTe/iU3wRAAiMdt/4bmbwC6COwAabkOiM3TLM/E22ZtgsIOWSX7OF1lCxjEc7akrYELWeR
IUOS4Zl47mWCIWSksIi0f5PPOTPzWpgo6CLdLxjiSzQud7yfomDpjEQCyDXcjcORBMQt7Cn7pRsM
uDQ1eouVclv3oysb45cpeNdPA8j2LeOSeTDe6fJcuXiamI16u/trGdqeRwqH8QHBtgpCAjA4ozCI
h7AGz52UxNqEl7a+402AvIJnW51a8rbhhCgKld9v6PoOu/jKcN/Xmru3g2snFsdCF+RBH463e9b5
TjzZCCIiCmpNj1Qz/Szcj0aA0H1uLW1VhyXNOxfaGXFdWNZPoem2K/0kvg+KWoFdMtDRsB+PmqOK
k0dXdVaQw69+mx31D6sp92LA3R0G+96zsjF8YwkzWX60nKWXlf5whhmZRLkh78CUKGw/bYr2Vnsq
Gq+vYXPHUZU7ToQ569aSdTMdXuxIr5czJXQczsyvz/ctrtyLsHbhlhph3xgKNl81y8OiMnWaHl7H
bJ5zmzWtBSvYHQEk5FQMs6i4qUWvN/1Dh3EAoVQROl7JFntov5/cyO3dxQfUSX2Gm7Uc2VOotYxh
MsTEc+AcTosWU/ap2N6RZSWIet4T3G2A0X1eaZQ1Pi9z/VYSq6KZO4YAIV2pSYwMMjO4MBVVG68n
yUHo05KoDscrmegWmzRFQqR7ZdCxcfjk+9WKNJxN7ZumQnEbRAHENFG6WaWxK2CaccrnSrE9ljfy
KchQXQTD1H3qXX5qDVNDM1MBx4k/BzO5Tp6XQVCMCdRSIfjO94TBIqaxotr3PeIrevRcJ8UkMcYn
ofPRbPjmeklDv6RuKf5O0z16k+lKz6MpBBDlBtvlu6nugu5fcTnr6DXOA8nckSbKWqnGljzhOTDE
THoZGF02T749XW1aujctRnNs/i1nqKLUZvsVd/JgMN0F+7hRgUzO6ktBe2iOzWKOpY7LcmBvR966
9X5SHw+V7QyTRpKGqgSKDsAPZfjGxKfNWE0ExbMJ0w+/zit5YdRXl17vCAEhmQJPPN5i6smZJVp8
r0AKD0v/ZPGgsbecbMF/Q7PAB+i3L/leb+Fe1nlHUgZFk0kfOCStLX601ehiihqN9VVVHpC3fsKK
RM+N3qCrkWbpUUgPv3Ea80sKJjpkMQNA/ZNd/EqA8hWCMEQfbuo6XmPU7h4nK13+TshkAegLuxP8
ud2wemr5vM1hpIam2Tr14edj9Gf2y/7wOMuiyqwEcBVkCoz3dpZNSdFpq32mbK9ZEoweDb93JLAC
XvdqSK9hEDZkoH2BNLIH3icvVEb4QIpw1jFG0BPVLOdmJoG1pRiMqj+sMqTkoNUMvMsTZ1RBTLNJ
7np/aKi7xd3u00qOjq0/ul9PfUXSlYHztwhVxW0rMqW3pTqNrV/RZjmjOR3BEoqt9LFd2jnQkr4E
oFAlU2+g8+MmhLErrejidZZnzpgaxlz/UX1PhZ4q1ccFeTCr2ZPT8gP35bjKOiVLJyjYqM2YnO3h
YOToteksTbsHsYTEMjYL6KEBYdff9Jc0j3V4AI8QDj8OdWCzgIy5Tk3smz+UTJOtiGLQnb5pHyLH
vEp3Yr+XzU9BiXhdfUFOoAQJ/hrpLwMJWjp11IUsqfODQmcz2Zegaa65swSthr0Vh3vWCQQ7K4IW
pSTzob/P0pCD2oAOI3X2NAfxYV3Pz20KGg7lv0pM5ORVBe5LGyG5nZzFgsQ0ZZONWNbpqi7F92Ko
b7KwFRs305tJSirmSiaPVMLRZV6eBFENuPkVdsHojuK0uV8AjclsEzeBJjurlIR9XSjvl28+76xQ
EERuDQHWPah7E+o++giKAF8/1Gj4uPvGfPb8mfXnil2s/P2wzjJTmJR5yqbQtviFHYSbm59etIY8
F0WlPSevATpNGCZi7HofX7q/V0p4sVCqMg22Az7CUxlOLLZMprwO5Bu1nsUHGJ6GB93EG/MObWYQ
Y4O6TqVZUYp6uK01oS1dk3zBtnTOQuhH7ltrTfpPirGeObBf7Srsy7IiUr9w0I210f8URzsLSb8s
x+/UWmTtPyzosj9G8+SSGLgXUCEIcmoyVoXD5ZK3aSkw6rG3Td62iH7KOItdQf+9vdupE73VF83I
DrFEnBqbi6fdeq3YSJkHf/OPugVrW0ZQhindO5wMBRI9CcKdi4dJCsNzakeZQfiVoml+gU3B0E/n
zoect0MWVeSPP6MRm5moTgaX7fSIiIx16upp8XtdJteQ3xo9Lv20eIOZ1Ojr4aV4516IUzQu7tP+
aXdwIvO18NsEk6sqYVhZu5SY8nzA2jdckcsgMNTeCfmPfFHH7DhGbKZL2IzI4aOpT4b/WGIa64oI
ZTt5+jxaakkHjCB31dcr7MhZPf4/FgsoqbrKfMHl2T3Q8S++VNjIPXS0qkjY1X+1NfmWlOchbCxg
bwHHzwGPLAkN319hcaJ+2pdmX4GeFuCaHZl1byGj0BSdn/8LaN4RIIC8IJdKrRgcoVcpzlCYrIF/
nQIuSnuvxPina2ilZFplDYxiWNuB0/aJyTugE9nNsua6YBpNrb/7FT7gpIxc/YArluVwSWLlnFlE
d4nnKhg+AADgygb2WX7J6bbqje5VKUWLcCn1cVczrjGYFMhp6eByOqTDg3Je2tqleFRUI9r9s5Tz
xOPUonDKuSrA3QY8RHHQA73F6OOYsvF5T10Z5ErucOWxjboNcmRQBK13C1cpknvw4EAddqMNITbP
Ja6mpsh3wBEGYF+SSXMVxNv1ol4hiN1ZOHCE+zMekLYBlOOEFywqbjbICmVyE7KkVB0ojijiO8Ip
1hfePrYuACUdajcxUCuJbXy6MHXQjKCOQFXK+FG+w3mqWjyL8fito5p4BxE5AYyA1gM6LFCqqWZV
yv/rcT/yn97j/nxyMB3+b1YA4hcZ9gPfvfZ/67dNND1FGfddldp7WMweqMHPzA+8s+YiTYanrKWg
rhdN9lwuyd0S98XgxUxT+LXghd77bq6rXV9ruRgnNV5HnaLubMWEXkqu6roTZ9R5NXSMv4IabY43
Ab1ERiXOlpMGOiQU7B53MQGq49Easd5G63S1WGZoaEevQYiqlyn+Qk32mZrAWS80XTU/+UaTJaKR
wm9rdlxbOfmSty8WzaB1YkpNq6lclosCxYD+BggtEjZ+RLn3E/U+iMpqXgxLQ1sM5YR1+LNc1pgU
RvFsD3HM9r94Gd3Y5/OrjsJX44mmwkGSxP9O4OlLXFRC5o6Lqm5/mwt1aV5mw9EwS61VEieBEj5z
zUIgq0doC+qe7yo+VPLUBoNChUkjA0k9vTOvUMxp9IyXXiQNRHMLlqUPcYHE+3oIVN3IU1ukufQU
HBMCD1FB+Gjtlnc2S7YetG0pjA0ZIqhK8mJJ78QUgQw0NbqXPBpmRT3O4ukH8sAXslHs0YIKO8S4
XOjbITtW0nx5yz/cignW5REBLK8g5pyc8qSWsqcEWHcgqVKUkkRybQUW5tVVXSS0mtDiGvYJjtRl
vp8SbYY4Q9EGPXxu/y5T40EZ92UKTdZqGRfMZpwrw3OXnly+DrZW22hVLhJW8bM7jkmH27GThHfi
Ea7Y2jTuBVNSSr1f9BMMxpjxe5E5nK4xHJqURCZc1NwWRXHL6HiZ4drqSKoeGkbj8YQ8X7RFQZbT
tuHMyI1XM0zgtwYWBQ99/4gSPIfWPat43kr6EACpLjnSrDUrfywTSDU5GoXE8kth/fd+/YUkabdl
iXrgub8508SHz0shY7g7C1lU/Jegkit9MvBmvMSieTh+c/pRw/6Q73+8DVn2W3/fDPZf9JWLsPfV
waJKZ1Z1h2g7S2rtIYBgib4gAm/0XJIuDdIJ16MriadlymKOR+btpu9wYhmu8fgHPTjGZqFHjRFl
Z/F4s4jv3XJ8X8WWD95FR02YAwZrHY0ZOSBw+DBiMAOn73oEa0lQK4cQ/suRrW/tJwDmkrKB7FBl
CKbI3cHap4rXCDnGkh9J0e+nYfwuSXVjzWreGl8EydoTvW1loF41297Wx2cNebk3FWYNHi7VZSM3
TLTVSOvmIciBQfboLdyaga+NWdXkO5wlevi4aplaFv64Eie1ZQJbUGh/uMUYqvHM5E1aD0J0xYPx
0gQgpnxJ3f6tfhDAdR28Hntikk8Jb3+pPuv2vCkUhdh4FlMIRmoC4sZbaVcyY6/pdF7ousFHDrqj
K3zTyW+/QxspjGeCczLqwB5ArN8wHipY8o34/OR7MdgEnTmGSIf476/Z+fHHZf4TmEgQiQocuBOB
LOilJuaBa/r/UMUymbuyFj8vD0mMs7tv5PpTWL/tK5x1La1sxfc8Q1uUChC+yMf3vHQpK5kOA5NX
/q7f1I4meHHmDPKyTaAE2VCI6osM/1SUs0NgaOIN8nc+eYt4UDuoGV3+KoGsal5jUFz4GrrLFCie
VSdvQiwk8NKRjYZ/JZlijVlAV4QGwyYaBfeK1WQ3qaSMzJXKubsFxx+KGctdvFfZrF9dNL6MMsqJ
6KNjugBhdF1eAN8F2bfXQGpHZml2TCqT0TmnykLSHowo7IpvoOthqjVM0q8rafjpvMPuFLH89KIC
0wbtCr6wMBi+WbXsRLDoHyXaT+GVVmLeJJtIzG/trgfOaUAbrtPtuWG0ohPXMt1rkK9QCBABtmvH
3saRcz0zKFb79u8/MHBvQeWcPcMETmJqHEKrpZdYfZHs3cJTBQabRMZKrYrbS/s7Tzqd7MGhvhXD
7Sx+CN3dO2sSKnKtYA9cMHg60NM0Q9C/kDwwWx6R+2rZUJyEoTwMYt/zKl3Fey3wJdQpyIW+lAh+
KT/2jc6JZv002Mne9JP5RP2bCFCLHRTtXAf+7Ozv5uWtf92Y8iNuvGn36DlIw3zp6OBs97lrJwxb
fmZEWGzGGwk0xDsK0nWF3NZhdYv9liC1KiwfsDAYwnVyiilbydE5qrwpPGS/ad5s9R6Q2q3A7wMA
zKe79Chft9FXKEBFtwCYj7IsOs4R0W/kSCM1brSPDKR0YHL9CfAw6gsALWIVyab6WfM+FjYlGYt8
E9rWuiyCdtJJEONutTsrOYpc+CVo5j3YOOaAN+tR7DHhzRdtp+HQk4md+dONcRMOmHeM88Zxd3TE
M2Ly1Rpwk5RPkjIjmrWKRuSTviurWwOP0r07y7LCrMtFluHDOnWCNQCNJifnqTLxNvLN7hkmbn1h
Ychkh1lWztGPL8xZIkdItGqwCm4mt6JaEyjsI3l0N/XltgliU7r7crwDscXfLxK7e4wbE6EgLkEU
t7uTllhQYnvkS13kxcABwuZY71khTh8McdFk7D+w4NLp171ZcDuy5vRffxVSgmlMwZeXam5SGmvC
/t09n/SvXAQ4sQImK5030Mr2YZWAlqmm8Sx40o6TYVxejK7UkRk4CKI3DZjWy5+tpVR3n76H0xgK
NZiCCuE3CWGTJmvKkjUQjIzd5UMost432HnlfbD7bLmFuhS2KjVV3sQgG1aw7P/Rj72s7MG07gms
oH3k87D0HCKkHwR1vCkaSXfcHVsMzrbyEc18xbXpLKvHEzpioAw9k4zx54qfMbwpJmd6bJ0iGjT4
bUIZWY79LUZH3gvujKUjasxKPqXdPm192fuEolwZE8DSWGXfDSgJKArzZ6NlEjYEz2EYcQ15qj1z
Zce/ZDzybNXPwLe91T2BVsSKJyfduiSkfh/N87iQUU6mnBjuK93DJvIzY6RoKsMGmcZqWVJ/6ndJ
Icb+uFT8fKlK9voEKnaBkZW1lZCCLmlnvcdrCiOfJ5s0++11DpKc5si5mkQ97yefSVcSHUliSFjv
z7RdVCsZKgCpprMtHM3nk1gYYrLBud8MS4Nvkmp2qkrYfgmPS4CbMg4OYYynWHiY9NdinRJpgpns
kNSTBO79HpJNOwxlRUZHFh60G1l60KZDq3Ui0ZO5qFVprG+CMCfxMh/d0m3aTHHVTXXm3H80Rj9h
h3RbKMyUvm8zfbCj3SAXhAQWrPUD13d/M5kZu5gq7XrAzmlPGbUsCdge8vXUvDKu9QohrcVx/oh5
1CrT+NGOwjCBD5ny9XQOtPm3E89h3HA9QbdRTG5P+HptOorqQbwaRknAqmh2AkbnbWo04iNMjPUu
40WHpGczXgO0et0Oc+fnwanifwAs/DeSvGNHXCDCy9vCkuQ84F+9P1p2yeDBXE3K9leBvNJjieiF
h99caaRbTgJ4lIWzg4ZcsK3NoVRRE8i0crCDQOKON4jgG+wrrYVpisebuofdWwCVBbK0/s8I/2ov
tGwvQe8ge1qjwfHae6gisSl5pNMhDfFgLxfNL5m2HOdZkDa1X6QM6Nrd0QRXsnNl61zjgQ9KBiXY
6XWrCszbEDgkRDKnaFnQCxY4h520NpvpolNcchdBvvBikjBSVsIbwXOcKF8oyQvWtSI4ZC+bcIIz
9rJ9Pm1LbZASTPK20wFM6x5HqqSUvjvra+5BpPZOPw5/XE+4wdofI6VHBZTJwUJS0PHx6nDmMLR+
K5LnKlZc5YmOEDGlbYWM/dWc0mVevgtUE+M85n7om+W2sH22pOz5PKMyTxCfIVIUml6rkCIfhvbF
xftHwq0D8UiDZ8sTJR1W/zIGbzgJHN9xohpCq1oMCITiPw1fuWKvoIC+f6/EJvN5m368DHtKtw6j
MgNSEewfay0pd7hoM5ZVmWkXHB7RPZ6ov2fge7ubTv8Y2SLjyEXVEuIlQSZfg3NMJniMVCnulSTe
ojiJedMkPZSHKqMTvzzxwRJrLuwEz3mBPYHcBnVTSgC2V9MY2CwIkMM6ZTJQb/nzmDC0meDDwGlw
Oydt/MRPo4Avf1OW+mxOAi/Yaz2UbMVyAgdHvfdEpcx05OauUBD0JQZUdrDGahuGhuwUeMP2Baq6
WtENen5rJOMmhZDl1ECkt0tfrRQ1zrgEdATsO8Uj4iU729h42M1RBBD4PwlFu41e8L2h6gBeTPQu
aPL5O7TYqfKn8ty0a1xkxotGWFlx+the4kuAh5SOfisrzF9QZ4ss2l34CCrN7HIoc/xMFD4wBLtv
AvfxsqnOktIt+CE7hZs2CvyjaUAhu3LRgu0obg7EwayIx8mRlb6IDOAnt22llqxiARF+jtQiX9ti
sLrWKDFhwGk50l2ZcCiDMwxasUjBYwblVtdj7lwKlwX4LuQXp9li5mIIT96tjmno2oFKK5meRBTe
m0HLbuIfz+AiF27rdSay7YhXf9oxq4bWdkLXby6/f6Gk0r46+oSV02N5hj2yFUdc2RjyYyZTRg/o
84obNSO1deKaXylS/xlSDCtNFdjxuvXNACk04cuXOgHaQZCazNu8m8hIm0piFaAKRxctm/L/sZHj
xYpcsU3625Tu0uQaujEn9h8i/qBkN2B3bHb6OsdQQHn/6fdEG/J5g1XuGLei3B/4BdefF5e+gbhd
N3byjxL+ZJkqJt/TKgk3blxgT3UhU14MThzRTorqNDuGwA1qLJhQTLqPiCG4oJM/JLKz/zLdTaUA
wdl3czLpI79DEQFFDkLlGuPE5rYHpu9quepq56VPAK1pMRUQGNrAPftp91J9mgGj5gV03nlIeQt5
K/WIndapgRpZAlaMjCYGeY84IpQPMaHq3yTvNCtFjkfNBxmjmjwNlxlME+LcdLxQEYFu8o/Fk6be
nLCcAN4JEAeOEE1ac5a30tGmliQM7tR45V2JsWOzHnwgRGSxX9DxPjJj+vWncpze38rwBh6SoAMk
Tg9m2ub6Ok2dDEqabweKylrMHyIruzEiOdMlBQcu4qIP2Osdw1mVZrzgMfilP8uGsr/EuE8BUxTS
qD783vfi1SvTjHfzptu6W3lxC31ejOCQTTGPbCgVTrOczQy7tXgKKkzr4fmncyq7bD1HtAfIgm6u
w2iOaqP3wcZ+WVxxjoXYvClljNycC2ZKy9RpPSdpebsnkix8PvJeFHswm4BQYwMp8F6PZ7I/8Q7A
G38FDXKygXOUwjdPMVZefpPjTTEC+nUO1gagZ3VY7yXgJZzB3abdY586FSOO+PsPUzsBkQaqmxMo
eYyMl8d5+aiOYvBT6bgKqPvx/HRjAkQ7NHrcsBkDgW7F0NJRRixOaOv1BISujUDtAMZ6dkxE3H5U
r9sUHXPkcHfPQyE0v8U5jzTr6Q9xj283+KeNLzRM1ZS+9jCp6TBxKW3NxO84ZKBLt2w0b/5t6oIE
w8F750Pr13wzLj0SzhWnDfsZtHjuJSkTAvMBWYGzMl6YM5dfOg76dl5fp3gMmZ/GQlFNaRdYm8vm
lmrenkVdq9QURTJu9wHcGH0ikFBedGBRtD8T7KZDlk0sHyVt3HLVxhOCNQuoRq0TaLcg30+Qomg4
zLtrRnvVXd1I/RrCJIybScUIzu7pybazJzw0Y4d81yqKmAbcis3z5AWDRKbyXKViT2f8mXzcHM0C
9ccAu4ElFQHPjbey8imFlRVwoRy1yRMBqpCQkcxhglFcbPOVbGHLY47+W2G0xgPeZq6zYOeYf94q
FNbem2+2gK4smwvg0EjZhq9AYcISx4W16klM5M727lrf3QqXfDTe3QFkj+H9GML3unQk/4duFlI5
kIfnbzXrLdMEtfpPHDNlzdiQWViTCjZBlFgRGohbeI2LRXxi6xNgKmoSsMuAy/GC60vTjUfbrNIh
S16UGh0bT1SaWe8VXPEbP+3ovb5yFwkEzW7atEzV+omy/r4lMxzZzORagHpB22rrkFgH/KeUlp53
SbXTzZl63ZiRcqocX8aWnwd+S+7IoN/eYlrTZ2oaXxng1bSOZRzamPPGZhi+2qI6w3TIRPKB2jyT
w5iFhNlmKbNM70DnP7FGrk+araVAOzDLDTWoJF4SFyEjtVvTgSjrbG6EWEFPHmxmI2d8xoBZDLOW
M45IumX5rGyYXq+WfaBkI1v/8EaZX+Wk6fOVlcXpPJAg2BBzdFmGEtTDuQ8NOWkyET++SMeg7G/M
3gvSLdkxbIv1r0a8EXMvDdTSwySZoOwxY+T2GssqUr/XFVOpsq2Gc3GQkpnHxIl4Z1dneDtNPfqP
GaL+e/N1kEfQVPWhRo9/kjB1xRShZM5oMqsxcDjTKNAiUzdIARwUsWJqyQBCJUIY/OIr0bGoBvbR
ngM4Gkj5M4Ltd0jtWBqu/on3AzB1+rX7nymZ16dzt5ngZbip5sbobXTPf1zKJQQiMn52J8smplmp
Pkc0GYIThuApe+cvceSP9+Es3dwo84+0HCQJiZhomgv06Xt8Yb3biWRvRVio/mFkTiXUEVQ9GA/N
TJ6z7iM9nGsX+L+s5GpRrhOOSQ9oo5d3/oV4KQoZlheFEhjbhTENMHtIdYW8D4UXxDorHAenLg1+
/du8l+k780YVBkkwPCoRILkVghhZ02F0uPOGn4nmIPuDrbta97e4F2MT/OuZfoOFEwXKBF3c+soy
jVi+nyhLo2vWLnjAC2MFXQnPNiYdcQi6CpWq+JyMKiiXwX/4cEO/jjVaFBeanLfBWNY6B8PLlcmt
Dqmtx5anO9/vgg0GNurQs5PWAYBCtFEuCENyc21udt/8E0mlTXz+xAtdlWfy02IbKXVCJ0grssvm
joyoDzqLoyDzHjQLUINGrF1KAtQLXYdjjpXHmzSn5C+L0HsydB5GvqGP6MTPRG1y6Cm4LdssVWVD
pG1yeJSJ4/KgtHMiLpaCbcajc+nGp9rJtpdrP+ZzIhe8pJXTnjTfqtz5JMIZbuBzV1w88FloodD5
BnwucGl+9VAyXm9FmearPcfxbTQXIwM1UrdLngeYPbzANY4ILsK2cFMzjh3XfmnuxK7d4xGYLM5v
WpqHb+iZ4o0gahhw4FAKa8r3skscCgl/G57pOVcjeVwxlWzgNYcqTXzW2BfCy3YocnWVivI19lWM
57PezixHfbRm5W/LHZO80WJu8bQvbR46ilJXDvMuPkkYEPA+tm0jUPu4+xQ61CMsVuHwcG1PbsGr
y3wAvP3tU19XhbTLEleeKW2ndYvtYuW4OupXBmhwuz6tWsdmUAtOnTgZOujl81ToXA09XoBoZKHb
7WmrHec4KqtIEoSyi4t0L/h/2mRdWxRTi/wrLJ/wnLQZ7N2+GNvM5er2Sjfp23hAp/q/BrVu+jVO
1mGY/3axDXBTVNBpkxR/Zc/Il1LYR7T8K5Q6MqKQeO/fESY4Yc9hIBtbNgGNxVonfU6k6U9NcuOt
l7Er2YvLeTf2Xoo1kryh9e3AVSw9+tQvFLvvoCZ0MSY3RjFGYmxzgbf/S/tS3PQC0UTZKio03/sW
Mb9lwwIJw9JIq/HbpdIHZwnufOJSBKpMghivrmw8HVBhWzLS3Uz/lqnURbkHPTiwwLNrrbBH8lRQ
b53Vq4fAq2TajVO2mPQ5FryqXspelRplCw64tZh7xv8jcG3tDs4DV7YE+iDXeayLKqf2Ll8LlGUk
LdabypEN2a8hLnQs6F+Q0y4zHtsb+iu5rCnypf++9p2OwMxYCekj/vqVXirPNcUlHSocJpFgXJLY
eARyl27bNrkRJa1gkLat7YLnI4dda4i5okLw1O8Ywq1BPbJ9f4iREbC/P3yoWkCL0HXJh37xP/he
WNiBBGwTi/dg6LXR221pgrbaq7698PcpIJEb3hSzUar39iyHG1Kv3JNlPNGSdwfyVRzzkHKlnRnA
5kOyWh9e9j144wy4g2yh0OTF/iFxXKMFE2nQVWxf78dX7hnYbY7EA6gFfBbVoKY3OubhVpOlPujY
6bDVw+/QWe7UC2aDGTgsBfIf76UAdhdJ5aQz16oSlONfFATR0iU7mFAmP/Uovnl14I/L4ps5c23v
85XxOiwykXvSoQ/F8uRuw+TVBa4Va1ZX6LrHzlebqsnYgPcG1zEcPH9evhb0ogYoJEMXDfA0mTLf
Ly5YF+IYJqlZilhSDTTxlpU1axsU/3miwqPsUA4zgjy3O7r0QsPFn0S0iyThkuY+YdBK4G4tJ7V+
0dH1dT4ZFmI5u5yj5vwizU20JFGcWu6dtTveU7SWAWOvUyz4cKBPzOyuGK3F7iUMMWQaARYg7aEj
y0QQBp2s7EoUdFzu+BVbzAxQT5jwnYa/hG8K0UXtX7poVTs6kA5yr4kohBS0f9g3+1VZVdX7rkva
alsqXYG46viCWssLitcBoS+pUmq3gH3+6PWLItHyGknJ1EyRPXB///mw5Op98uy2+f/N3QU1vmVW
+qV/ymvK1bhO5k7XgmYPUcwMZQ+mUu0oYLCR8s5H7V87yD8WuyWDZrSya/PbCc71jYftp+iiT3M2
1ksqYFTw9fBWSWO8jp5FxD8YO91rf1yMeyumKRGmwCSyYsMkckB8gAITzzXprkiZ97uhEqSlkSaD
nt2ozJOdOrqVTZmFAd8Uwxe7l3BWrvtGDeGZ8QRoV+xMv1R0dg0vKf+1/QL7d/Y1P2tj2HlUUAwc
xPSdpKDyf/nxp0RM4mRECATVjvTQCNnLx0K9LRurttqy4YRKYLLmYi+Bq9YHjwyYKe+hlKbiVfGI
l2a1zwee48E6Tup15UoDfopW+oOiSgtSyJ2hWWwUJi+2SRErUy34W8/9JU8mS7U0vnBdzsvf7d0d
ncCjJuJfU9SFmgvcoc2o1NMD15bkKfdal1KUpu1wazlG0YAGWuff6bCftFQ5wOkNeM0TfRcqAJcW
Ozv+GIkwAdBDJQ5JiDW7MEs+6PPmaGC1aKrQQl+85TGgMw71ftXpbP9wGArq8Y9V2MxLhQbC4NGk
XiYpqaMOSfhSFgrfEg1abTFaJvxg2iubgntp0G3Oq7n3+4un5IWB3ziZOp6fJLgmf3Jh+PAng+k1
GoLXC0vfQikA+wgmfNQ1e1m90ymCeu6c0RKvWgxsmhnExZmrDFCHseURYo+rUpFDeVsstI5COWAE
HWaYx8+He/dLPLvc4ku5/LTUPMUwAwYxFLa/sKRm798QUi0/DEVBEdZd7RRUrKOTkv9sQ8J2x6Ot
osImSG7omNy5nFWfYFy5ZYOlynVBQ9ggTbtFU1R5tFUGQirsSp9lnB4IVDc3c1iMJ55RkIWs3Ccn
ccnxyW53PQOSHkPVeaUYq2KVoPetoqm0HSCB7hQ9A5hSCIJdLbhBhBBV9O2nPIMwll5dghLFZxIX
VMmQIeUmrs8SxPB7cyDrFzn4X2pNQFt4iEZxIOhwGthNMy5ZGfkbY+IRRlG/CnYn9rVpDX5UlCIC
irenvkN1krk+h8QJbsiKRVL3By+ITASqwK3gkOzDtX85ejbmrs7rkinXMZwPDHtmWqknMAF2RnAY
1EMeNIlNG5ViQV/aRIJTrccvHqtpBr1k5LUOA7w6WasskS1JxVIAMbWTBYABDtD0+q2WDWJKEyYj
ER263ZT3cHhJnBJ2jUx895+6tvA8ZUYTyrJ9mOYBSwWrVNNOBaIlZirHmUUK4RDHsgBwvczjr4qp
R1MPhdeWbLTNR/apDHMyi4GNBXcYjvbKC1ApzuTeL8RmLY860PwCi2m13herNtDES1zMP11+/vaX
7dxnAf2X7/5b9IZJietMJmg0iWgCF9beI3VH6OqSayNuBxkuHxN/NswxUxR6VDwG/KG2eLSbTcoI
AXz3z5PSDOYg8L8a3KG6ha3WagJ+cowj849yorA0YveAJY/pUORw5kmhGMFqGElalNqQgOM7s2X7
TGnhj9upP3rQvpJ9fsnpPmY+3onrwqewTEsIwJhSd+jRBKiGG5zXLymQXNUasalLE2UJDbV+Jo3b
rfFxYui40QZudYVapen4h/x+a8NsUy3HrXLupPKy/rZEOCynvOOJebvrEfCWHJiDTwSSRoljctbo
7QKMCwAzolb9x1JSwpvdLjLF8Yut6QPQNBSlNiJoJuGjYgt+gghXdbBdM0qUP+2xE9DYT6Zl6ZJ/
DaBdKWjAuSSD+FYBkzA0jiA5NGAsKaazybMBfhFZg0T77c0PNlyoiuJNtKyD3i1jwt/fodBr+lUw
NRjlkI8msAO03ywhwPzk0VUFO4yQBGJkJLWf6J2NoePUCz4dd7O5FnxnSrjtrjv4BQUZU7Nv3kwU
agGTt/ddTFJ8RSgqDWoGts9yP10mgz+Di2RQQXBFSob7uj3R3IX7WQ82VeqbclP0P77tZOi43Qfa
WZ/dPRgF+iB/G2ax8z7brbkn7sYtLqgakRsVFwkbhurLpKhZSucY+EuiYZNCUgDxsqKDceEa+nWU
1fgN64oRzWgujOW6ezt7HRFAqadOOoHdhzhVPfunnHofbcesWZb2mRHuCOCyAQCZltfwu72WB8nK
DWz18JIgjAp5joEJEwZGvSInLQdmeipaAfUp2v+4JVNfqBU3kgqTXe6YceC/RN9DnH7/oCS//D7r
cJpHCOFhmByunxfLqeH7we4Gu2/lVJCTNQv5o+WE87VpzI5eslVm8VhK1DTXyem4LceTv7Qb+FwH
eeg3CWcivPk5VBGIioBCKk3LKbQQdDHAdpWqlgFc/WDlfbK9ugtxW9CiZutI7ng+0SsZZ8S7OJhw
eitiu+P9GM+3kQcQgXG4DxkMp/c0VGpJrTiUNpYBryUi8h2pAOD7CJHIxfYcm1TA9FggIQFYyLMY
OQdGHQHEe2uwPD9xA9vaetoUDmIby/Wgv1KXQSm1ww/+kpVE5kUCtiaG9FuFBcCddHyjLSTtlg/H
C8ILTxk6eGhuHGWwlDKUan+9e9noWIY1/59uL692WKAjuhJcHm/2mo/z7mgo1cst98tMVi6E+n7Y
JrCclQ6orZahTdkAmZybR6IQXSj37NhHutoDKBehPhv/ieVo1cwFGQBlakOQ37fnjVYG5+yXcceW
EyJSuDqw1+Ezlyb4BfYj7LFltiIezbgs+fpnVjcP9rqR5uooMWuM9eTCkm13ILtgFYLQGjKpuqKm
AlbUNnt3zcksJZQVi+fcPoKD3N1JNwhv8OHqfbCw+YBVblwAB8yGfNOOYl4u8THFAqUvxfX3r35m
hY6aKyTl/gjSF6AGgYEFKRRcanK6GNwGzwejOewWRe73c8vMlwqjZQKlF9/6NGWB5c/NUOHHl0p8
e12ZNqEhzAzuzez7cYAEhg32Lh9lL7WGnPP8yM1Cn6v48wXV2zGh4qr2aO7grsSl1zbCjjVYUKwF
NkU+rWvDmdOBdMaJDL4hwjHVwg9Zj8J18EDepZ51NlX6bLYTTmK47sjH2WE/dK8TnUNon+FUaeqc
kL2zqtciEmcBtwNYChsuo/xTXP2T1QGpdVrPPK5BzF8/vSpb58okZbWq6FmsEbAPhtPLrTOYh+c2
fFCLlvlELCrkY+Ay0JvNFcf6hDg4CfYEmKK+UEvN/BTYLwrbG+d9JDeg0mHbSSnc1jsO7Z2Fxksl
BLSm7JkX0oomgKoFpxlLX+x3UvR6nlB+Tmczw/AC9LNNgvtDpdrOMlao1q+oVTZZYw+DIDzvWy5i
CdZhnThTf7HYXxfECopiTmhMZqZbzuYhmAd3TizDxeqFRpSA5t4BcfwhRw2C2tmnIK/zI1zxYaN/
S7ymTJXwsRjQEVr6a+PN5UdhBPKvMt1i6jbsEY10wBtPjSmxkH3KCxcJlL635Kj4SmfaRRxSqZ1T
r5tqbS1XhL9CQrkbI8imqOxElrzuRFBLcOhUwGqNtobeRFabRGefGY1zedYe+bVWUB8aNDKviqm0
IIQHzY+ie3/CEcLapg6a7MzjeVSVQVgjHLJDORyy9Pybx6FcZhpYUBTdWO28zS1Pn7v7tpo3L7oI
3X615MjoBhWvr4ws8ErclI8+vPkqkzhwPsAF17jViXJPhxXJeaEL68Yj7YMrW05JCxNYTWNWQ+e3
vtY6lvokVeoZbSHmQ/dKNrI3NAfnH8nxgxSyEk7o0SwFAnbyY5ZRJbU/YN+eqBMfAWtbi8c9C+S2
BbU0Yv8JxhuN/spBxI57FZYDDm/IAb54m4wBKDPoskFwrCiicle7ylYqGkM16FNsQcJe/Sr0NxSV
I0KiOSZbbo3pAowuwKDTg6GAdPqwOuXVlD1kwuM77WEtGCr29bBwNOKxfvsTleZI0csMmzhE4xfY
vetI9hB00C4ABgEN6YdtbGtCKFSLegU4Da4DkoWCPFCKv9km/Q6wL2HVOb31JopMkyP/l+saGRAO
aX3VvNE0w0MCcAXIY4y5tamJLxgDf3MrJ8BvA7Bz146mZlg9SJJTah9myyOcskNuwvRk+Y6BPkfx
QXDJHXysRMBCUYPhJvAVGgPFFW/I6yFRUSJK1nv+z5hvTysQSlFL2KUrN33vspiLCgkP/E0A1wKH
g6DKxWAqvxuowzG7eml/DbXjP/KWoknKNGAfv1L0+w6ywXZWRWqJtx8DAL4vptRnSoQYj5MDODi5
NligPYF5c0wAbnD+70y8b4UuVRbp6a47pxXH4EL/p0QCA3sshLvxZl/AwqmiVLEwpobcd3sgN3uC
vx9k1B5d8m+DNZp2NM0IhklDF8dDdHuSi0rQeNAPMeMZFrSRZSIATXszzDPZLDvV4FeTorWHsW0V
LKN/5KcldStDGKQmgLZtVIx0sIXE+Z42AsFvfYPm2G7U/CLL0Vkr99KYt4+Z7IHOVqX6dz69Pier
EnXOs/qFVJjU1iF3nx44uRos+5k2NX6a0qeWPFsRhPzXNmZ9fhySrBGzkhYndchXf0Mnqy9UpKdR
+LMcr1Z+sq2/hd6s0IPvhHiMxn9VInMZTCzfTzceBOFWwd1jFqBRdKo9WvhJ0+2SA6/oUwG1SaWX
3tpvyswSf+adBtjW2zRjB6ATs5oRuu7Ku9gd8MAijwv1P8hdt8c/mZHpcTcF0IdnEDkI0QFVAy1Z
0XoCehQBOl5ltPiFHmzoVKXpVKPNwQ3li9ld/zrfVDlySajbzN7WsCEEFoqi98tPTM5KzJJsj3q5
tf3uAc/5M3la3V6LSiuJOg8YLFdQhQ9FQdjGich6VEgWIx2i4q/68YFx/yi+wbsODEqVMf9uETyT
CoYuTy8MhU4I3gYx0XR43m1fsqXi+fpXbwCdB+vy6Yzx6MGo2anG7MSkYXMicjG0R2qF3Fv+dlg/
jGmvgnpYAmcFx0OIKIo3WnD0jps7lR9mVmM3MUUsPIbV7JlfEhsja/QKUkjpRIeICIZYOOmf/Wy1
/qdpQARIeiBVUkBoiZG5JGhSE26KB+m3tV2SquCKicRgkSIZfw2UryXHjT76ztusIbLrnMkAAeLU
xgQ9Tiz3+xsF7sEbdMmE6YlMuJnoSVRw7c5nnbj5a/OYYyjALNI0MlCpXlvfcgOKeqWCNuCWeLve
bC42BFZezqmUinP7oJcO1zeI27mYzebc1n8SshTA5Kyq8araoE0DsDzhrnlv92BCYSVCThKO6uKV
MSrgMkH+yqAXPucwWjOxo3LD5EEfEjt6hOxrq6LZMcHIc0FToN9hMEaTsNqvY3HU7GY4wB1noBcp
a62wWhoYrP0Vb4i+qxew5c4ulUIU0zPBUam6Qw6UDKYp2voz35vNUg2/szicOUNp07g2EHGFYn0A
myqUYNJEGYcZYr90aG3bUrK/w7RH2gt/3/9GQanTdXEg2NVDlQ1FgJTLNDxPQjYnSpVG0GSoT02P
Q46RtpGAz/sDWevCbCkHnqGJlRpMgevNu8B9RgFyD207cVqB/bDLFmYfn2mlZ9my5lAhzGOPxGn2
XhBXW4RBzp2U0ydryxHf1Cnqhn4lr9Mg20vIUgnb5oaRW96q102GWhJ6VmfONpdmInktkP2NZBBW
4K46r5xN3WzSfXUk0WM7FFNSiRaxvFBj/She0Y4C14YbMKyV3HcukQlS+kkpbFW20bsrHif1eQE8
CU2DQADimOpWi8kIVKAMV4l5axrBT9uB/y3DnLhWeksEiPlbpWMxbCgAKDbBOmU1EV1BEFS/bIxw
+SBrMOCZeYmsNl23AU3OBVwqyb9/OxvOcMFLsS6PqD85RWnePLYbHEQTFach8bf4MnxExw2wcgOl
z5yI9gAXs3ciL5+MBdCU+uujwS6DXo1N8tufgzxcEApcvq92Zh8cfenckRBeQqRGLw/MgVzKMX3d
5s0yrezmzmRvXbKJyCJer7mVMI9nFQHdBoolyx1IWROP8BBaY+Rc3CI7vClL6OcKjWqBakZcKYHB
l91MI3mwHE6yI6tch+rsPl7MpYERIBWlVKKE7Y/6kGWX21UeWMWrnAkqwwdBmQ9LAbKGO3+qogzP
+bRhDQsiKoAN3V7DvzoLcyDnKgnf5unyw2I9pg3fFac+AdD/RQzEeBd5aCKQZ2ZYxsFEHWyjl3L0
g7FnC7gaTLxmgsbPb7A5eV5DTqZ1jHKFdDg9x7GzM00OD7KgOb9wfaX34/u8HnOAtOhJy8rGmwEr
sPbSWP7t4dU5wBxrvH0n3FgT2Ji2VJrtOMznG/DUzrJfrKXQymGE0eL0v2qV/ynTsSGpGT8V5vQE
VE690eoovQQs9HNm7Wexgfi5FYsN65x6iWGQekKqRw36aA/qBTcDv9VdDy76rRXguV+KjC2+NXeb
GX4L2WuHEs/Si/UP9h+U6YsFKF5yiarzfNJZxZj59vJF14XZw7UNBhbU4GL9XAzaXsAfz2OyO20e
SPyG6zUqjTkGNy13RM7OCIQc8ZrNUGnh5RSFl+jgoQrJT9g03Msqlcjf4CZ93puWXZWA/ILkqG1Z
9gaWCrJUALWRUU1XdAf7pBHbFGbamGTLeeXh0cBNqVbmyienCn4Z2EJKqB47zbz3TfoxKw/OQPIq
ozWyNciy7kfgdrlm2LfuIAkr0QvTmc4uoHq6RC84qTC+yBJKxVJwlKk5ElQO71gkOdJ0RS1ftOcR
Qjy4AnOiYZLcyb+TtTtxdDMnVwk/2U9eXnaxwLoZzZiQrExSjWo2WvdmCR7EeMIZWX2ZjDSDMc83
CuF9LaSO9sVLGhlMCnn4hy+7QQ0nhQofh/SVekf+a0m3wbX+j3OfLQrPQERNjWjnz7PfHE93dTkm
/QqBOTfLg1mgbUbOBrxaxoUNy3QuxEtppFOhONZgXtM3WZHvaDIeBFWk3FxLGtO8LdD+FwDsMzTx
x5N/Xk6Lx10N1FzYhrKI/Ohqmpit3UhO2vv9KwW8PHF9cStxZAipdJFHNeyKC9UxlLG6zJnFemaV
ILH2vcrHDff7tOFsXgzyTl2Q8q3Fc9EVI92kcfWio/orRHPdcb/yjYoaTLMtNnl7UBRnQIM5fjSw
UXNBy0cFM9YWGhPcjKL/hxiy25a8n9NXLMxbTa+I537/4Vj0GJjj3Dxv/JT5pPp3WwU3d1R7m15i
BRF5dH6bzd6GWy38fHDJ6qdxjQoAZYdP4WYjuevg+5PiCBPPZ2qWbwIU7f1k/xzxUhukjITM2TLi
qG+anCSE5egTTdqiLG8x39ReHb+Ii++XalP332DOzwi+mhcLYGZx3SrTl9bgkH9BH07b32javGn2
9tCJ2Nb11AwH7HeOgKGtEN4t9iLtelyWW2l6W7zBmYH5nKItFfzK0aFk82pXg7M/ZW8VQwrX0ojz
HCTKrJI7Lwlr8IR/eQn9bXwdbofIO+yjrfF8YjHswzoJlUsWJhbXcxhc7W+AEgNRFvDANe9pxYQH
fy3CtBkyWRkL49v+jrM4s6ZGn1YekN0Dn7Fyj0yAaDY9HMwiTInJ3bwSc+xqFh0kOcV4n35jk1tC
voLwSuyGGXK0m7gH9t3TEL3FEsVq9O7U6DGm5EoZzpBbSGPmEYJzENfdKGaeCX1ey1GeHuA5Nej9
5wAzRN3kwPPFXl9n2pD3H19iRQPK3TT68gfs4Hdb/YYoeh68rddmIIq0NJIN8tNNdJgj0myDjTT+
hTpOnM2TQAxEUFLB6gfemAcK2yMZHcY/1AoWJCdVGDqnSM0xpsckxPKwt+ZoAXRndFk5QwV6Tsj+
5H2UyfN+qf5ymFaW6nhKsQ2JrOY7q5yApPLctkBiqOc0Wz42WcrkapdTEJgZEYyhUYS8eRNNV/+t
en2iSOVzqJdEl4bkomCbvImHEk1l3PB8JZaWAcK106cCoq0IkwqPwrydzy2XroCpmvxkT0OHvCKK
12WI/QAdlntIbsUmZPpy2srJtWh7ui9kBFm4/Kf8zRZCgFTwUK2PklFoWRIZM2aIYv5vOpPgynOm
eIr6KYH0PKO2bCEAGMZ5bes/1shiawgvpUUqzuP6RcvWlJqMeaS2G+fLZc4AYQ8t7+t3encLIdZz
SPwSYbbmJOMgmq0XiKjz1SVnxSvKKC/67pIZyr865YphiohO7CFDsfq6YKtFPJTaT7rKubMxo9V/
Vm0UO6uDnl9gVP4/A7B5AFFmwy/R2TRdTky+KOOk37XzvRgavoU/Z75Cn6dr4xAnNaeSbs9BUsBl
escmfp3zUM661kcDidxIlYUWlsWRw1Cfeus9MkwXZ2DFxwqaezdjaW2m+Arq6o91SmDhWyT3jbU4
IhKJGCI+e+T4e6muT+MN5gpfDhY+vspJk9VcCNRUpfGoHEg/wtCY7kY5uxY/5c5DV+euSTsJervU
rdFGBOL3f28HxqTOyp9ZTlS/E/qqaguZhsJzCGFpvJpNA2zf//ML82mXPZYgUEl4oJDD1DItHd07
obuYvyiyVQzsHB7cqKrOQ5hpe6chFW/qJ3/5d0BhWU3UR4WeLVCAKnMDb6bXAznQdEaqJB/1+th1
dOEe7HBr7m4sk1Bu42PrG2SOzOZiFLWohYxBT8WjKh76k9e61S+wi1FYmurKNj0hNnUSldzLBQ/X
88S9mz6dKd0UcvtG3F0/hSeqtQRO9K/1nbMviuGLIG7F90JdjuZdErWBuzXt7JuqJjYUXa8+0WGN
pd9gtcSw4bzst0TkgFe6bgj18vQmoQv/qKVuWRZDaPxNj7TMMA2JKWbh4QwTmdqwEGPJtaGgfkrY
Ur6O0HMXOZW3OqQsUZKiLEYOr5wpao8pBl+o5TzTkratb8ANtgtN3cMHohu3i2uAjaNdRnIfeIMW
kGL64ox9PmIXpHTOOdtrLuzWmG4pczbVzwqBGQBSNRueab4oL7+XOIEYPLle4h9c7XWyhiQtl2nX
dcNcFwrL2xOZM2u2SzRqh6flbppJiaQhlYaOKTwiWOQH5VmT7QgMqW13hSE8To7wjdZAYAJAt5Up
/F7mms15cIV1trVDomDW1SuN7prBzuBBcKMJUptR6yGnXof2mr0HFQiDDx4fpxhUCYLMYDL9T9Tr
OTWRQC9k6qsVQyO396JB/zo0A5coACPpoij+unUZlaC5NAvajLez4BOqoi2fL86opzgJsnE3ZfmG
4NBQhsX3BADTEQDEsJ+xQLLZlNmE3rhmlW7rjvTHire7LqrE+wcdxJoyRbOm5+0ZtbVtMK0csDQF
xGp6hywz+19SeMifEr3nEbL6NTohQIDtxy69P7T1qI8XOz2TAqD51Jjz84rVB3cJVDcFXx2b2hJs
y0Z0IfcOOgssqm2zgMBnperqcSMhMG0ozt/N3ND7bMcgxRomWigW5alOkdKDHKmmpWviiPO9h6ZU
xj0Y8me593eUmEHTZ9+dGweh+2v1Po0GsD0p++TWHRDmNFSC03G0G0wZeT4SZVyxsw8WAjL9VfuU
qSmXiZ0HkXr/rqAXUq7ZoXYG0vC3F8OTMKhDqplPPk4EZaCXlESv3Tbn+LQdupQkzLPxSD8BqBHi
SqXEl7nHhCSKYObdliY1CkGQFogJ0/Tiaebm9HL3JcTwYaHl/L4WV8aIJislPH13QK6EpydxHmyp
ejf2uijuAVOvb7vsXkhZbqdHms9O2YdeMOoyJaV2FEQiBqqW1cWWkxJYmyRIro3gS1KUzAgTbSTe
uKe5NEWrAHM8ranOtmw693CJ2iGLAEJqmJaOWfQsOdA4/Cvroesc5w9H+TsFj/UNwh9yrHe84R8W
gj7cxXGB3LjfqsJqGd4fIYsIR2QZTqC3gMg7qtptoel8BmE8BtGCrayV7qV/wl3uzkzz6Q8tprzm
TWwHxqGIuLoiqzqVF31DR4JeqhV7u1G3O9+HNFrwewW3PjkknMSh/87HZS3J63jZfTrl0/qt3iAL
Q45lit33MhplrTRPCh4H7Pyb8FsFFT9VLg+Ka/WwGDNQatik7OEVe/zcobGHr/FDGOV0+TUFCmZp
/H01bGQOU8ySWfUY6WaRYrOWyJgvQVHrtBAZY+ygSHNV8nNxnm5BxByMRFZbs5KgcduA+zQcjdfn
1aatDWttvLxjTKR7/y6kDElMirP1WiOPZ0Bq+aGqUfITm9/iC0iTQRFqkDFTjWu3dXjWZzBEFGkZ
0T7KN4vMS6kQROjCjihuyZSrgFbQqRy8sEGIK+E9D6BoTigVuiFh/fTHhcK0V0k6a49BdOSR+P2X
6NMfoR1mEDj++YIaNk2yxvJ0hXg71UvzLZvSwwLVCYLNxO8k0Pa1dYiPw4xLXwpWsPFjySVoHBiL
UKU4ZSayUm4/1nL9wwTcowdvQzKx2gnI4JOKeuR9bYNPUZIaQf7L2+15Syk67Fl+RRzWxnQB26R+
hCzvCE15lQgy8GRH6gS4JdlUgVA+GvzvwRM2GQ0uk8pBUOnf5obC9KpoVdE9+IRuzB5jv1q3YZQ2
hjRaGoaQ3fzBH1EI2s2TaisC3Idxcp0CsHK7QZ3NY0Jq0WswDAAQ91hlndLzveD+mBsEx6u7JaY2
MdiyHeTbwEWgoSScT4Pdon7UEbWiDfakvbW2AM8txkz6u40Jfj1wIwARaESD9UuCgGAbTn1mb1Ij
eCgXHLRZN2sB7bz3u2KregtMqYzK9Z3Ko+h0E8XaWecqRnyiGKHoXawSlM9OywPKnON19dbaLAgh
bRDLUDka1QODVaFrQE7O548IVlNC+zKbLEG/vX3XqYnFVBs7TYUY+R/ox5rSVrcNay4Al7anakbB
H9YQUK8ycvam2CwxsktJwC2G04UrRSSeIeEppd/Q3fKeUyZiEPDpYHJRI9aZ5Qb98ekadwCJ1iTq
BZ0VRwShv72PiYdnkiXaNZFMHUUiskj18CuuQ6OPe/9KPlcF+GvJZfQcIgbMzOa+ZmWPx7X9yUW7
HJxJClJpuy/jVFUWKTjuFIUjl6C7yajz9KyzpxHZOryZrBqzy9124IJ+Ybjbq6afRp5EZBCsWRYP
gp222zYF2oePS98ZnkqntIvy0m3ROgQsRwIZ8VG4P9viOBk3xrBhsfGZ3eX9vyvLww2e+JJdYqlQ
PY7VXQTaiZzGWJuH3qkDTcIb/6R3gqADspoQlewYs020Gdoo+HGI9gj4tmO6v7GvajxPNxe1X5fo
GNiFhS4mc8FTr9niAgUn8u3Bn9v0ilk9hRh6FRk3ww1w6MoRr8D9aeFcGySsBBW5GuIW+Ayflzt/
H+xE5Iy3qOInwTJSeN+Ayr6RjASqlI8Lr6+TrmZy/AKFmCL4D4q030Y2hSksTa9fM9UawsjslWWT
5m4hDrQvvqJ4+FPUHEPmudzITUBOqY6HxTX2um0mfx8mccWyKRv0Tp/E9HLjwslu/FrIKlykyfzg
wRiYeIcL2mCGPjXof4KVLBflGVZrvGbJ8yeRaD6gmLVE7Z/NHvuz5zx2pgOerNkY4RbTUJpgtv8U
O3iTSbB1leMZa+nqxeb2q8nEA1T+2ZuuwKh/WgT/Oy9v150AbuK8wO77LXKgAMiDgdVqMFN1xrpy
4gfKg2zkF6ANQDn62QIC6O4+/nsJQg0CI9gv2yfH99ev8WKv6YBoawbbXLcYI5hV9iGj+pB0mHkV
pFI4KTdq+A5KXL+HWAIveE4eJOr4AbhZm+rpMpQ+cxIBhwGQOYdin+S5RyCI/IhCx0FGXY+vrank
xIvoJA9fzU8C6b7tutyBuiB1XtbyUOBXYCkACNEsZ8d3b10TYSLrniCJN0XctwKK+ZZ8EE6O9dtX
b/SJOSIzFxVvdgl0lan0npcNQPcBAjDnp1c8oXTSxwpSUjd7ft3qbMpTXpqDEgXEA4ptvM6Y0HFv
w73iPTHykz0v/TTnSjuJPw+x+UI4gxv8h7YMyOMJHOH7QHODkBnqxbg80AMajom7O8gMdC/pwoWL
8/UugdRamgaAQ01sCLQ3SuQl887w6+7aXfzlQKlqOK59MMqg+sRuJLbErPEmWJy9NEBN6c7YG5lv
G1LvbZXXyQl+JukNPIq3bbRR06a6IRx6Et8bDmQ1Wk0vuJ/XjL8Dn6/bFIhCLdMTYJVQhNZi8nWo
fKAxqZmeeeZ0T9NAakCqVcR+TDGIN3PDUZi6dSkW3XRB75y59dykoTIZlAqxiCuWGe4SJIrELyht
YzMQ184mK5AnTY1LaCD+GCtm85YJOM1yvyC+E2PXJNz4N3V8AFFOGqeH6+iWCDOP1G3mRAFT6xPr
l+Kfdbwa7DHfh6MOdnuq3Hl6Ra5sJBIQ0INGvOkyEMi15PalsOnYGf82SOa/tfQk1uELWcNpWIFs
GwbazqknJ578LU8UDH7pXhcajgCMpMzJG49+S2563ODxLINkJObr1Bu0csY/p5pbfBIiX44UlOvi
NKDgFvqvpRTf9WAmJgIjp1wIXohzADEDLnzpArE8c/2TNme4ncyu0APyg1b418NW/BTfXiX6GjuD
P7GxVZBGk8TS/4s2d0vZO4dSbiCAsSSScWAnPZol7NCuEGlwKrzWftRx+d8KBZrMK4BID+BSbRTZ
4UPDzWzmsU57d39Ioq0i771PkA/Pi8vjC9tSFFy5ZIMLfmCp6w0/kwKJtCvpsjkTnZLnRGWVUBuh
ZNLigwJt/PFh4k16qU9lR1CGyKvBqntKM7h3102CAUQyTbLK++mF9pHSic5Kx+Z+UEWKNBaxwiLB
i/udYlLwKXEdW4TOQpwqiMmbvzPTJ+g+/K5DsDeoC41pLbgL8Evdoj5YREqyBI3RgtaId1PxgpVQ
uXwPVOWp02dDoShog0dQYg0C3Bgnu6xZihwv0+eDZrHkmeZxvPWD1iDNl1a5N2XoO/y/BLPLEJ0r
Tk55JZ3DVz+bq2Aj5eRM9aAGazFcA+LUFeqDqGda8usWawD8Q2eAlfFU4/WWbRbO39oONJUXcyVi
NFX31TjDH2FnjFh4LIVzyaoAIVEggBKS/+MxcPvXLq+334QCZjfiJd9YI4pJesSypORGLoV/YAWc
7wY/PJlV4NO1ZDbylXeImeQPRQ6MWuciSOE6hSmRDN0ssfaN1gkXlEoXJNZ5kWFFoHmLWIPH4mgL
u8PlqmCp5MI2nVanNv2SPW7KjOUaAdJQg8cLSs0hKH5M8gf0nse/7Bs+7Ti2Ip+R5p6WKEgtyG6h
3xgQHy945OJ4Kg2bkmhUZLYq2wS/mJd8/NkQkYlNMJCSGIaofwvbHGzGEvHIke05PpXo3g68/g1x
02zZ1oEc9pjlH1dpJJlCxtY5V9SL+MFqVneadxErM0twI20mSXK4YU4289VdaRMrDj5nni2iY2y7
mwkAtUDmk1ijp6UwGJXIGMb4yDSGxpl15i168fUadNdd/6+UH93bvhwXeYc9jLuRclpwFZRUIh2V
1R4OHPZIG4BfGl8W1vsH2qnDqbsi+Dk1yp3sUkOoGEJhLARCico4zM6Fts5l6u7QPI6K/L64bFUp
RltewccERWPgSWllebqgZaA5ppDP07ecCBMc37jGkKamphsyeAcGQM0jAztX9a5Dnu6bzswCqsR4
akFIXRy+T5UNdB3HW7MUqLgp43tUopMhB51LcTkbzWse8edSuvRZNXJR5eDN3TpvhOXBrplDTDXa
63G0vzVVriopTwF7qwuO+enntDnNeXH2wbRSzpxWaMuEE78ibSPSSweqQMiwhABep9P+nkrq7rUD
r/xHobQlYfM0J2gMJ3e9OPOlHx4TymCkNoUNqo7dUZEuJ9Ct3P/GMXo/U350Ohgk1xs9cHeaTxKL
qByjCNZmcUl3BtSzceqqYuTBgkdfcIMijveOgT865VRWEs0dJ3FVpTYtlOwVIsdc9oyTiy+5p7+P
uVBEatXCYZIfbliE+xSwzco146UagP64LP9BER5DsE1ttOv4lVHUIURbXYoKqPueysOkChQJl2uX
idtDgH3eCKIw8GaLWx6w5digtlKXbVRpQiQ7NGhKis+baRl7OdXG1BQKwevFccs/ldATgkm3wj8y
otdt8CSzcPzQ2goQP2tOX9R8NUUV7REiwM4ValJCIf6SMpDHj3UEd0itiMmgjtGRiw/jc1iYgMFJ
DnUOb/jVe7SZHiQPlmaenbWzfPUlFo/Wd7r8LwLnbXHjtPs90Zzcqf78ot4D+Y5/cM8z8PPQuddl
AYimkSUyjmOOT4r7uftI7FxARFsUxctDlejP4FCU+LwlDO0dF5UzsEAsn6iALdhEzlZrh9/7/TIG
xE5fvu8ZfpqnOZ86ZcDcfpYZA+FWdPsbWFEwXzwJ32EnkE6uT2iqx1t8sKsG4Jukp76gdZxKhaPc
iGbr2lqjUnfPUZW1duwyMHqfk/Ym0RdGGoBdhpOf6nb30qU6BLa3kpkFn3YPtX6r5EEZ0hAykmBD
c6qq5Pb6x/XP1oiqMTr/4U7NJiUbQ89MFoMV8Lnch+RGnYfwzIlMNqCL1Whkx6r6zb7YUD6ewZLk
8oDClr8UD9mC2eprs6sSYsOqHLNjjnPHsDPn04WaLXl2r3nwwXn05z9XU6eck8HpvsLWE00dZfL2
NbzFp1CRWH5mp1ZvA3/tfnj3RCo7/0QYbgoRERybcLHUJnGQpBNhnACjLSk5AqeXQL6AY2L7quMk
tl4lG9K8HfEdsITQ8jxwJWzG+t3k4+JP3mXBywLXzbJeSRsFLniOaPmxtg5V6rCEBnpzjexfDPoB
H2z4oZ9+lMsQRB0+gYXrg49aZQaf5zSN2zgo4RTWy/HeU8WH6cpARH3x88c4TSjDuXTZ3nLWOEQt
7KIFQ4jIXL/ql0FKKYxNly9a3XgmpPjMogTcP0FejgOeez0AsZAzSutrfzMOgqr8Ak9D/zoPEKvG
qXS8Y1NXKNRefc96a/Qzt47wZWGNAFZ/olOgFuud+577c/hwGK80N9DQRzTxXEmWqzdqCafDiAlB
liGT9bpo6wzeN0q73BxGIvlHXx+YSOdoMoSOeZlfFNclmCa+EPZdHECIC0ctSjfjRYdoKJYXfJBQ
JJYr8mvFOYqwsHsBB1HuBA/5Yb6AEZloEyjC5BX7bLQjwZQzR65bZQ8Fp57Eyiigjt5POjyYj48l
jHF2DOLDWg4e95wXYflu8SxtO8Fb0iPyi28GizKx+Eavutvak6pAM8ceKj8NcB7R/JvoV9lQSFKC
mcF1WEzFcfd6QAdXvUOYuLF36ltkG7dqZRLMBvAkpzgVzHq5bF5aqLJbfoD5YyJptPwLJW5QOZ0q
kt5vDCxkmztzeZq3rOUHNlMXOYf00suDajhf7K7+pTNDq/FcxWRhyTp0W+DXfVy0D2Raej0vKwXj
dgPJ6rQ//HHwaA6f/m+5CWxST5oxzZY0t26bfDwCqk3rZ1lrt0AHOSReGNm7zuYMNZK6hqRYNHj0
ACT7r9NpOVJE0hR3gBCXMSZkJ3IKDZzmhHgH4mv/zOrv6KbAsayFG9y/z79O6D2Vv+hxtWHmtxKV
PrXqibEpOUPd8e98EtiJUl0dhRv85BcFRYCig9b2Soq2LqnWQNNngPO4D25KP0p6zetfjoHbprd3
thiC233Vkrx3ipoOtGKtqiy7qFoTJExfugy6nSl5K6Iw4/8C32DXiDD25t7xvID68Oa8btOEDm1m
VI0LbZHW/JuCGuEyZ6kOTnL7G9xqKGWOTTJDAQmN+w/YS+8rU+32goDG/P9WcqI8aak6PkVbtVNB
WkIpX+hm9scm/xPX+CcPMrhbg92uM/VdFJ+NGGktiUD92iBJWU5eadFr809WmmqJHIZvsjAPqS/2
6OXP8fsJ5u8ROuAuTzyjIX61EvdZ8Pq3pVb4CSoxjezeTi9kMDDZYbf5Z5tnxUEbQFg6sbSzip9w
/bp2Tf9+Dk6izOXLK33jzoKSxbcUqWtSiqU8VNiRVqZgpyg/Fbyzzldb4o6awvqJCxgvM+skfDbC
PQEWIDjj2BBEYRLsBG5cDiajegztKj/K4j1peQQ0wkjfr1SjT6SB3f69pG/VhjR9nFEs1VuwyFIG
UDY/OLUBK4IYJ+IAw4M8e49zE6dCsJesLfImFsG7mQm57q9oWZllD+NcqOAWB7ygJJRThqOISL7x
VekpzkM+ZpzgNm2LeplmOQNofgfNL8W+ewwdXoNSbFvqDdfrHFSi7Vnh1lHDrvgcVThYIaTxzzIj
9tKarGdFN8PWqCNMPS9Lz570XdAaOPdJ5zZDDmkQHqOPeR3cZpE8VzzkI5H2IlK1M0QRI5TbGE+u
YKTPs+2+jyuWTsxU8P+zQFzv3yTt0y4UGPI53rlvuJFYmrBL/4JEJiNKaj8Hjd+mva4yysyz26VS
PAkvslkMmQIkRlggyEc7j6ruLacelFGpkgUHKVAll+gtiRe095yVi5z5yjDn2FPhyqBoBVw2/bOr
OhDWkdzLxy1UN5FK5h9rk3w6zFCdW8PClwculEMTrLSF2QoHfXRxRItZJ5PoM5GCkKFN5/p41BNQ
PU7zUBjf3Bc6YyQ46E0hVqOzH26dbhO6au66kkp469zU2W6DwgiHzAvsO8kjZrPohiwMz6TX0lb3
E2tobpu0cFndn4UYM89AN6RsT57lt05cVT9sesSrtct9hKbDL1cSLkMmAmVAKIEn0m8G4aEdipod
KYnigtj6OikMWYdS3mnHRB4tZS037oN/fVqdPK2OJjxZoTAlXMMezE9rRUhsMa06YvkxAvgUTxS8
wIDnZrHx8NHhDWva+8E6NQ8fEzqXdEGjDR8965bU4k6JZmFyoXzN9ZT4jmPlvsQnzvxiAlRuDCZn
LIs6e55ZmVmMY+PDmUXLcatSfARBuzoquBY4OefYppH1ArtUy00DYoPbnHgiyVCremxqNeVTR+ss
dlThwnwNPlc7slmbs+nhi2uzCxbBrPtL8xcAW4fU7lenbf6cK0qmfcloQHRT8M/K66ybgoa5mf1P
3igf01Sh5CUb/O8YnCIf41mh1NDJF2XSTuO9rCybuJRtLgiLPy1ZvMasHUMDpShpfFaTE8ReaTr4
A5bwj8jr5lOHp3jIzq4K1GnNXEc9WICRqrP0JIcbXvanrKH+kWnC/ST43Lk+JmvuV6VWe5CGanp+
f+qU5fvn2Cci6MNX5AhiIwc21BfXhl5pHJ/yKf4nydN499hj/Sy7NZYLsgbJ5pjF7Orh/8vC5wEc
0LNstjx5rtNMa9kO2b1UUtxb6w/VPYANSN5g6mbMKqflf2VOyt2EeYxKfG3MBHvaA38LEQKctXN2
WDgE+wO5huIAiYC3wWxKIxMFynapzjCPyQSps20t3JaxwlxHySd4fpqCNKzTP73cJiJm25aoMUJO
QOikq/m5GGy3dgqoJAZbtXIHOc3yvEF7ee+ibJzjrbMb9T1tI5/1tCjvvKnHcYr1zdLDvVgGITbd
a4q2/BxxoIwj6z3+4ByidTKT/7tvdsk27i0TnfENEdlZVJ838SMmz+XI1mEgaajroCFFE+K2rXv5
0BCVj/GjZ5Cn3Xq5FXlr7h1Gm9yWLfyiYEol/NYtEoqWRAIsRyFIhiGdbz/dq86ij68agbAbfg81
+OkPHsffJ+oTFOYjTAoKxD927wBTp6gpQqU2EJp947WPWj6eaHoQO/WhD/04OFv555c4evuGGZY2
6dKEtGlotfr/XhoXxYIKm58j4rblC9ajkfKxmOjSqJEX4+Vk1Ed+n8Os5ZQKp3bGCnt5bumG8K8Z
rB5nP14Y1tF/FIToTlyWhqXErEjG5e6ka1hAr9wa4BerpcPHQWxsco/+I9Xj+2vfNKSN1dLQAOk8
vRu6SznWcVwEaoRf3SM2c2s0AV8dw2i4nEyDuaDMTbrK5bn2AwupZ2uEIpoTKOJUxW+6BWzkjX6q
U9ALlX07emPXAu/ZnNq+jskbV8hoOAcLrZJWGwPGygafil3fh3n2n1aI0wAxRrUTMUAqqfzFEep7
T3hnirbBW4SwGEzvd3K11YCIp5x0aq1BLDekkg2h5+OokemHcfeUIYJCdRfwJeGgpmoL0F/rtoP0
35g35B9RZsipfAR+a9n9RnIz5TAM6UlNL5l3IjcWXLi16Sf2XFVK+HXKB15gJsOvoNzDtpsp5WtN
RuQ+O5nGZD+/Y6hk5ThbZwQ+FbcXSubsBmuXdjgOfZRoiATi79RzVf23v4IVPpXrAj54Qvdmo/MB
w8Qn8/fVkl/1+PvOpwg2jEVCqllkM+nFiDpPO1zQ5d9krYs6KZywd3GVGUZOVtlpY3UDFg16B86O
YrjILdeBhKXEvG5jOun3xin4Lu1q4Z9og97X79KGLgFgrY06WD+jPKw2nrwIGQGtOqYxY5He8G5h
dgUTKWi44GRead+ILmcJJaPA+iZmEZDNKHTjkDWIlozkyqOGIx9OJ0vvIoWX5UmTcWqhwWMiOmey
WE2P86Z9hu4BVYbun+LmBFUdCKYWpxdHOQt84AcOawCgh5oD2wxfhKgS7enjGMoOpfyHZq7W7LyD
b0CPvdwEfD9FmcUBP8r4qQ5ZP/zzZPG48dbJSZssDpy351ebURtkiZecyBy+TInY88DohxaGLfYL
Cb3KfdPOFxxS7j433mEu2Z2iMMjfcg54JlL/dpHtsxLEhCVujEvofMAPGDgl17D7KHc1q5OnD4PV
S7Y09Xm9mQDWSmCkOvbqwbJ6H3H1pDakvHG9huMONeAXr803KpUSv00Pc5gLhuCPcPf4ObRq3PJj
FiqOhHZsfk0hmfEe1rnS3dPw8Y78IjP+dlX4grgz+x+fwN5GJ+wXvRXCKyzLIpU2bcyGjH0zy8yN
uF/wMB2P8Z6BU5ffv4MqfD1B1D8WLc/KA8o3p2ULbELv2mxrXelFS2N+EOdpa2Ill+MgU1X3uxKy
SsXb4uV7dqUHgrjDv8RvPOsG2WJsBZZHKrOfuIZyU/DNckxLgaziu+mSIBRtD1USRRcFA1vb1egp
lgybgX7hCXyQny0ZvoXBCku+CzzUQ7XBHPgaf5qWxgTw6qn2vI5hdCZWz8IK+RHVwORPIfq+ER9a
iQ7x5WkzZsTk6GNiBY8KC8+2g20KzLnx6LB9g1mGlkMCwpayZj5MFxsdMiHL4reEm0JSeQNXasEu
cKj7sTMJ7oJ29eGOVrIj7CnktnISCLz0+O6ZHTOiJ0ywhonb6tbL0dZHrhEyj8QJ9FoYxeziX+QZ
MO5Rrgk+9THMDvTy4Cr7N5GxhXjiVLvKtIBnv09LT3voir4VDUqz/P2sh+WOky+Uq3FuSp9nt+80
kMwm1gaiC/ieGiQUzpyoMM46PltUlMXS9o95s5zq5a4XCWsKvAx0+TaNRcyupyWjYMKHItbyt26A
UOOgic8nD0HDWdSAZo4pUph9zvB1xi4xW9wVd4KzTMafr4Um1aVP7NJAT35NR0QJHjp+lmo0hbkS
q0jBrlG5A11yQj36dW6GqWkl0Ujje0CzrDp5ihUUEcGnUlPisRcYCKgUWc093D4UTPYiuuhnjE6z
+TBxOTIydPwTZo0ZpudFyc8LEBDl3Jas1GHU7U80Lgv2RNqs1T0P7A9NJrxWKnQDk5AnRQL73xRF
LEwpxThbDu71TplcdGtR8GfW9zcOJNOqBVZSZ49tAldzG4p4KzDWmsjL8y2lfOqM3bKr9ezO5krr
0Lj04SEDx0EOdTikfOKQ1vP/csbErdMh0myuhPNihO7qBoSVR9xSAVuKdtRN7b/kZrQg8dtUktgU
YAgCgcg5TZmHdBAL7M8PhtzS0pWEathLR0TDHSiojqG5JDdNAdP4eI3hvi1rzyDew6qLOQsxiroD
GirAYjKq3qDqkBcPE4PnuYAdGfZ+i27sbP//S0dbjEw5jpuSXLsoD0r9+m6+yX+8eQOrvNwAh5P1
adzJf0xKaMsoGznbguhPSNRLJ87w8IMLsZ1reZM3efzljJwFlc0zDdwM2y/AwjeH/aPMSompJo9I
EYNa4L0gBGkaI93WT3kqto8tH3tD2p9cBRdM2b60ih+Y46oONSxG1TwS4uUeDv7+ELqTHQLnhHCX
FjTHcxnn/ZwrRNvvGStMt7k/mRA18RCQmhrm08wB/DV5l3Dz9SxS62jAOwbOY/hg79FLwmv/doJW
8Y13TSlnju4F6nnQ2ABEsqt0QocZnWZLB7ZdZJ6nXDi+ghJY5X/EvemBRXBBdZDoFwn/cKOZva58
DpogyyNmOsm3nrXVq+FXnXfgAnjBBmkEYDM8M98pha1VlCvcyStNyVbRRltvJsAg4Fgq139zP230
6DW6BDkU6TSNgNcNGzMa+y8W3XajmeZP+ZiNJ3wY+IMf39OID4N4z27YrwWbPAColJAGRHIpBCxW
f2wJGapFKefMu92TWk8JKYn9ZxK48E9NVlNt+1uUPP5CnyM035CzC5LZ7/Wreb2oshCXxDJKDaIh
qN3BI37tkQLerNsfVzq5T63c5XQMGaT0IMmc3q8NA74ujgM8g+hUDQ/7CADHkxR61w53tGVsP690
RSTjcXf0GpxbWEWHO73evdozH5crIkNTBbE6+ied9CmKKTLrB79IKa8rZ7Jynh0SJ/nJHkhLYoJo
oXuvzPNsXfmIQXpWir1PntRcaLL7ThIcyp/GiqLTztd/QXalT4+LM+Stw8ReZKHbbi+gwWbz2yRU
oLlIBtwezXr2sVRqBWyXQ4Fz3Y2gA1LsTIObPnI9SBgM7Spg5b5nVgno/26Ozeu6Oe1+1z3j50Hj
PYW1zFmAtnKJwmzPvC2tXHeof/92oB7x/Hbksa4Vnxy5b7O7O9ArBySlv5sXoBeJSM10zeUf4LRy
xv+J+zXmEwCbB899YGa+UwcsWKsvLRnePWFYyVNjYJRfIg+ytt7p3r2ZxK4MXyLt+tJ+3UVagxBQ
5I/RavtXcNyZtGxvfs8Trgicq1LuITBCw+jnOr7/GhxuBaVldHk86ts4rGCT5AEgR2Q+KLp1OYmV
3Vz1BZgisEUHuVV3E0lxgFCJPqjD5K3Ku5HW+PJV/vXSzyfj+9i6vC3EPJA8PVRfDLRhaE2a3UX2
1vQADcEQXnV3EjAGlL/4jZfHaAnJmLHRvLyv1U62guxJkYBaSVzjLwK6nI6/eFavRh78uaD37/GM
YTnD+dIPmLg1afYxH49cv/bN4ohxoJrS5u6GGhXZUqZZLzo2cREXf0UbDrcPvSBqLGfSdI/h7yFW
tbj9Ceq8o8Co24bFN26UVwPbVTvRdYcEsTu1bOEjRarpp69hNY8VcwCOjg5D4RTD2qyY3aQhUbHJ
zsi9I2V6nODSGVieeBGlmr7yIFnPf6DbAEKEuqkA19W808EMHo1XeyK4P/hmpEQQNoW7cMa7RIqD
Xe0v6Fwrb4uLUKqlHlskkQ+wAhZnV0p/+u/l/XNL66NXlXz/PzD+Hairy4mZ0Xuks+lNvQP/iyeH
kCf+VP0COeIm04Yz6boCREW9/VDPyU9/J2mM89NWjaI+JxR7qJfq8ONxKiMSxfegfJt3BLt+IV+A
EuJSjt/4Fpj+9ypDtZb3ezzpIuatv4Gd6b5Cg9GVIagyypREOsvoRS3L5Ci/mG9DBu4K/ZjNbyAD
KhemzwKpFV513XdfgYWW284disJURt1p34tZ6DM2bchoQMGKRiE9k3eDkHo5m7L4H6yAyUqiuyTg
+Xcq56lic+g3UPJ4Iku6ocbB4QQr7RnLOKmyycANXQdkoxQB6IH3caWJSwc0H1iAw6qIMIe1UZvO
ym7hmR0qZW4DbO4+HQqF56GUadITlw7RnfHdqDenNP4UJsiJWICHRtjLKMabqdGf23uAR9Dq6gBX
afhjXIqNJuLH036WxqU16WQ5WHQvMC+4T9cMax9qMnVZyycT9GCxSujX0rDurgBCQQf9EQDNuXxp
4g9k32dPVH/CgncIbNJ9ea2oPJaBX5yXZRoSJqtez+R+Hi/ZSb8gyAIeI9waQRXgi8LB5erextXw
j+2eK0c4+Qe4+s3U6UJnqaT2QYrhBbJNCGyIhyjSUjx9dEGDWWsXANMWcUd+dhEN2sN2ztlRojDa
4Rq0BOhCe8PzRdMteVvf6SWWp7K3vkn6BNtvt95zmAlBbE+9arJv84M3c4Rv/sHIF6sTEFR3PCs3
uCNcIgIdKNvfd213YendudmVnwii8EJn7ebb9pgE1Pt3PALU+75l7jyoL0xR4c/oRvV7YeBGj5LX
6ix/uroq6p9Ou/wNv11z4Bzq+HYXmC8c97AG7ppfRBbFMiasJwWrN+x/LC+Y5GHdG4nRI3axK+So
CFmLBgBm3eLkh11250znXeH9h9ohajV13Pm8ReaA4YgANrkKhENoteKL6Aoa8LlM5FsAdEL/e2XT
XHeS/G5Z3S0vuvyF1DvbEh/WPnZbS7IssFSELGl6VZhg/SBb4l01eBFXCpPE3Y8xhjgKwNRDdwDD
kIiRI+v1YYGBYXldtAAYEEfTcR4yr17fFfXXRjuFCx3rEe0ZWtxIM9fek0AaFa8xDZTEkzA4I0aP
9fEByYw06PARdQ39E2CsrwjsMT9Mt5A+GPZj/K6c7NhRa52UAvRwDpBy/jRlx+ru9AWrsz1d3Acp
gOt38YR9HOlmVXfPmrSxZyfadHmGQImd4RoVShYZbvGE3VaiZxB5ncB74vg0Zm1C97sgsdSaeyOl
yPh0F83NOp2TSblorudou4C2jSycGHaqwqRq7PF4MxIQjoqTKo2KsVycFuCkk1HVWslYTnVW717S
0xZRPxxI3XlkQy/Fd6OzQTm9NlGGbxuZIuTFpFr1X/PXGGLD0FUrkISwqlTkgovyPZYr6WlgDsEr
R4TYZOCCqwQXsrb1hlBYBXASXOe7h4VK1siFzQe2UUoHiRBoFJFNwK0KBWWgXxIylEqDR6Sez1sm
OS8ROl+MrG0RoXKdTW7a6IeF0mxPu8Rb6519RT0nPClfUg8LcNq1GUSTTWDKDLqUAq6duRRAjmmd
C6gnLjbMecOfxxICB3JU8egXsqqCiW/Gy9tlpRr7GsjBLU3W4DxtH/35647H8mXVWS7fg3V6H/JI
1INy+W+CU0i878rmVb/3iTqy26Qalb1KQsmcnlHaT6NGMFBfjdFrjbUGWx1Z5yx0Kbo5p/Ox9byG
8h/l817Eea3wxqdp9ACITRltPzyaWFL39I4OWwmyj6DuEomOfZrSVYMNZ8xknzLRfzptJ66eUOWj
bixT3zaq6oPrzsb/hjkjGNFI/ZM5TyBgGZ6nM3yG4Otdwxi9RNBLBJ4sHQL6C7SIY4K6hjeTns2X
fLXFT/1pnuC6VGaJF9r8dachIY2QeIhfPJSlNuK0l86zK+xTnZz0FFAgnVb6mj4NFjmPB9DjLWhH
Zcxt0yR0a884/OKfkdVQv85T223gV0cSy/Cg22O0rmTbZ6HSN4D2JSBGzvwWoHzzmvLufZAVAiao
NoPjp38T53uUAK3ff+aGyNYZ4bdzT0euh+7bYNIfxd5i+23GIh60bcKRztnNF0j+3kFSHU9zEqTR
OUyWPK4MLWyzhUBw+MBZa0Muh4DwIj2dHFJNwJGeL1ZSn+nzOK+UIg9F4AjceqM/vnjYzk+0xcia
GwK49sP0jPjLEHjkpIS3MacEz5X4hIuBT0PGcNRlTjWnbaBimT4OUMvnyfw+/lFDWnF3u/oXZvNU
9hVGUn3dEZaB1MRxiSCLODR7hv4pg9lz/UNVbFNtmBOJ+g6+/RRm7uuBU0WRdzsXqK3G/CtVYuVg
C3k6jazH6XR5X4VaQv/5x9+DEwpe5sh1eJPfJvhxKavO1yZ+aOI6AMtnO/cq2W9yOvAFdhEiSrKp
kiEslTqdm1LF1+RbkYupo9478MieBs7xxzEo5Qy2L+gjEF1w/UtaXphV+e9wwid9U51W38huNbYy
auhKw9fRzLgS2vVI7GhfjDczzwFBAduXCqK44+v8cQjMhiZByxXnN2tlAiipqYBv+GF7meg3lSX3
DVfQP1M4q1NB8CWwB2sqi3oru/f8lZks1Lk4OIcS5svPJB2meKPNEOBYEeAUJcmmUZDklBbu1HXE
PglHUOJBYEvzLLVu+uuiS8tM52myPCJLrW/Dyr46XekdjOX8dja3Yn42og3LElzNY1TWimgEKA+y
ja0b5a+L8o/zzaEGV4NVgT1hbfmgr3h6/AwkZuc0jEjWDUFlyp1sjqo2XIIwWqI4EGkc8XzZZzsG
rEP7tYZHoCSrpgTe8tYsPLwhXES1gSwHv0CBvMJi/S/M/C5Ew2/n1KAZb0vB/tdHTkPO82ZV1Nhh
+x1gwip3p8ZuYB03SSRyr+hYApyf4V259bTWaGmy22bpqodkk6Qf/5UaJTohul+7izfuFDoeCsOv
1Zz25i//Yx5o+uZ7JTnQg6ZU9RSzct4txuE/VAq38ezJd2AUpWIcDAbF+45toOQSjnfblWeCKGbQ
dRhOnPFRI77iHe86FCXiuSjz7opzQCBeHfI/g+UmlaxwYqMm4qcg4UpH9K4CQrNX1pfrEQnJ8WrB
qhlOwMlMf1SJxsM6kl+OHawEhXL2xasEUWfs+5BPp1K2DFmKIIbjxF2ipnwcX5gKoMkqiydpAEyh
FED2clQB8fmi5wxwIfi8DqG6Kb3E3pGi/St66hBGoUtE47+IEC/qDxvaao3s7Hz2qXC/ak4wlgob
tNIX8a97s1N2KuRTJSizIYZQWlWyTHDLMMFhk2BRzkYtu0Z4wW9a5rVWnFqaScmCS4knY4+RKnYP
Xxa4qO8Xxa3dmMLlcTGGUY83rUkHTnJXPjFAGD4B7FQgLqKLPOYEMjl+PdFC112D863JIOr0pkhy
NkSQe56UsI2E0ALugMxLIrpMoukc6cpRoNMJlyHcHBZAmygUddjwX4ZZKzk3TpaZGKHuxMqtqE7d
0Ls3XlmmPzvVFiwPUI53GtQfJVBv3iKXoEoTqz2+z17gG9TsUJB+QVHqu1EJmdKVeKwm6FnCI2MM
opyvuRDo6zZpj2fnOl+VdgGWftv1go6NOvLE3xsWkkEOKZipgMFkZR5vAHMBaQ5zYOr++PiOFyY8
r+4jgxQ7aQMG5Yjweli8zVB4vy3UpS6dr55I0MnzYe+135wc0/p5EKKLODVsN6KF1/gWJXjQ60lP
hSkSP3LvEa/YYWo6NjsPD2dL+XoVI9SjfS7uBp8Hi5xMetB6sklCXmvFFN7ixBRSJEaMfB659c8N
9kCek72z6pDhCUl/JzHWFsMQ1YSuE+x0LpjC4tOSpiMkYNEGivF3WQ7vsfvuBfFQU6mT0mVYG1Bb
YbxAVKo/QNr89d1Ffj7u1F1bIzjzgvxR2/0Izejpy37vSdXtOzYHnJphO1PHVyX9H/M87HBLZB6A
BcavxyE9Z0dNsruzTD9k3t5F6tSlpz8UfDMDpIk3r0q/Mby0VmvkEMUhp1UCE4CJsccqSeB6kenL
M/BPHcdtZtFmoiqNybaY5KkucYk5fS6CZM1K7O/MNyD13M9QKgwZg8uQ8pixcsleAAxIUW2vUABw
fubPznZ7AjKvfc1nQnVgrEV021DxnCo+1RsHhcQxlMeK+okFlVbjaqPT+C8hgNpZ75U/X7KIQYrp
PvojOtRoEWZwtmphYc5qHuNMcocgQ2d+OzMkTRRznS4m0IHHjI04V+GC3KVqqXMFM8q2W88Lupjp
k/4pBTg08rM8clW0EsFGCtKxFMy/aciTXq03ZuIEjmnSajTVJLnbuf20VEe0iE0Z7FSkupDLUAj+
wM/WetdZAzE96I3RY44AC2ptvZEExSB69cWScDPfcYbrCQasHVqphofHdyjo5cExwkfkFWak9H2h
9MTrHjBqV/3Np4m04Mk7/oT1cJf3p4nqCtxrzKVheSiiPxnWV7QuS12hVQV395jWq07SkzABXizV
UeVuw4rsQoc7Yovi/+7Z65O0DJUzQRrO8gpFtO5KD6M+DLV3cs3BQh+vhaY/XRR7JISmN/XgMfAt
6PoqiiOy9uL53DzhcDKXoU/ZEWeMN0TTSBAPxfZZgW3f/hlM/MhA66XQdYw72xOlRtnDBG0rMYOC
c099D8GgsKzkEM5KVkB4wxmOgeRUlPn8yTg2gFF34Jl5r1H7QLKD1E8g6wedsnbnjVH+Ft5wXnJR
EJit/5LXZPgzyiPq7dDmmNG95mSwGpbYdsEQCPsDKztPuY3sgVdwSQ6AkXRH+Qf9pAVksjKYmyR7
QPs6n0Za0h2G9YkIfLzzhqSrSn8MYBix59wyxCDh8KCzU5yEtH+opTlVPgUOHqpd47gNHxYh9U/5
JIB8HtThzvydRMb1vb2q4WbuW3k75ShXtaVron4cj/2Njkw5FokNQ27iyJpwbWab1zryoSHX33pn
7/jyPiJkdaM7rStE+c+KAb1rDgzKK4Die+RGD6+bUe0tmjYJaFrvkoJaezMTP3YGOlb/PLF9FzIF
net1vTcvbI2RvNDQzzaOm3cAFvFJay6HwodvnhbKRWTkOp+5MIjKiGdyHogKCYrM/YigTqF+cAOc
3FI05ac9/OajD7uUC+UQf1FuQ27T0Orl2Yaw+6p1lzMyHK0XVVdrtMi6Ju2UaVYzBxgWHULP7CpO
lw1jH1M/HY34v2vLSP6vym6W/e5FjPnjWfjaygz8HTEzRlRoxiB7AEJOlJCgborueKqcTUNxBuDL
P10ZSRvUbhb1h8qyeHQ8JgUv8JvRL0GcKhuIS5MnWLyS0jFa9ebb2unj0Fh3B89IIQ4xBRayF+f5
lYoBwK7ajBslsKP7pnTwZ/J3J+FOBLQYJXggqHWjI+85n5tYfXzavigZEsi3I4UFeNXVuhNlwAIw
ag+bfv+jPiCLBsnOeVndgxc4S6iB28A8LXXHflxHAC0hWhGGBgLvvOYvHdlh/4FYowgV2MvJk+gS
J3XqxV9+fzofPolGzFzwKa6USWn3bskiENq9rpoW3aAm6x1UIAcw7JpXxBB4EUxYxCc4xhIHyMYp
i9inQ3VU5Dxi5AIXNe0aJENMlPE+S7O9USbmyYfz3uUDkTFvflI6L91izS4A+Jfi1Y1WkSFvEJpW
hG2v+9zRSPvFxrhJewEhQgZ5rWgIYLSxv7QRt9ezSjzv5sfaOLrZwCTO6wFFRdh5UWH90/saRO0Z
fo02/EMOEGmdKe/SjB9/oCowAsEg4NSThv/rOIXrwL4ze+rsZ3ElqyN5eyRESjPUY/KTeGUGs6bt
7TYSAFdjvQMJCzjv7dOBzcA3yk9FdyGd4OoSCbB+Jz1CBtDHJFXr5LwJ4GXRzEoCgqYy9Yn6XElO
3rD+j2zMEiC1exAziPVggrmK4aPUr4D24FUKkfxf0anvfjEKTg/as+xSQIsC96x/Qgx25AG7VcGu
/UHkmWDk8gmmIRsqGfRmmB1rVBDJkqCpG5cDwJdVVtEwZcmNQcwQtxLProfOB8l+ghliL+ik3TDq
uOd8m4++tPd+QhfsWcO8rYeIp8N+PL/x2FVwUMPEV5T9V0SvfVWr5Rl91Ynk3gg7+euYptO/x1WC
Jwtd6+6ZjnOrwyCcUL30R1BVCSRr6i3vDXgu4thjfO2SEMnC5NGu7EU+LAk+yPC1org72E9aXbL4
RWbzl8PuIRh+IbCIzblsfrVHWCpGw4tHTOROOvKrnIe8rx25GQUEm/HaTl8aZ5i0aWM0kV7pDQxd
fXL3bvO3tRg4Oo6KSUeh9SoUbJwlU4grR/6NI62+nmw7lhxfOhE+dD+guQ+MKdl8JjVhQMCFEFd/
W50wlSu/0Im7Evnynk2U6Bkk5ThMT/xwEk5/Z+50fOtGyFQvhLeH249bTavlVshyUMyiNn2Wi30h
1AkSkER9bpwkjCM/1ZTv85iV2gPW3VB8+Y0lJARdVnJnzh8vw60oEKHSIpiLS+czEq7ESMNs3mTb
iiHFpZ/wQhZ9leEvfwG7qObCg98SJWp+O4QEA/lcLfzpLOPL09L35MHxVmiAlXek0HDM60KtxMLj
9eBv+sSMt9fX5qlWqeNeywrTMNS+rE5bS5Am8lUYLzq6ii/FzCc4kZ9kZwqTl88BOHOMrmomgqY8
l4IRgEXn62x9JEzDNGntNAgSwVRQiWZ1P4KUOzxzfX6Fp10AwmhZu8gpB/FGEzcRnpMJitN5Y0LP
P71B3k6iaDyAJVsbiob3wSjUL2z282uPE27+3d39jpBWKBrhT9pBiIHYqW5qr0Pwy80b6lksme+i
bNkk8eAj5wnN53ilKGyDMPuIipCCQuAP+JrCMlneuQbUGpcLQAm64mNjTGKfMRGitTtgiZwv6nIi
1WJAiuiZb8PzXkBctSVEb07TBgwJfEXsvQJGblIh1QboLbJaNOVGMNXgB/45AF4UEsTUwiohRoGZ
xlsxiwlFd+CdhZHoB6ITpPzpazavlzkznbFCvyLYEp2SSAEAJFMETWs7opk4Vs279BCMC3eTwfqa
7zoD94Ybtj43i6KJglsZYKyHLZeFncOGemrD2ZOk9cSpDurIKJ56AllRQlfMHvHfG5QyrVBZ13cd
KBh0zvEiuorvHU8kXfnORow4WCWLKSLvsOMOoCaQZs6XnIBGbsX4oTXV+VW1duTspW4Xo6Jp5uVP
ci0bSpHS7RPtLE9fsKunOMQN7WKCY1aZ2yB7+ztmQHbPrDFGBeeLcHD95pCRIESBITinG5EVrNDs
cYdNpqy1YVF29yqDrZVt4elze+ZfV6+7mTM8CTcw+SG60bWx9QfQkB2Y6AXuQyirgLo8KWkZa8t7
1dYUyg147r9JhWlln7j2JNWwdT30YZ9Pv71wUKvkpuXL/RvraNLiYO9O73ZNAlk0yJnvZ7mOas0j
t+DL1eA87Z0QPyOUQmZU3B34kfLNVz13Va5GZFsO6b14Ms0KhiYsZEDW2bFAApLYn8WK0WWQrl7f
OHW8T7MSKS5gYunNwNZiuE1gvJ4qVwbAso717/sKZnrhpa3yyrmMLIgyidUIWI2/X+b7k1V7ERYr
1Fwde4H2MOvnRmNuYhAf5bQOh3tdtZ0goceQRpSXoQD0djM1956H4Qe5blIUGIra/R1glc43s6d0
4z7kJaNNkn5mextjT43m4GbDg5ZEINOhvBxpEaw5Z0OkXqdVrn9bJysdypcvJQwGte2z0EIFIbEw
7AWcnDpZtBFlP0gUuZ1sSypNyfmXLD45tWzkgAvy9TRzdeiyLYQh0GBBjHerSz9V3iNqTbvGAAnu
PrTQlAzZ7rcyP4fwU/Ee9nf4KVVELe4OlTQd/pe2AKfRSdOe51uVGy5er+QmXIGTH5cK/P4aPnuV
hUkuZvqpXOEtfEc3KCUgR3mpaziInit25pzXC4fE+/iNuJut3oThg9mxhC5LLZrxQ9Fin8T4ujJX
woz+uv4CSH+HT2zhm82I5rp/87ssXz3N4tBXyEEklscjxyXALuRL+EzfyiMBFA5uS8JnJV2wEBhA
dmuy7Uo81T8IYaop+6rxUGshvZSk09oN/9EsUmorwqmSJSIEC19xpp7tvfl7ZLhT7WXrsuep3jSZ
XoIqg0evR2TeGIC9c7bYSwG0/PfYX5trxIuXCN3sHBFDa0GFczezlm+Gx0qZvHQy47I+mRYhQaTe
C0L6qkP2sXvmAMeAg7RZAobPX+5AY4UHhBbsEL9uY1ZAq1+72BhHwK9KBxgC1tMqTq1NW56O0irb
kmXGqIzuTgrxT45kWdxyOh7r+hgoI0exAbkm3m7JIWDHiFGGDS5/IahrHQpBx9wNr+S2bR9WouEB
Oiq4XnX3KuoIK0kIT5cEe3u93CVJlDoYJ8NdppDq/Ng+tKebY0AWIzK1iKWGTxce3iBzkaWsvuVc
vH2sm8pjhURJvM/Gkg4J0sjX8FhTQK161Fltq5EwbLIkSHU1QRc2+DEksBD6FT0ROu7OKOJ9ErcD
VoUzIMlO0CCtTpOmEsUF4JxxOQuxjJ2UCYMQF1ETxZNWhf2ExMm5ZAH3XjG1ac9S0s4qlvkbik10
EUbtKvN2+DuvjCwXWgdXHi+bND8cc4gcLZRDjhuxBc55o0VaqaqpH0r55TUhN7IesOrVIW0BtgIO
DPfP/9fqvkIXvDB7w571yKeA75qrscog1rb0R0l6aotMj8osq8srL+Wctgu/8vlA1hpD+s3kRvCR
wxA/GOna0VO6WjBeaowGpB0el0el6vpDs/4QXW+wnDXSF9qDp02REOi4XyjyVdd3Dmr3BvY/b+vf
JJDJhJiShFLfGiRIRepSAeay3plhAKC26rN9bs5mK7XipHvLp6lvv4YXz7AlcLqfzRXdVglUiDJt
WubqkvZlxTtP1wgDd13RiSraPJwHO9v68RwEMWVJ6MMQEK1HX6L4Z1c1rEHYOZ8rP3lBeGColOMJ
3MfAzz6g1vZTPDaZYZW1nTMyRLl2vnLiKXOu9Yj2leyW9tSod6bD32iKE0pfkirqVXl9XAzV3QCF
QqNFQ6KS1qatHMzmIs/gIT7x7uFIGg3qaPyHK2k6d4zTmg6n8wbzAK/9eaoSGcfKr6eV22VaaF7M
yx1FAboVJu/7z2XsOf9rl6nbTjWTSObz56TgyU25vbps6RVDdnLMvr30UGiJPxv0Q96/tafztS5E
SJAbzdy2aj3AcNUNCuKdjwIoXthdwwa1RZP1rmsHckJ/w62mr5uZUz8rqTsjo2IXpVQGChbIaxWt
9tTmpWpBdi7+SAE8XjiO2v+mnZ9ehb3dk9vzUY5DB7E9rEOulWbipKU0vEibUxrNGY/8fApRb9zy
HGpZoR8WwG1uOxWBsrBr3SytfgLTyBHf45thV7IBQHUsIfGaYIyp/HMGl0lDtOdIEoaqyd9lsN9F
A0O2lFzAfQtBipUlVOBp/SHBcV7boruhgt7xxOxvPOnzhgvZdySx/9+9IPNioYunsD1HZIShaYI6
eU3bFSt1VquiDmWMrWW5AZAfR1fLe8r8fEhg6ZN1AcqXVOS0pfRG3jZrD9oBKic5rARFjCQTvq+1
JIox/+viHVTihFB3KJ8CWzXzC/ZoMluR0ZG+2WnKyX5gR6221M3K6cWbGOJBo3Olr7YdfRKS/QK+
UJCxQIAP9T+CgJRfrzAgSKNpuRNQej1TVm7WA2CNwc2YlJgG9SJNm3p7XLGyB3T6tihw8vJZ5uhT
+gG+XOTawBF66z9oSvOXxNcVh+lUtrrfYPy7jpIgryYOfueHfLdcfvr893nbZtKtoZPLr2PvbTUz
zA2VZldgySfrpgHt5QlP1VWkreG690+e/In9DYwmI+H/COaMxanydIVvnwlHvlgoQ/R+k0RuyB4h
OhGcak4U5KdGqHnYdH6ROkc9PR3vINGyNvOrIQhN/GiCuNBgGUYdO0c+Owoi1qf1x2/SvqoVnqFN
j/nYKuHvuh6ll9bAe1dOMHMAKkIWcFR4NNjTJgxeC/aWj09uORqERYWCibC5md8zaAY8c36K8pPU
ZLJBwHUdZaXWnxfbfkm8FeYM7VxRoSY2IB//bOGYRl2ujISSZB9i/DeYHXQc3ahsXypSGAg/sig6
+mJtJw0K7jgdehI4ix54mqShr1ljxpZXlNyKSeNRuOw4mdZOpsv0G3T9+zySBE/WWBwKtfGH3DRC
rW0ouo1W0to4tAQBcj3EthOfUQDZnRz69eRrp+shgKRs1v0u390xpmDTjP6vF7VniY06WCwshpsN
esRbKVUMeCFR00dzvBTxTK5MMiEotxtzUWeSBTjSc6Es8pOUvZ4GzKPyTyLN1ZBTmVlJRegBbL6T
r8I5zsEtIJElcLgOwTELIqn1ciVs9ZwHO+9AZBrhYBguoihQAp9riD3hXfZ1rBj4ly0sIooqs9rj
MZXrHwvJXpM3yadCwe0eAvMdqIZUJamr/U+cuevDnYChs3GnnyG7fIPKcAWRAY0Ru8fDiBhSqbUW
bzF9B13Q+jywH4jHbZKX/9fQneaJ8hN4GXZjWp1qACRnKvHzqeZOV9rfpBpXNKC8538u+tL31eEr
f798yzMWh9snwKgdFjEFKfkQJ4Gu9B0To+8/N9XKFz1jH1IlbhrUI0rW1T1H0fT84VYl2A2O+346
XY33T17CRmeT+BVQ8C6b9IQRFjJbqZ3YvI7XjkAzdnjJw7EmjuhuriDcGR/0xy+9XsAG99q9lD75
00wFzo2JRO81JP3pvpEg/523wxQEoqZFLYoUkkbRaaB7izxwlO2Ng+9gj0puXq9pU03pG/Qb1v9n
Yr1IyW4bNfSuGizFBT0MVDwZUgFQjnsBtRhbiZxnb9NqeXGXCXJIAnO6wAoyCXYKpHZ1FV6Eb8+B
wZUz4ocZQHPABAi9XXpzfDQewIErJtzRdUq13tYaS0H3ao9SHal+wwxVc1tYMxjgzjciBOPfo+vX
XJCz4QZ3brvcutsHkP6O8llZPwtfl/osPWKO0HRsL1zACf3QCcYyZNDLpUCIdBuw3pEwjovFKjDC
Hk0npRrhUIAp0OGtEyV1VOOQlDijSZrJtTHHLOto+4/Qsr5iTULQ7WBFOxCX/zrxVj6E92eu2Q6J
gJvGKAi8XOYp/LYgRYYbMQVpgVEeCbBo+t4/ZekAAtJqPEb00ghOU0qEWv1rKJZEe9tcSSaC5DE3
p9HSg1BlP7RWS1gElmy7eNp3rWj+YJhC4VvyxF6ITL/VLL0ldPdp9Cll7GPW11HQ3VRS5x2K0yHy
hfJASv2//2B/f4PW/eMSyHLWDfw1+viEak7sXfLldDysXcFGnSESCaKRyDV/y255Gca2cOQb5C5/
JH21X1Yowj9djnLhRCelNc6g9mFsZ8X2Dn0RnbBhZC3WUMpa2XZ0lD3fKBfhLBAg6eDISvonBy/I
RCM0ov1o9nx7sD96LsJXELVDFs9kdJF8Pn/Z6VXy5KYCMA8hPow1SWcsv083OlJqk2fJ2e1P4vyx
LerOAcUtSs9YwsNSpAQrbO1oyzG/18mOl8+PNTYffLeRb3rcuX4ENsiahlZBa8AreRd4bx58gHdi
Biu1e/3JTevphA+dKIUjeC3zdxwFwfAGSEX+24bDV7iWxN2ZRFHPjwnpzcgmJyOoN3kfR6TSHVI0
FhOiGbYumE43IcobceUF8QbhMS13MZbFGF9NqPNOh9kQvpzxE3Hw1XU2PpraL+etSQJXHyJGfpPn
0Uz3gpuBOpXzvOYj6VhVh2yz/3YTCMUggInajwqZ/0PydJkhI2HtH05Bs7Wkp1KTnIRbjcjh3/+S
FbohJ7g9rrUTKKo8Kj7XljAUn4mv1VBXhbze1vT08Xh/UeP8sFTmvGF9L3rvWJ2AyyJkOOdf2Kxd
nqBunLubU/+XiLWNqUfh0X9p6503WCSU2mgUUacDLArFrZSLdn+LDJgjCa3/qi8R+C+naDx2pCYL
coD8vywEwEGMSBnuNy75DFYXPlwAlUisZZoTu8iTvbQb8sI58xlGS6vH+piTGid6OdDDNQyBmN2W
IB4/UoKEyJ4RgBZLlq0wVmG+VBVRswl/JF+9CARzar21iDTI9WkmaQq0XW9bWqWQCFkLrtUptevU
XRM4c4lCar+sIpiYDVaJiPbhdUHsF85TjjQWpRZZijD+BfOT8cuKL+PrT8wYzWv/OBlYYTYT9ZeR
GaPiaMnL3dj7zXiDncBeJXe4BmFudifSNZuNneA6nBjCMS8PKTfixa/uMomAQK8KTM4BG2Q+f1TH
Eg5KS2IxlnHmuLEvEfxXLEJ+qHs2ToLG7yCfm7hVZ+0P87wfCP5kpyz+mXqivcvmC82NBJLKYMOJ
Xq2Fbjn7ivckgomZ62sy2ZJfxzKzmi9t1/6xhmK2SXUnga0axb9SwGFL5Wp36OTU2lSPTJHkWbwL
jHy2AlcfNWmohELa92wcJ7/UNHxt17v/6tBJDIRa2RLX+cKEkLR0yXNRq+cyWhP3GorDk6GxzBf4
bfpQfOoatt/cgBdZ9f6GLhdzMpiWwdvSkgv7MFcTWC+XDVVV/cyp/9TkrmOhQfcYrBJ9tpAO14vs
vsMVaS13DF+Kjs5KIbrYVyLgXKJpuDWbGXpy3nWoXiQo1vUW5BoXl8AeXnT0+CuHjuehlSvP77Ly
GI2q+AQQ/kzyG8wWFiwDzQYzHa3ZSA2rHNzHBgPVeigML4zR77eyaoE3MQeA4hK2Fq4We6A8x8L5
SSHkysG50jS02tcx+BYRXg4VadWSZVDGLznCROz8UDtvMfBocSKDhzl+bFHRefeR7zcryinmZ+K2
BY9/x9nQqqjh6jqtiyOYtcCWcfCiFi9ICQKRNOhMXMXp/oeJIRBmjonee6EgRu/oWKKm8gvqCCvH
DR9Oe0gfP2aXkysdCgX3CA9su0Qgpw6KqpGRExErw6jcf526wEb2zUze+5LYKTYwwqYmVSolrQjO
nD+7wBBQ9kthRL4FqfxiMcODZvuH3HcemSJ2sp/YWkDKPdQGTcP94BboGjWjgxdO4wYm4LmHrUXV
bHFnJTFf/f1WrHMk+gtEaJDH3l675PT3HKSV3OBmSt1O7NimGDfUExsdURjEh30R3LQotyHRyJGh
v9syw0hNoUd8f6cKaxNio8fCl8JfdRIIm7e0eWkIbwJvqTJicnC0ctCFpgn6X3q2cM/ioljAZldp
GRKjewIWsSltbL055qEeWiR40HEJrY9384OrkBcuqkRZ6rdYlubaChQaQv1FEaTMIT4QKukm2YNP
UdX4e6Oo4zhByDOX5L/NTWfphxv2xq3v+gm9DLb7CvGdRTCpQP+dmETyEG80zJMfwb7Pmek3ByBd
MqfoSglugEEc51Cc0K2fzASBFKel9OTyGzjQfeGRoGGL2XrwNr5JBdPCPAfnkX8YiIHYrVP52f3w
D6hiotaa2u2/UUaJ7Gi/zh2rXudZUmQYMtbMoEZgUqJDkxCxwlfvQQXkDY7MnLuR0yNt8IIZl5aC
TLLOIJZ/8XhCwMvj8dcjA3W29xYr24o5ZRxDnpjrAsVnu10/pvvwWUoDwUkzr4hzu7P0JPLJ8+VX
wyP5riAJ/8+UAWAPNwjKu9WgVCa7sTjrI6k1Ou67SPZEo8Kp9Adp7f7nqym1/Dj40HWekfS0tnJj
UaGhJSze+jbZb9ZzgwAZ5mzenJ49fqXUtkQ6yY/YXYafrkOGfOGPVRnBx8vGdJjCSuyfW6Bg8vf0
rKI67jxsi150b8IzVv6wI3wfaEMVeqgdpHRZPPJjC0AR0YbIpA/sqDt++1Phd/3tamll4uDODfcd
LOevQQHLQO35c2sHavhLevIfHRmZSvEbFjvjSW5yKpHbSCGpMt8Ryzk7Xczn6mM1cjXmY652QeAX
tkFLaA2lT3yPmIYwPyO9Wt5HArwYnW2VpJM4LT/C//z1H6jQs1fp+hTa8W5OX/Lx60QWCADfoHhN
EaCCQHqZZZO9WiP63f8mFoCCmKTce6rS5yxcARHmZQpX8BShCG67c+lKjHQgYGOHoubJITwqjPq1
Jpc4Go4UmsUqoS9525Fik4SNulaKb4YghYUd0Xn+BBQdWAh21hacmVTIiI/i6yFAkc63yCjtEXe7
SJyXTySP09/a2OoTTRL3pIFwisJ5BZWK0XfYmZSFBT/dnpHMEjZTgnVQyljHNNc0eoDvfW7qZBuk
byGeNl2y7fzTEclh1fXoakH+5GVW7oorwVVZ79zkxGWHuXaBsaqH48DnHpArwxw9P8CZkcIrUPQm
35fgECd08QJTwh7YZUCxfIfT/Oj/g2horsiToD8gqCAKn2VwAMzbWMiWixcQ497talrfCc3MXJNY
YePpaYJVlVNkACJOPswgrxy0F13BdNF3UFQlGeJQD/eGEBOrmSH0I1DkC5CPHU/VcfKTOa0BS0Sx
FfnWe5WJebobQZIcAUsxsjyzxJGsENzeC9LV1QN8pq31kaURcqjVJXzsmgYms6jwClE52JPWC8z7
x4FV8WARSw5aIswV2IknuwMuiuJ4rJmDu+0hQ+oNAxXX8NzJex4htXSV9UFfVCeaq9HYmXYMU7K4
f/UDQRoL6imtEVXG2ucIg0h/fXPbGahEnTNnxH5UvDmOAtU295CuQDXom95CXSAK7iJLfwVSrp38
tLlEQ6sgkvZjknvCqILzb7OSmn3Vc4BKpf3ZWnw1HVt5TbCNsVvSYlGAdJ7KxiLaf4aqHj5ZKNI/
AksX4AskBqQFoN/SsTax0Oc/U1T9FxCTos1YhqMnESy+la+RdTfa3VeUVl5h7PNHuux3iP+Upv21
wba6dJFNFsWS2seWh7K/NlBiQaM1QNVfgLjm8bKxGO0LXEXz71KT3XjE5c9eb1LVy74PfNRIoPEv
UgxH6LUsgdnTCXCr/eDuOOzklYjfNLC2TKBgXvyKZrQCuIWmJjLwo0QlX+s9D1oo8xSQ0wU/dHt4
uENB8tY6v/H5npCoTjYVR7JYgWbljk1FostkzTUrfcPhxSup82Yx1+kjZjR1/8qKj/OXKcw75eZ4
oMKJJEGo/scdQsFBb5IWZAwEPfTkQvEvYYiUOWzLYGbDWslwqX9Q3+Zbn261PLezN/EqoidG2P/X
lA1WbNRRiRniGgx19AiaayLjaQDnI9cXyAD4lM/JL1U6gtp2UkuCiv4SFXlKm348cF+Ii+8Q/bTA
2DjFmlp94sLTBtLTVsLCb0RTABnvuE5CYkxGV2ZZL+7mRoinJvNR5Yf1KEMu6O77gY2YBFGcqSSR
/s4StCoCuPZmuf3kWC3UdEQTf4kGgeacRc0a/uAnQq3LrlwSCO37ilcfihySnKcV5fRQpVE2X+yd
I4tpJBUctVPL4q5JV5rLA9vbZWL2EjRM70qqF8kJuzfKZW/9cF32RCtiV0YLkw6xFbNMberDDzqt
nMIEaNyn2D1wI7y2P95xpe+579x69pNMHSP750Q8aYi0TDLDnfw7d7FSguME+JYMKV27HAvcAs71
GHrggGzYLTRyxUPC3M+IAuAazXiW7oHn9M8YNRTEmdy7Te0wfcwj39CjH3U2mn6KAyQ28oXWy34w
9OnxIRhkBKpXR3z+iBZkZGm8ji3fXY7MUHOO70kDAWziYA1FS8aSJFfIMjAEKLmTwYC+x9jLXsbG
2znIioGWH3rx9vdpcOzHpE+f7EaWp5z6BPBZCwzfZPhN79wPrYZbPIFdfR8zKqkeGk0uo/7dRtyb
AUXqUzOBQ0BknI2QwYQ+0m+zY8QoN38opj4760awKpwWDirsZhSTFGzBXN0uS1OG+xcFAr42NkKB
+Nu6b4JT081qI6EmJ+lU51zW76Xcf/S31A5sPrKpbSPuyZFWCz2LoG7J2JnS9q4zd5NvCPvOj7Km
XultMcAqLvdEx4gIr93Poc7wgVF4LXy8pFml3v3GYF0UVv9D8zPXIpuEbpXlMXBlE5mCD/uW3NBg
Ny72WX6CW0P0quMYBVdNovdL8dkXbc7eHgLJ6uTdyGqAKXCYHvjJ/TCl6C+fKfVZ3socX1gufWZb
gQpvupMB3afPDmFRgR6jnsQ11y8JMdhUxLLbP5fvnqM0v+LRwSICD7UL77KyKWnmnmQQRboJGVbj
JHV62z7u9pRvPgJC8/uQF1F8ykU0Z5N1j18S5Mgj/s3Im2lQC9mPk/KyF1798mNpiGXwYjAPrEou
nQ4XxBSSaWhLjFjG+NSUhlkqeU2+mz8OVWG6Jv2zRbDnpBxzEoRa7iFmoJBPO3IBYbZ37kYoUiJV
IsK2iw3eTnWTEBxjxBX14vbGUdGAOaMKBk/516+I+/STV9g3r3qS9tGFmIlCRWR4leEUKuxVKC25
aacZYqXuAVolc/dc5pJuGvoSIXtWzsIShQAB4+CIdiMEzyYZgrDthf0U52zkPEaOESLb8UwY3hsB
q1E4sPazfXHWryxsMZ8z0QKSz7Rbwr8QBMHF+osMgyUyqJAbYVP9HmBtm4OhiVCgiL0d+anOX5Oa
CaV577j8ejbF2MrLEb+DlSNd4Sp74SAvutFCU+dNXR2gVplPzaoFiuQa7yxeUxMARKglrp9qSbPQ
y5UroaWa0tFQoUwNSN0YRqB345YgLFu4naY6k7Va57EPbyw9Msn3cqQl/aI9y4aZsmsXhKZD1w1l
6SahyMroHNBA9skR5MNHi5Pan742Y9FBfBrbNuz48ekLCoJMmNGuDGlX5xboc9iCokkixOa3GbBa
BLdYJMYHaRLAzqZV4hg5iUJqrP29OeME7KVsvTcM/RxE7Er07ODKNc6ijG1uab9FFPZamD6pqfjr
zV1IPCSLWxc0KUDX4ixDaCFuowFKp2JqogJhBawYjWeZ67/toqAF8TUL3GI6UuzandyTD0W7ksJ4
kbd9AfQYIGAZVJjVPUmdVa+MxLPVLaz9WQuz9/G23fpemCtKZ2YdqYVuCEOhl83CP+OYyKpnpDwW
YWmswgOgieUVKE/fXquCXZvrqxJr4HTgCFJk7yg08srpl/XX9L2t2K3stN8bNdRU15ilDBdm8pRv
r1hG37Gd1AlWalXTHVuRE0KH7PSaRsOLYyr3r19WGnnwazhoZ5yKEs51ws28AAEsQAy8tlSIJ8ws
kiUdsBi8tVaO+KLbgB7O+PicOq9ACVkETALC/dSTALagoodtdEVJHV7NeStf6zeFY2UTOGkuuYqX
7FPFL1epv/m84x1qFdE3vwgJD+U8NyrfIJLZvavaZ0UBRHBAmC+SNM0b86ps0KZn+Cl6hE8oyUxD
ikk6UAW9fDcyRlw/tAijGnNEXKt8H9WfzrGt7y9yXIBf5O3c2VT1caF0r7AT2Vd77j0xmA1r7xoL
IZ7DTovb5ajL9e/5CSb2NwrUhO7GumURimA53fm7JWn8SuSqwZ5jieG71SXdE7BpY/xhBbrwUpDu
Jx0u8FBGg6uw6U8s/LAdsoRnjSFCMHuvXYTj5MyZ1LebQ3ozuxW8O1dIZMYKrB8gZmEgsC99nZ8Y
4QG6XnTnmVeZEGkkQVSukrJNn9sRB31wtNs17Eyd8jiAUuqCNBKuw1qwAYKee0og2+08NkX41VmK
/FJgvuh3u4E7ymkHZx+DY9XHbbcxlYqk3J1KnYwIVvndSVFs2VGEVsVx43hPQaK0UfL1ZqCc6eox
Pa+69rBqq+PhOA2ICCvQ4GadsX1zmdHuEOEQBdHObDW8Gri3vkl2fJAJRuY0haxTjlNiWtKzdv7k
hJ0loj/BjracABbu40TLI8zLUcjWMNg9UiUn+3Kxz6MmCQgClbf8dz8R9WzqyNby3VJdtw3smxyo
5egOaIUF30edTnhVXk1v3n+lRN2YSmz5mnFyTSGUxBTTm/HIeizV/R68p/yMM/jSiwDVkitURUVX
d4tXnwRxveQeQeVWOD8dwPemxEjmFdidQgU45AO9DMDp1FhDUJVQfN0/7dNYjl/WeWIHGkAGiRgO
XHqgkf+qNdmL4rV24ptko6C3ZpNRSG8T32cUL8g9bKuEHkJmStic+bS0G4lLZJc8k6k52osQ/oql
O8fDvMB5MghZl+XVP1wqyvYkZ/1uoC65LU0k2JUHGF5Lo653IKP5hT5bY8p4MafaA9J2W8XVJST2
5TcVbRbtpUEBbrcoKFjrfmDvVrvXnkVMy6/+gvnpuiBmM+La/IjVtAYA5qgJiE7YCJlNJ4kc8ZT+
FRimCmpbLXZWOZ+Vb+fz6JI9P7RJ8oVu8YnFPDmNs0HgSaKH8F4i6C+tmiyZEuwsblNiId2S0eJl
WNvjZY1nxX2SRjCkQroo8kRoHuBcSxR+FQCDWTJjOcc1VABb/63b/0owpoQtwKoVjVCWz3nCW3fs
JKgifnT0OQHjD/jM3TgDEqr3DWw+X041N+KcfBQ2Y2FsQvnYuTpWqB1dvtY6rjldfmVCfRD9vA6y
wfspVcbtoQszToUSsBjvmj6o685ajGErqy9P1PSOJT/WHajacnSyO6jmDLi+UzB2jzC93dov0fDH
hCoEAWL3KrJ09O5p6hm2MdUxTzmrKofWvR0/Pd7y+yC5zWFra3sj35lFSHKA3BgQ9CUsaFadpugF
uTEKxLI+gN0TWIwafceiEvrhS+fr4SKWHHzROcszFVnrpibW6kj0rE7in0J+6ne9ml/Y6xuboFxi
PuqcBKt6EBG/DaE2mxLojVrOP32UQ/cGrO3+EGg48HdkzHJVGReDL331Em8XetZUyNpuEMTUCr2P
QdPXa06KrHOqWKAYjD7X8aFarx0nuYQ0vFywwvPh7NZSCCJBhRryDRhbX3lr/pNt1aSUY3SDXm8Q
pRNzR/3ZvINHstzjqrrcPwG6awEclKTaF9hjs0K9iYUJVbrza1tpB2un4wT145LNXV8SF5vAGZht
FCmx4nlAClu+IDoQxMJiT9FdS0zRsMP5dTD68Cs48RBMYoNMOz0I6fQW8cK6kKQT9qPXNiVod14x
8zskL/JSO63lCY/Xzh3Kfe0KjfOCSQOAV1sbtHgHdFKw8NkGUtZfZ32b47WarKmTIpkZsgap8wWU
BM03G45Fzb/WxoxmHUa7IfdBndnuUjWfYe2e10Ny55w2CTUBScREgCIDVovUW8JF0q4pNbmQid8+
d9D3zypl+UmgxxzdnxIV5K0Rla4RFa2Gcjr4vWk5247NFqUXNHnRoacFgBWw1pDLlEmAwoy0dR2d
LyvCSlZOXcBDeLHiixC/Bv0MegEmvgCflU0o/jPZvNqcC1KbTysZs2K7WP+XOFkWuLlJM//RRiYR
+h0XfRqSgtdlDWuzCEjl3/H/ZRAemZddGQfgbBV0pBJopsBvQj0C7906Nc3+bM03dDUAgrFDKSZH
+Z6rXscrPB0S4LJ7TOB0KfIcyu4K7FCkzuaWFxTTC9vVV8qD4aV2oGE7w1Utug3W/yC61PEm8DE4
mrkLnTtRTERsKhD/4if+7PN60C9Ij3mw4YWW0l+87/dRk8tihQh27a2EUM7rl4vtkv4AJxsT9bTu
shioPrTR93CMjTeIHmRQ3enFhBILpdX6RqxchZUbvfAnmEr+aOyqEbr6mwBBcR+5OZWhHQfAFBEm
OmU8pi4yMiWF/BtAMlzRDB1O2V492utjGT5hMgJaM6SgTJhmI2LhfSHVHV1d1/BZarkF+WU9ZzdT
5bTLRKNYG4+ghd6K57pHcAIJfFoD3D8Fhy4ZMfLLSDCKw1gPnjWTua9icOhOBxXYLZUKuJ22XfJu
UfoXulYFFvEE47aAwNlJAJ/+680PdOnQxALu/eUz+dvvB+e1KK4a+Gat9PaMTpAeEuz7bVhYN9Kl
005Nh8nFsr0Lc1wMA14w/5iDWSuceW9LvAIp98EjSy0bUyLG8xQvhMYj7Q5E7lww8CTB18W6yogr
h7mMQ3Cl61xVkI9041sxfhXweaN+Tuy19n/T24TUEkazYW358axb0P3ifUSJCggbwKCcSpCXxi6M
T+tUSQQg71+Yol2dKQG42zEuV1xGbot7X1rnoRtTSNEoUnkLh5WgR1tPi5CxadltHsGclIICFTf/
9sAxVyc63gR+SmcubF433h+kmRCWGJ37xLkFUspgaA3fggEX84lfXL5JeTjOMa0PcK6oFS7ivKae
R6BT2mOpFTzU0qY/77oGLtmfjtkU0cNfO+8KpwRqsN3z9AWIDdjPqj2ZWsh5Va+OknOas/u5v/Ph
fHZTPCwYzl0ggqb/aOjQtXuiC4G0rGX3oVjNVBoNZU9KFevwwuPcf1F+Df6SmEcmUTG8n8PJYplG
EyG1ci1SCknhhvhm4Gim4EchOZt8CKp5Pe88794345U76lVFc5EhlhH7w6IBQv37Z3b7yBa4qJj/
FTMBaxDXGT+Vv2vtaChE6y7JWgWbXRrHyRj5Y3vzTTgsgBWmMlMcInqYnBPtOIwTbCPKkNAlfCx9
Mt2SXwWSe4eXHaQ2OGWcJNXG7VP0r5Tvoc29ILtfs8kaXz+JbH62JfnSriSj0FcgkdXm3u8O9/DL
tCLQk7vMl+nWrFBZBPwf3GhMnGnvdec9KYLQD40IkNWRQTbKSd9lT2fIk4H4KvecEjiubS5E7T3c
tUegC4DsrytZL88PjkG1AFmthPYCfjaU782y/xeHEn4UYcDNtWV2XZhNKnTeMP0YCMtKp+vKVf5S
HkQ5tGdXTFxtKtkQKeYFWdusWcABMANn3coC3jD5DfQA9+SVab98HXWBsOsX5Q/tIW8AVRstKHoM
VXe2IYABNoP/o2nRkhdFmdIXC3CclFQUC4SsWqvNnk6efEUC52pbxVOcEWm+s08kmDJcOO6PYeat
2H8uP/5ST4oeBh7dhWQNEsu10NkbNY7sKdyogGcLDcnbriR2UklprZfYoQ/LxF0meFKnb7IImWFN
tSeUlnvSWkaCiUqqAoLTRd/8WHIyD9g/cT/zFyoNWijV2C/g9EmdAoanjpEP4AIk94lYxYlVeAFd
7R9rJRoh/vKOtwXBjVBOvSFKb/yghnOlwEOKG7mll73suMKaDprxgyuDLlxcu3Ej60DGsbI5b6+3
58BLddBcrEZio7cVg9BDw5Enq29NknC1lqGpoq6bqpdqa3XbvafkeH66U58rutRxxeXvpMGNcZJT
N/3usLMFJKtc52ZfLFy/C49uAycmGmIdHi5MSF9k5M/0eJ9XEtZl8vMLymPyE8jatMbGgLe8KWX0
blLJskr9gseiRjSBBaInAeM8aMfOdodR8CYPDgwvRZMIlXAaFg/prlLdHalkeUkV4NxtdiUaThzw
PdALVf40bnkkysOfFALLfveIqck7qcKCRfzgQi0g02NnfsWpSTIr8E75itd+y9yLi5Nv+Y2JnMH0
EKvteQxvQmyn5wjVCaK6S9vfGjWaeDcVJ0xmr+3yvwCcIrb+NIn0DNipy/qFltESY3gv8bQeECPB
3krA5J+4ezjLBzshlCU/zHnznI/PRk8nAMOtVxpKJbwFgv8V68GDFmuE3KKoFwlD7RmuTBewMDII
uU4ByZM/zwJrB7MbD6ZN6bmufVA9UDPuXik48BqfMPNbDpw26nSPtDavPU+HfqFEqMQGo1+ayjA0
365X4HKlQtpq/+YSMaGF8A7NFaMGDr3cnPPSzTMsF0ke/D8mjd9Nd1NEIGqDFMzmsSdYAmi9vcBS
fN8jz4ONPDyFsEryTed45b6oZDdCQLyl1rHFjQelHzILsnKdyl7wL37D35l0i5DPHuEw7Y6AMDRC
C/8o9yGJ0kJzk7Kd0kXtjOYnGLpKYeUpw/eLHwMngcUhhYadpu3yE4EC/047sj9B7mepy2f7+HAG
AijFG8kg+I/BmL8NkBxbws4qaIGoYw5nR9JDHnxobeYQzthNgwqnElLwN1MkouJFzDfu2xWzT1PX
j4Kf0FKMnTe5AcZe8COiT9BiG9UcFxTBpCGWcPx74pX4krrRMCUTaNJ3KRa/pGfXTw/KebZR9g0Q
eXdHYh0SUkzG7h1ROmtuvXh1zeDGKT3WlUvOIt7E2VJwPmsGxaxZKCCsna8uYpKID1TOnuL0W7b+
ClcixcsLd2R6vRqo/nXkDnSlZfJ48zqInvFsmksXIsYKIh/ldq/bTSnktadLAKJL0CE0adi0DzbU
zKrzDJ8D6rgJgeUIoDTyrOCQevpgRJMcCbhTaX/t8t2P5K6K3qHOG/mZ6bFHo4uB/E7lvmUW1TIT
n4guJ38o6KRVJIK9X5QJxGMJI8Tn3JIM5IWam4RlGMk+GumEGlbAtSeLw06TEKVI1LwoF9AJ+oc3
aSwKWQ4AIfSMBDqnbljIVIT5UypIq0gh+Glsj0Ae0mK7ydl/wPBTQRAP/NVWQK6QB4uvwvE6AvH9
7s0c1TlEANIlVDTddkNGuTFAq7n81VE0zfzftadVZHwC49TEoU9QZjZs85R5NHqKJTH5HZuqQrdM
1bmg5WYEXlsIgJTFV3vr5uDX5MeYm4MgIJNlKbiUumHQINOVftfZXyngCUQz5TG/YiOjOsjHAUhs
KBmx8JJC5vQChOvA0eq5EvXQzsGfFif7s7MUkNfNvDyX31m+tnFJTHnDWKwHMvzubsKDxRBRIpjE
n8CPV1VNHRU7/GrsQG2zx/BF7HbRqJ5f3ClCE14q/nG9sGCPR5QKlq86jwsqFLvI/HYilbIpVGrJ
wz5UoKocjuzqwBXYrPTcmLDJdPMs/cjRuMXBMzhjMb1l1hD84xl1vTQuZYLU5gsRENQLxBq5SQno
aUIBmpRQe4Q2bUZFbz+Y1g+7dfPZMi/QnnaleGOcb5dvVXHG1T/Oiq2jmULnByJpRwyBncDk+Yqy
i3HXN1F/IxzgjtQPjMPwLtQ3sMhL3JIPxfYdj26vBM08wbSQEfa5cTb3jA9a9qERkUFBnJ4mTuar
tIDnq8WOS8vliewfWAV3ReNlmq4g2mQPaTTdTx9ZQx2QTsFYplvfPK0EJ26PtChXT7ZwoMxNB0vz
dl09X/qAnqBvPDth/4EqBbl4ch6Y9wfvfdwCDu9v6ZtYzMegnPViXRFDryQvKBR/aHpj6NJ2phjm
JN7keCG71hdi0VhDqMV71CqdbCcyXqkN4x9uSTAxr0RvD8gOwkqaRjbK3SZZ5lNcvl0heU9fWUmA
Dy8zRi59QEw7ufzNkkLTNL4E+bg1Brp+NOGjRyj2EFO0kl+pitgiD3h5muIHVPvku6nzCnf7uhwq
F/c9SqThVa4d9t5plz6nyIKB6rVm3cce5ZTYFQ4mdTP0txoWoRulQSqPRxvLpaNAfJ/iC3EBE4NC
Y3mCOAJ6qwMdxYccQBQwHvm3wgEq6s0kTZTDPkZw48bH2PpKpbeEFh4t4qGhLJluNeeo62RJCX7E
c+/R7qA6h+8xoIobxJdPEqAjJDZiD9977snAbheZuuc48lMVQwj6sneocVkFQISvVTy6hldRx2+A
CVumWiX9ZJJQTjvbAExPiYL7CLkbu0c4QRocZTjsxlvEoIjV3HG9/H/l2XnJTlxnLRPPe4Oyw3Mp
tvHUBf9rW3C9e7rUYoghIvm0dKOalf1FV36MCSYp9oWBPHwkAv2w3cVl4p/mXRWbgn5XxPuk25Hw
XB3Zig4SbYyhO74TNW8KCGtPfUcneUkw4g6wHb7Tt2RtE6ahIG5N9Y0wTgM8rOQ7vZDcArwjD7IZ
fK6YshhbLd5S/XzXwd8l65Htyo9Ch5dvvYFH9q4jY408QxeWBh8YqfOF5MmRydYfilO5uG023unb
lgcKG6MnP+5X3ztDxpNxZYVvkQjk/+8LEtR7WaC8cIXgK772kythC+EJ4azcUvi0XvPk7ME2O4yg
hA+anzdvjKdHr87/YJKOt7KLJTbf7BDXf3/6pP59GPx64e2zZChpQcLKaU3E3E7+rILCcct1PDkn
jn+gcbYU88zvJepr1oED1KSUBTH0aRAfv+0xaCVrPFFhNVnoD8XTIr7JkI8/jwAPxikmoBqURiy5
g1k5jXaLvlW/Gjy8cW71hIHCwcr9dmZxN01iTEDdyeDcxf+5MfMFhozth6GCak1ogUUd+XLDk3HQ
ETPLTV4ucFFyccU6nvO2zn7QGkGMVkUfjlmY0Q4jz20eJbByG2ipJ83TMTZAYpxqq8LOUsPnJ2Ze
/bioEyDV6XqhTpt1xHKRtIfEiZ/0diX39etN0VpWKUkfAWKfrGFnzL1KpFfZuq+EJqLDRP2t+0ZE
9GfA4rOxjOYhBt5ULku1aD8itclskLiXvSPj4mt/O4tamiM1pCdAi+rANeMjfoPW1PyF1x4b418g
FAG7H5bI+Yz8GzlIJgiDzdzXOXUtdO2e10r8358dRXAclfiszDFb8FtV3tYsK9mY8zRZa+ANKJs0
8vj9htev6JtKSYMK11WOgFKHNchz0DbXhKq5ib1EYoeopScYS+ISoyqroshD1Yz1E2oX7u1QYrTF
qaVJ/bfjh2S+olxEV/WmsOnmziVuPUPkVv7SIDG3dmPXXXUn8eIVdbuacF3CDTgA39g3z5MsQXqW
AK2AJ6b1x4Pf+FzwRg5qb/5ZWbHwwYoCHQ+cyfxlDBlYSEIwFIhSq1ssr9tycEsHpa+CfVi/Mp0O
nsOUE0liMja6AzzSt7UP+CzG9eNvpxt/saUozQ8hCFHdUEwn4QFeh5OTb3eBys+jh2psfV2PU8QM
LgMByFS4d903WKC8aFcZ+ITBKZtAgmSPEakn2Q3LswNUM5kxujIf8oBZdFiV9XivF+wphaPQha8r
qrVVh1awll9E1IfXEN87JBDQs4w00ro6dN2k7KocNC2YNmwK7SvaQqlyUesMqrCkHHhbUQs23RrZ
OZQRWl6kJ1SsF4bgPqazTo+9TlSVeu87GeyQmi3x+1m8wtUoCH9+a9HVrTyA/t7dP8ONyqWJ6if4
rhLnRLLfLNh2kp1ObRfjflhJ9ROHQ3ORxxeKPze+qIbfMI32JijFWgWUjCJaTtH9Bwny0SnJq4sD
m4NV//qJgK7vIarDXYWlFIFmZN5ewAj3DoTAzaxz99zr3ITMp8ACIhlWr2cnJK4usKYR2hL6Hiby
dzIKx8YsIq132gNsSGSmZgZX24baF2kWJoU359y+vWAGBb+tZbQolQYBomLdQdxfvbbaIAV+dI8V
91vGMZ5Ym2uv7kiGTAo/UaIkAv5yg2wP1IypSWlgJ3NMX0ZHG2oekA4aelQE5jNLBnBEyZHmjWaT
a2forhyHoEfVQ6SvJ+wBaFbiFWe7JIrC8NwbFEqYy1k67w53a0J08mLkPyx+aL18hBvJvnYURyGX
Latk7/okhooz3RDQEh3E+Pxqbp6QOWvCw0q+K1x5NoQZBdUTkX2uOGonatpdpgPukpDH8pMKFleq
2mDfrdp2647y+rhZOQTGAoITlryEEqnRMlN/qjsbjV1MYnMEjD5m5EgmdCJAAEays8FECYU33cPK
Efiy74RAcpfctb84nw44R1cJiVpfTm0N+jvNGToeZDXydSS92T6JBr1JFpN1446sNjnRp3jECU/z
Gtaep8rRlPZH4MMsBmd3RlwZ6PeaogbLw+ZzSpv+B0JnD+gaz9/R89s3PwCDS3LAC3YGxqul4ciR
6SKRasdSzfNFVOBNjNsvQrYEkfmDj3RgZMd0O0cdVYDsEdCgNU9Smj9AjdDbY+YTsmzwbni5+Jrn
pqCYYHxqsAzuhM990/efOHi3H8arU/BUZxsmC+4wBvLqFFu98xD776RxCirV6e75f/hmv6yovBuw
0RUJEGpphmS0uqGksuo1nNyWm2voGNqp+U/jkV87Dmkvgfql/yHdPj4XVtI+EvTT3oS2wHzyBUZO
5snYRl/6XyEBsR6TmbMKmU64Vw4JhgBki+8WCGj2L8ju2DSVVk7MSnakBunP37QPlD4Woq7k8i0i
oAfV8cl7F1sWRXalhx5hSRvTTYEoxjuap9OMZFkLZoSo3DJFeKXvijVm6KqEPVgMVS3JWkh+GJVu
z17ma9rZmR2CndJCqHGgleqC//6pkk28HWmipyE9ZUBqptSBogwSvTiYIEmB0JotDkq2Vpfi3lv5
IZU0PfSOsfGlEEA/t507hj0rKLwS9T2sjqq8DBm4oFeh+TEsrRHIEySjhlM0eBeGsyfa9/owS/DT
yLqWCJOmkwZFoRCw9r8+2jvKqsq+kh6w5Rjvrc+RUbxiXS55RpV8nDvZo5L0NQXaa95PF4qX3Rgf
PsuqAfUUBbC/3wsnrCo78iovk3Gb/od8pTK9KuB57Ktxd/U9+DMsUZDrpxqtd0s97yC0xnIgOWvR
0P9Mgl8SzxliFCuJyu6/q5TI9XDeA4jJ0lSYNUGibd+im+I5+b7M15d8/wx1EuaGrNkbT+U00Qaa
kujLxZI10imXQJFg0N0ginUEuLRO8dERLN2sihVI2cZ2AhGOn/v/eGJIxPeFeUDH31gOxdWjMvPS
QgNICuh62NapVBik1Axmw4M9++q4APCYmie0iV5wxF3JCxVHKVoXbpLnTYP7miYfLvA40a/m/Omn
5ms0as+/cjfdWySvYZ4OqKF9k9iBcLs38s8lyf9U6b8C0spWicXWVg4sqCInNTTE5HTJu2AgPfjg
5Ynzm1n7ATOGN0sDn08zAZoSi6FsbluwsDg7mqseFdQ9DhEHSZi96E7jRRqfvhjiGrJGrS2r9OT6
LS4KYNoHlmTdMO5tc2ZJNTYKOeZs/GEz0mS0J9DhtGK1RXFEc6DyFmFFQqhZo2e5ONLxe3jTF99j
7MluIOx50QHRsmJjV/BJn4dWzORwYqKhGIOn+Jr2mxjUGMniwtJbkOvj+oudwoW2Ca3gAgrO9sQv
Z2XUjYC69splicw2OP4qNvWNTic4hj6aaDSbZwi8m0mnYfHXKyRywXLw7ZdlvY2L0wwsMcUYRr1g
xgk/YlOdSGxumBDeuShPcwkddRKbypnsmzdEh9BQYkHKMLh7LRzVhwatSXlw6JTycAoOdHNoG1a6
7Zw53wkTrqEyi6lRQSQD1SQEa4q24DYLvAMCVBkJlXifsK8C0ylR+IE0R++dj9dQQ5r5dTbcu39y
RfVwsuloPBPxSxNVlPv9bAmdT7LgI8Np0BLXF8l7WjqrwyygljaIrr4GSOZodooNibmIPdK1/xXy
Muv40fZuhDdKRDsJsGLcjXI18E+h37turiN1f3xP9cyjU5oTdGUahaRd0Nh/daVVW8r5ZGk9/D0V
itLe01Wa/ke+nshUvnOS0Sm1o1ypirHrrNypTQ2TIWmD1C9PGknlne3Ehx3dzE9NmPTvn/M/SgTV
y+q+qiRdro0PeoH4t3WFNhfmHukjGE4mIDqxDK3HJltXiF+FvAvlcSzYkSAi4ebjI9V5A/b0RNKz
5eR7bUz4s5ALg9d7h6+0KQ9SLReuqEYW9TkQWRq5TgrJXH2WIMkdBdhnHhEFwJwwECIfm61w2fJo
njnxf9pd5RDl5cpCLzYuRfoCth5ObJpvSO5akB39C3qZebKmIkbNMV4BB3rhzKEU9q7k6QrI5CfK
R9JAXMeeyDO9hcwAq4cCnP0H3MIBl8hRq0pVuExD0HWxHk15YdF3zOZSDM3DDTbCT5O7hocsCOKS
NgbhWoG26Wpkwj61HsR8GUG4lMM3gabmvIVmsVvZZ6I5BUWQgIkiYYAlT6shUWV7FfNUR9tPIT3T
uY6UK1nytmeKayqUDZbSCgFZckyio+GeanJBmfr+A+5gbnhHr7fGioi/rJbTftt5Kk626vO4C5dG
KvCj3lxKpyCzfVvEbStb5blatUYZenB6wu6+bfkGYpbR4VD+zQ3CuPzgct+vpm/eRPnY6cLrrDbY
ZugE0cIs6Z1x/zgoK5uOjTXoI420KmbwxutykbGsyrZU4dca5jGlHw/ahIPPJv81UrXBeJENu/q7
G4zBsQm5ryF4PCTJEqw1o3s4PVH9kltTf2lC/0LtswLLqf9DM0mcehCPwCJYNQOxd+KXiNAR3P+8
Be6eExIAf9I91Y29JXRA0ZYYKBm1tTcktjYTDokewV2MLYA8v5H8DLGaTixRBIyppWY2XizmPO0O
1EpGiti590mcNCs+9gwg+juTbAFBlfDjt6byukwkVvMx3PSpohn5RliDTqg9XvuZQJhuO4XMiUOG
7Q+hEUyUW5LUT55CF5HVTXpWwx6O/7k10HUo67SI6le5d/1tJvf/poFPvj+nditwcWwGFKggB+iK
u6B0ejTF23Twb5QOW/lJoEsSZXL5AvQqPyhyTlyMdC0YaZjEJLHkS9eyqBgHlr1SemsRYCJSE4jM
lWI2eBHBlQo5u+KuNRSXAhvObHmiXjNQxkCMVlVFdNMq0JsNdMqyk5tlZnxd63cTbqrcvLiQq/fB
7FvCyP/lkFok4VDQCV2yQZWtqGL+Omk0ny7SzclPISQFWP//Q+Zo+wvTkQiXrm1aMos1P4JEZhBv
syb0CmsRN8b0wb9Jp46qo/uxq6H6fwQLDj0NULEat6n2Zt6FKIFUHDeGqO2YRzDj3um+yAxMBrrN
VOScRGBBLMfSxU2U4rjjlNhZuGeggN71MhTJ63nW3eSsmk75V3CG2uPSOSp4BlpOKVXv/uqZhVJ1
eWShULwb2uIqW+ilWOvY3ZsXqAiN3oHel3yrjY+pfns9QPGEHaht4S+/vpHSmZTx2kTfyHxuKKj7
feXwKa8wGPe0tznXFfHbiCOGCJQbgL1lpbiGeKT3/W/6kSLsNxjpFvmyoik0/mEQ0yg4/hixy8Zd
hr9yv1FUk89TJ8w7PhuE5MrH/fAIEfM3Yl+0Xm7XJjp1YnafcCuolfv6JAM0AZaknO0dBrchanb9
X7YcSQyuHNKOXPLDZX+N8GadBda30UYILQNM1QNSLvVM6IpZvVqdvjihTXsRvcXw2Ajvp3oESI5W
dVDvCq9KVtvHank0RnR5eGGsbr6+yzd5UcYVnvfca06ww17UOfucuvKxFEaxb4iV2EjEfhT/hTGc
hTITsKMiHKThXcOj1hJeM0lEui3EoMJPv/SxQ7/rbmpms4UEDDMRR158xAETmInzjnmqB45q2eWn
9eaVmLtNhmES31vKUpTD02Li7Y5A2QbJ1MQiV904dI6IY+3OpgsoDzfvf4XZfomG6yin8vpX3V7e
MyoXTRhyOHF9NrO0Z52qn8plfRNBAscVj75Q2O2HfJxkob20mZhiUA/uxnl3USkXdBDbG9ZCYXot
nC8tj+vHDbF+TKUzdsQIBBl3wy8+JcrEauS8h+lo37Sie8IuK4Hf2FwuRR8t4jMKRruPoiveD550
j6nLKP/9aSt9R+Js3nUeYAvhxP3ENCTJDBFFJU2tYJqbzf/KIg0PCp8tpoeslOzNwGvSbah0/EXP
6DbdIalm+EcEn3T0Vt6glcvN8pka9nNJp28fGmEj69qenBiBSxKtDqQUYyS6DbtWcp22dHL7b3z5
cBfuWz2NxeuuAORKNcU0jGHp4haf2l6tdJPRty5B5zHJiOFwjkueeuyL0XJb2cDchhePszKQ8Tk/
0yjNzaABlJkXO/8WJ3Z7ONYhMK+kmKWRtqiplpz5edBAkY1IYCiB4rzNtffWsMb+MquNcJ2WHQZd
lJzqQodM8yq+vOcT82hp9nlIbWY5PbLg2sLbE7ElQpY581EtbGLNf9XMP8WH5MJf6v/gU1eU5DpC
DKISHPJTYI13VKQQ8xvT7VuTIQgIwSGD5HJwPdfnertsZlxQwWYedZPgjjOcdCCX1kNJJdF8yF3B
3VXv5wr53AVp1A5fBxqRSYUPgyvHHGNktMUpfLHY4vis4KM5/HMqXXbmxayEJjVqsIjcSWPOoYGJ
NHkf1cRtLmZ6r2ZeOt65YB9+Cqz5hWvMifXOkrdp00zR4d63cBkNbhZZa4QbMtaSibUzCAiCnObY
Lmdg3r1GGoygFUJfEoAnv1RuNa6jLmu29eSlSf2Zg26PkKQFWGJ+YYoM4rK+AxaFoGdsID7eqbt3
EIQ3V/8pwpjXAo3PiKHyEHVN4v16b3+NEJPCc65fPJIl3tfHQIr9pRv/1xzD4QNN1f3ycOPZ4vuo
wZDRk0elW77G3Af3gCTBo3EEzGZDP+2n2Vi7FFih+5D4v5TSJLc+yzp/ErpI7D1q0RtAWVBtiA+0
1wxNjhDAxYGt0W+5+tHkHnMQyQU6A0aX7fHy1RTFNQR78eaqmWHwBOtoXBHAVYQRMPwoc9SfOrA5
kFTJUE+SFxM+ZVH+t4xfJ+Odyru4huImb6B7wc76DvpPBKErxa5YJhVyXmoW5anM52n1d83y+hr+
ZPCMB+UfwRGcWQo8xJX/kcUa/Ecqnt1iEEXfBxc0G8GcJ83MkdavhXgulIV/oPiKff+8Lyw4Tia6
YL38H1ywrgcABSRtcWwW5Vtnx3zcB/L9GygpeUHPMo9AvDcmjMoVOSwefR+4UGK4vi+qsKKXh7Pl
rJIlbxGHajawgko/tap3QoeHsulKQx1X+3LsjTUoQp5ftnLdIAyeZ7LQI0mWfPOHDnW4P/Zu35fl
XWS+1VogcHtAsHRR1+B70hhPYD5xwrXL/YYwQvAkeh/dJ9KQZUJqX2xMCoagE2kLWPucgp9LcEGN
wtVITy0w+v7yDZfi4DKwt9okLvkrFnAGh5macVcFO8qfDbPX+NRJ2k4SWBEZka9uMy1JDAm3U2+F
EIgjJDb/G9hpHAf+Apw08l1X5suGENi8ZZjmqxBFFsAQjrrWzZR6PMeWbGu4bk7+S6ko+MuCL9N8
d8xITQ967vs7I5RnHKIqlIGDfw81b7ywQiHhaZKJ1px2fZCEhFY4j3wGQdS8Npsjyk7CwmttXHZE
hE65Fo/fRrDTVTe+bO1wl1j7JOS8OpjZTZy8pReiXCWhDTwru06DGwLfTirR3DI65KL2aKFcJHf+
u0k+eDerQ61Jtf6uddI1h7G0IoHSZWokKqwWaPVtEQidfNYyG9GUpBdjA+YCdqsatYtDGTd/vWn1
jrKiIwT5RDenP8PohAPl3XWHIBIH40Gjp5VVOB4pPf2TUCHUJYVzCn61pGpZObRIJ2JjR6qeyeNs
suFpJJkmPsLPddRVJvMpD7avB7VpMSR13sLJE6NsqssS2kiCahdH2lMlxYuZ/xhj70mqEl18KsTW
a57AUoAIym+oDcKL7RL4y5PTPDndv7m8PBXRvHl6WVpuD9biiZnDBjMdwqLrSf56i9VW2g781l/4
dh/n+Z10PAILvyNyuNRC9cp4u0dIng1cdJqjgBXZaN+Nf4PBLvxbYACMTKI3+gS3ynxQ7M4EVhMt
ZrFbx7ZE2ck4+4Mt6vhQF+T/F179MOKLWZBA/2gLOxBi6JTcROwi4zc2Q8urtficF6PTqpDVdgKg
HuXWdi16Ewt1lv7OHdAaVG8mPh1pxSO3jF6V1u7NEk+gKkXAC9IReQkpaiEbueuJIwc0nPoICifL
2OUc4mC+ZbtZCtmls5ZJTpQcBQ/BIpl1eNy3ZYd8Ih+4+lc9EDar/uzQH1r7Nst3BmsIGe/PTrBU
RS5nNy5S3EKz4C+Y90VbbtwDv+ww/e1id1/1v619t9CExZHeEfmxvwD8IyL3nT0EFt88e8oKIi5L
qjlWG8iVVllI3D+iG6Nvciv5zt146gJpdpg7wcwqXsb6g4qBF6y+g5YIJO0QRi4CId9wt2OfhTz0
xMX3jPPUu5qQK/4dPjsKCtD5qlpDBhF4DMnpxVNS9rKWbb6UAfYRTW7kHVexJYp/9serF+dQjBLR
dn/GbZ7tTbBkGRIGjUG6PotTCClKj/9NbLmHJkgfc99C+LmrnvFdwilGwQ6+2pN4UW/s3uAuf5tO
EhLrkeNxYvKt3aTuiJENT0/9NSheXnn2IDdsCbVFwsDIBYoWOGDO/Bngsx2PzjbIO8VtlXA+sans
O6B6XP9/F2ae3z8dhnprBUmslH6bZhGYANzZVw61K9rgm+FsUGz7CqXxtorzR91dnigdgiBfW9xy
FrnTP3JRm/e7SP/oS7b/hhupJ5crgkwd2E9Q9K2mtc8gcHXkm1L2s89kVMnHcadS/lRJmhcZ0CIB
YWOlJD96IcqcByv6L+wTOWYVE68b1+pXcXHCq5R82o9b37ZZw1Q0ijc7LubCgUmAe8BTNOd7o2TF
5GacFcm6KlysiUv5CdiZ7BHPxicNPBh7g37BA58wobfGYdE0tdK5EHx3CfacoQ9UhziyoptXx/NB
tFiSymb6pJOufg1+ozm4f822iDAxmH5mZGvqnHRDzRRkZEotwNyTTRdg1O2nOCsg9McCfAQYtZhg
2erZPfiEAnuL6Pd/NxZ+jt3o3PFz+0VLJfx6RAEZq/c5jy+nbUkbMH8eLLj8pS9hVqvnWI07waAF
42BkmSQ/kDtAXAR2W+cZxnaCLm99YITcYLifLSf8ACuNYQfufvJfBiyRftwcLLVOYMkQu9h05LWy
2mIj9q1iGPdaaeVpjNBF88Y6e25DcQ5FDXDtCEmkzZ03LcGPvM/jtInUklHw9g1Q/IU53Unp7c7l
0Rdz1CILfhaVmVmQVgoUMg2dDJkKcvFnhtkIMTNnXxcupfmhblbAWEAoTTcZYJKNrVXdNytgVRJY
D7WrP8Ksr/C70VhPCdrg5Tgszs8UqOsxIv30pmGcTB588411SpVYQ+bTHZ9BRclXeLtqli5Uj3az
fOhoBWZ41P7k3tNlKkqSsd9vUZGPFfdTmizn6knctWGxbYWpszG0exnIgL3jMNeEMQTZbVJ4+8pr
+cRSam23GmiaLdrGFRxGd0iApYhxH0ae5WJiRbFvfI78uRsONeFK12u2YiNoK8j/q5CTGQdNMm1o
ElnZchJO+QLCwhMpv0gus92MQftH6OU/QtxauwtsgXGLSqv+0w0oXYwNjH8C+c1KWQd3Hj4gjDf0
oa2qKiPp9QD1UppKmTKuyLnszBBkqPBoOdjOuIaIJ2rxAcckXzNwnNGYOgMbnQ5ZT2zS49Wn/Rss
iUO1fYuW2bb5zbBlEGut2b6Py15mWXQrSsjKU45Wi/QJApY+K+Msf8a41H6O+YAB/VOIwmvKrToL
KfS7yzXVSgU91jzFu3nt90zFpJWJ398TpdV9ihip+ka+Y5lItwnGBjqJCuuwrbI+arU1jEL/NmK3
eecBTRe28iCNO589MONIzOgqeJ8Z/i7ZFAbzJ40Lj5KbfTKWPlhBKP2Httv+d0WzftRzU/S3MoJy
X9EVmDmaxOXAjH9JeGqCA6/tt0dPVlVIOVTSVefho1nOALRP+juCgL3T53NKihAEPCOjUFD415Jh
K922F3I8yimDZvmxCTvpSK1rXBxHIyBfAwZh4JBuY8asgVmee6QAyb7bHkAnON7NmYfdahBaMNC4
NQHvdrZqDpNOkLcGy81lDvKWZvAE6e4ElugFEPZ/uYkJxS0vM+5IqpUy/q0bRffQk4bOk3eJVoMe
SFj7z6onxJfAAS5YcsbhIYBw/yPmFsOWvLPKMm0K6rR+Tl/U3sv0hJRx7d7WgfhYq5ZRvseXYwg/
UH0SsNhWcb048o0nASjmo/SUzhhWHWyBdR3hv33znWiDoM03X/IbO9Gg1s1ulpaoqhP8nZKAfE+W
C1Y9DrUjEPUs4Kn/A8dxT+eONul3v3KOhbjwKhguR7d1xLZQM104Jto1aGRLiq4ctcjRpXgm+RnO
AYM+SyxfbWC753xI8CE5vTvTuZ/zDMrAmRXdr3SQ8kJQeKmW+MQPwKdpx/vpckcw8NrCQtPzocXX
kasu6CKgeJx5CK6/s9XJFciYaSNj4hMYonJ+rMd0OQHlqPsg0ml0idKiUmepESfJL594pEKL78em
sTIAt0uMjMfVPaVdCAOnwwHXNroVZLQ39O/hBgD7C/IuibiyuoYQeLk2YTjmEbsxT4kDbYUlC2Ai
O0B8BjfHcXZgCL+jemt2oOm2J2ZXrSmyoSfb2mirEJ1yOcXQacjpzDP/nQq7jMSMFyRz+q7VrTKY
yC60POSBGrtwg0TSXcIcDBGo00jzR4SpUywDNnF55RXj2RO9SWlgbIDyHAjkY00sRMmCwXVSrxCR
9BkM/q068NQ2poOtgcA+mvCsmzu/xoVXQmwFgIMzOeMjE4RS0YtrhanTroS+oBFdygvbx9tJ4Tcn
GiZa/61P+qHWeZLfTrXmpY3dUSutHeRIq331mjpqB17iOZVL9CzxaD6NkK2gqloGVqtkTkNZU2KA
TrRKAmrRINRlY2Gmfg/oYZqj31YSsDkeoh8BXKFMWaWbgJ2WH08rxVH9PXGK4EC6Im32sBOvjHzC
wbrHzGVlnV9J4x/y6y79YrMxfZhcgZwzwiuSnvxwwn295QetxG9TDcZBpj1Ea74liZQM4P0TXIYG
zNZOIxb3aICSGAsjIlJCqBvy0vqd3FELMl0R4Q+8TWdNAQmy9t2BtVafKAEyHCsyeJwtfluB1Fev
d7w9DYUDMw+TYyJOdiaDFQtUQLpFNEO5Mfdm/w4BWN/9LlUS6l2AIjAFq7d3dyJdk9px9AUG1zCk
ovHmJFkiPm/fnKZX0Q5QCAkN3gPvg0GAAMMKSC8cyika7wwnYWzdrp+Fn2hs9UdnOV9LhXsNSLL0
3kDdMvwptACdtCbDi+lTMiXjsUt1P5nqBJpKbTLrb/Q3LsSWxm+ZXI/evCdTEHkg9iXFZ9GkoQUp
tl60IyyUl4zTGw1HlsWYUQFxp07xNlootI4SvHHoNsjHk8fkdTgFjufWm8g1BeygoUxJGZUfNniG
TWVzcPjrH2C2f+u4uGTFfVTZSZqBzDbKWKJSHxwiS9XlocdGKADsC8GmT213uHvzClYRnYOWhwkL
Xzeq/bxhUCaFWBKB0DKLNzzftLPRS0mBWK1LHG46IeRMriQuqkaZKdfBE7OB6t0ns6BPDXg9VUKs
013P1NJr5/fa/34oI1VvbUL7uEYZPJc5fSQn9bKOl8qQep5IQbcH7XBewrFH10VEiSxwcXwnXjGC
LytPwmsiInwPcZkDyeVfrCkmbBD7tokbTr7n3lV0XMAMHxPFNK+KEdgagvPbFnTghHeV4GSSeVts
6v6d2E9rIY2P09FEN1CwzVXU2IbHHenWaiKXGcfcB6hg6+VoWYDoylllH4ElruONBKUYb3s1/iqJ
Jpqi5n+5H1usBA1SzTFlezaGwrDh74Znyv8onGzkWkP/u2+O1TjnnXuw4dtPJxbZtV4swkw7As7q
JWaOh9L9Uo+fOiQXxZcTUdD3yxlWj+NhMIUzqmYmcoqhu9XUOz+6ao28aKjhE7h9iOeXjLHBIzmB
14I5Z6kwggJh0necWElgByzb6N/FaG3GOU0PvFJaOzQTT9nOT0HB4bLWLXBuZxX3D0cBwfifxY/u
DcHR0PzrR2+uEzKMPdz69RFW2ZTm7KAr4yAcviiaAmUE8e2xwKZ93I3rVelDGMsWm1PClhh8q2i5
mg4KtFSvdwqbYyOW97nKL3qFVbW9zml5HGhK5CCk1NNA5qF9pwxY5H0rKu+dqXE5MB25xUTQ6Rvr
1ARmUh3Wi8gTO8jb0AB4TU+/vZTVtgxCeY/rEvKrR+pREXOZIg/ANqAbq5tGccdWUCEihorOOFo/
Y0cSH3YM4zRi0VRYf+fxYLNNvBzWnz5dAC611FRPmniCCXQwYnj4vHBjepLf9neGu15OcpfGXnDz
8leV39YX3L3BPGbiTBXm6pVX/4RdjxRIafapWHuExelroz0QrmWT68X+9Z2dlIpzm8jPuyuZJauW
4pogvsi3SR14BMDm+JA0XZfAMDP9i7Af2FvYPic1hdNaZZrh/ViWUOYeLkOiKCkPaQv811xzHmTY
3UNwiPzCkU+pNv8/A31dlADKtcM0UVb3ir5f/kaE4dIgcox5nWB21fK7eqDjj+S6EY9Tz+ZA7x2q
xNRZ3anGS1wgMkFtR9H7Q7Y/xQZTwVYCMV2zG7pBa+P2qLeZifBiAjCZgs6G1rtZBwPXGiKudHEd
g43u883dFZboA/zXrLwKOytawgrtn9EagUKkZdAaj8PoNXLtI1GBbn9i9KEDzZ/66V9Gx/WvL7/8
hv1I4K73Zbx73n+Cxi+IyR6nIq5uRbWietktaF+cz3oZ7koCWfnviIzUoxKG+lzY6I0HpxVCJndE
uXKRVlsBwiCaOyc9IKZXrR0Zq7aQ4IKg8vzV5YZWbzPBuojjbCf6OtIm7xeNvhh+N5batPRla1yv
m3xtNOE69WEox/GgAkx9jQ9E1jWWBpIzNfXA8WXA/mze/WTFDKSbeOhhNJwVDOXNaEmzSN+khLa2
m4vW12O8jYf/5Ak57ocEXU++csL7pNBDmQRcEjSETXJ/jMdL2S7rotpPC7P5j9buUbHDG0LFvhUy
nOZ9xZYbESjDoKWhx5pNb0o4rI+PSOrDEn6ASQM0UyQqZye9O3L6eb8i26HlBtHeUw1qzqV58XF5
ter7vso9zUx6yAaIuaNtBMSguWxZpS4hAe0CkQad8b5kuIZqs+mnYC2abXgewLn78aoahai5fe9n
x/ZF/Ji0HXthgKaA0hWW0oXGshk1yt69UsXWDLEUTOj4HCRgKkCzjbXcuub0mcLu3KejlaxEFwC/
f63BLVQ/sJa8xissSBeIpRwYrCiqkcFf0tLAXI4W9INSTGOxCTakoYRQsWbDelAhFk5P1c7ksmlz
b4mHspoNSRmtPxNa/FS5rmdutRd5h9ezLUHELPd6VdJVoMXMt4Zvub66KlvMeSb3fSaAMRcO2WCq
4kzn6kGmH2xx4vhSc3nYqrEYkRnF5dMu2MDDwKXePll1tWzJFAdzpWw+ryeY8r0MVCGN8i1rXI1P
BPsqlvwoz97DPQ+oJrJTPDabKwwq8767wUerfJk9cgw4ApKJZ7g8FG3jO8Biku6Ge/ASMR0144NQ
3JPmL9/YXdkDl1bi+vL9vHF/BNIH81G3kbTmHtPReKgXk/CR+WXliaieLNvW9f094kJcyAc63iBt
jH6nPx/JHFl7az5qhBaTtqsEMzSv1q4ntvSh5lZKVx9KfCj8q3rEs8DTa7smfQEeAr6UwbuNMslx
P3cCcvcO1klqj3RjzocLha9FuW/SuqSOgMvft1LRzPexi5jmvzpHg6ZSNkstP/X6Mq0A1ZwKZGOi
9+9MbtTTDIeg5Mn/Q7vsQL2n8H8FbkNj7O0IaKvu8ZH9dNX0szx21j7pUpAstdyWGg/IAOaZM1qx
ne+C0GEavRzZ6sTuSUxlspa0tltmTgQIBPnopqSh8T99arwqny6eEECFglPO6u93XNQXoJJlmq31
63+3X8F0GFYddPH5yEY3tFNhtAJN2vS9qvcheqRt53MHR7EY7RtREpb9ixmv4JazZne5RuxbRrhK
vtMA9oah6eFrPxnou9IGIMDYa8t3/kFYEmcoO7WyvzZDO1hqjuPk5/JH/lL/74h4nz2i/TO/gcUa
9Cr5M8bHBlzzrt4I9J9EhFQGyHxjU8XQQGGdFMyE9Eg9BkIg1SqvtwbDdUwAw53aG4ufb46Man93
kAAbYK90QSHXkYNLdVgimpWNnSi1bBUF4tBuqxnMCs6QFA78MjwpXAnYF0ezfsw4G7b3POJdhBWa
uaoASFobHe9M27vWLIaIrh5jyJ1Uvco84Hrk49yoAKQ4sjDGCM99uV3zmZUbvcDyk90oqgutKnpS
T0zmF+XYkv6HlKCfnQRsF1DYcZWyDdMwF8k7nJiKsETABrk1Ci3NaJawU4fezSYLQR5Imw/EW1nO
rvLyLUbKQD6j2t6HhM+dVpCcU+ylcb8IR2QO1ARRZ9HFEeREOyMz8vY9soOFuFn61qXkKmMse0qL
2P8Yv8ie+utioyRZ1cXO9YxU5MAFECfYuCuW/9z+aRFJ9FCWCtG46GjPukcB/6nBkF/Y0aUXk8Pf
mqeLlv9WROvoxe1zyOUN8dV3L7xzq9UzzDl9G0o4BJ9Ath2RUCLksI8owXZ+vmz+WX3kDkE4RB/i
WyZoWGP6JJQ4x6/CzHYVHfZk5gLcB4ICTlZYHu6Y6DOW52ZufsgaK3SdGP+xDth0nwuoGag7BO3w
iupKCGLemWmUV5MfzqAur7RzdwP6P5GfiU3QEpPa+cxRzxOQ4KXc2W2ghNfYroSgvBgCV91cGTUg
fMpVE0Hsiet4JJrl9LV72rwl9BzK7rVpoiFTerkctPQzuZTXGLOC0UYf+2rrAmo+gtuQ7zaRY0VD
NtRJh0yipSKyjy5z1oq6PbpbUzcqIaM94nM4Q4SJZtppGXnDIqzCUvoADaxbmuQuPlRw875HU1V3
2JOsN/iWDn47tl/6jyuEg7vU0q+IWeAhd7TqD2e1zxCT7pdJsRrSAq9indDA4QPynWPd/7Yzcm5E
ZVQqyWmsJzGOgxG8eqpOrXZ5APrGGVb29vSDU+6v38/V0blWZBD9EjEuSA/e0WF3cVTU/VhohseA
nqCpWvblNa2J75ww4h3H9usAUMkY4YhsBh7JV+YSPnPkAJYrN1Ec4YDWxkGcOAt+nSvVIp9z2jw9
EiE9Bl3BbEkInOg5Mwlf/TTgQH3pERy+9CHBXlY+JhTPUgrUjwlHS9paHs1jRsYtzEj8ovHjXIwR
17YkKGDvRy4jBaDsBJi+utSSsV+sHnh7Gsv7vaCyKu+oEBD9T7+eYLfwmMzN8UvqbhzLQIh0PgWc
txOuWFwNf7X44WN0KzpxYY00Ulx8+Qdw5W0U0n9NBatfNANfw9nIZmns+zwKSgbOsK+f3o2nxxal
vRNxg4dGR6hYjApYhIif6/ViNkSjVFtEz+YY4br6VbXfscdf3bm8+47deHYTlkHawbMUsI7kKono
1+Y/9uDDKDnmH+aQ84yCVLxLpHfFXvG2n7NpEgY/WSOcCOjD4NgaYjTSAeM/AmHVZa9QlvgdMXVh
EiMv7WCKbJqM/u2dXToz23UH0rRpq9a7lxWtBwpOaO4EQ8oVrJ2RpDzZJ/ueTMpmzGYu2herzdsk
wAllDTiN+aT+uMK0zs7UbPdR3OruCTq//b8wW9N2pmttSXKxkIAR1DcgR4++D+J+9eONIl88aKvY
lYKZmuGYXYU18Qs2rBM8oXbGoapHpEUalky/DptPneIDlERu/owY2RQpFIJfYolPnrmLjj8jiynu
XTD9kC5qm5ywnRBVKYUGaMKfFzksFZ/dxQzTxrcicoCA8hifM6Cm05i2nqJxJRujm1/Cn9kNbF4W
AUupSYNTB63AF9GHnzpFRL9Ao3shv1qTdqbRnFIFO2QNp2Uie2JudRVBqwMBFBdiuCyW6fsHIISL
EGEte5h/xrdnnIfUdFvF9Z/Hm/0/utwj3R2rbtu8ZinwRVK0zNZ2VrAAcCAVmLpsdBAw6mNOYr1H
5NRcsAIfory/eFTxgTU6K5asjuzMPQM++7BoAbwHy1qVwzMDxBUwNLnzQxTwBllQxM/bJZqbr4Ev
1AdTcptBjIpsgpiNnlzJNZmcfZd7zoih+smqSr9f59Z/pInh1Ei0DbFgSRdbCJCVBpYhn0JkUMI8
7RvFkXPU2/kz/Wrx5LVumU9tUOdQb07W0cTpURJ5EFFWQ1ZbNuOZ/WCWpKrli28UutxUjm9qMnVC
eYKc5VCI7SYkXnsXfmTR3exXZ0hspWdt/7nl3jX7pKBGXs2pMPL1sCot0cwQXBARABtzgq2lO1Fn
2tSlDL9oegTYOe4vN7T+lwYPQ1cFdJ+poOgIg9aLy90rzjxbL3Jcs+s0lUioztewHeIEImwzFmJO
RQ9fcCgZKk39o+bR3AUBF2ZnWpTClmKLcvnzDyh2GCUl8PGRRjkPL/geyW0yIuKjjWSgF/xrwXPi
XGYGABKGV77Nv0vSJk8I6j6JFQp1cCQedcjRlQ3IYJgrtvsfMrX5uSoAqc5qL7O7Wk5atiLUT9zi
SpPzniSmy07rQma8pQZMamE//kpR1mero0EPAE7+J346UD1LP5h46t0qtFFeR4fK2Hq1+uGgOs5E
chtwej+rvrJTau4fmtdbVeHN3EAsgRDlismwVSx3Ur1d4E/9HZHwII1E3S/5UkUvIb2vR5BfUThU
RTxao21Gu3owS1Jfnnk9atJDp08Vi2qt6J4Czp9mAEnL35D/MecTRwFcmbgTcqT0WQJfrxhBDOzi
hmFTgWT4WZwZu4TOnv5NqEkMif88VA7JEpRIy70TZE3rokKd+t6zmlMaLkJijpacU5TIzX8KaF56
OtbrDV1F+KiPl4nsujoxuRnRTMKdrgWwQNFC+bt30wdlleKHF/vRimqkoA8S5pmV02JsRu3DYxVy
V2BsHcDVKPknBd2uoWSHbF6ofhtLU6EIVlK96FULqNhgzo6iR3n95UVvlmr9tEU9IP4pDY8/ee1d
2oVwcYU7RKOnHzSJv5AZUe4LAWKqBeoR0s5VRJtm1wmNCEIdUjeaprMSgiYRIo5ZeXFsUBKSGKj1
ygfDBhdUPCjB2f8r7jSOmwvDGnVI3soJYGo8ngJFOni6tqR8vdKG+flx7wkZgT5e3arAn373V1ik
AHibOTwBI4KttquoUwayjGssBROFsShEf36/3eFfzMnnro9BikTh51XZkjW/j5GmHku6E/VKTRz3
s7qkK68mT/lOn+qWQBpFVO7WIKtylzt1McwNawgJO5BWOktBGyvfRID00IiUTqJBkoYYsuJr7RSs
b962Lw6EEyiI5j6cO0Ri7+MRWMXZB98t1SNgqmJyaC4SZZligL7H1p18P7IWc8GV6N3NVNQNcL3j
qqbPfu9TGLi1ungat/6HRRRwup9+aJ1Slws7wVdimsU63fXY07y6MvTYYKKoL7oFY9g6BwDnZnBm
uPJ0uEO/AJOexM/gR+wLZqqBqF2tczrzKeDJww9kxFzNLyU7DL0tUQwhIq2mbL1yCKvfaVPIDEUh
6GHwVJsP/vvutf/W5IteQSX6rc9q49ohDYvwPQGN6XDezN1H1VOyXRjT1+R6fNehZW4MdchpeHD6
mjvRPFWCkse7KvuFZ9Rz6VJ6XyUim4EO9rwWHzbXNOKtpaRl0ns2xIZ91G9F88R4K1muLZlQAzxF
rkbKPiWTE3/Cywb72uxg+HG9wCHV6zl/3MyY7xmeDmwOIVck4Y0zmMx/NGMwew8SqCUA6JcVdiad
IuDyf1oVMPk0PKOdOIVH771+AFkL6D6HSLoVOsN4nIhrRadIoxoMBWlazAHGYAesSafGIEBXhfMC
a0AULD/XjwGUOqrReEV2Lgm4z5Z6KIBsUsjnDvKYKAA5pj/pNIQUZLWtmYsF4+cy5VRHfwV8/K5g
OSv1eAFTA8nV+0KZ30NlS/EZlpIXyeH+tZP5TYIpKyR2AX5c69vk+dDAyWb0ROVwFn09tnH1/329
BCnRnwG9SDEEZSq2GvSg698XJMNUyhmgdweeIPed7IJ8ZXKQFE+PwN6F2LiSH3QCBqu1RXP9TYKR
BfzPw6pGUuBdJ3UN/EB0CxJp0Z+Tenl9UTMsf9FEjOeWzOR5PWROACKCMGgwpkkmUlXaCwykJlYD
AsA9eHRfO/ZElERj/u9K2yhx+XbQquJ3eX+KCcFF1WtShUVf1ubElRwvouv+nDrZEa0Le6Uf/5Pd
ProbhkaBcqgidtBmvUvxc2ll8hL1wG+aoB/2lNg2P+9k3TAiK/YY9q7f8ro9f44RNUIeANEesCMN
enxnkYol1mnJZCij4mX4PbDEcMIHSduB9FADKvHBgTuXXfWwMScJASb3Qo8PO44bxbrSYadTs34C
vDKffuMJmfEHGTUfiCg0l7TEnTiwSOdC8lcYCCJisoP+OyUJYWK3EDvaAXkyGrqlUV7eqZHyVN2G
FTgiyV5e2NST+xZyiOpAjUVrWRJ2lsVESdPoMO7YjKIvUrhveE8rrF3P4sZuaiMgJrVyzk6pHV9v
kZDmsLAVd4Z2ngD8Sh7XEv8T0iBqVWA3yYaqaVOxtjug/fdU7I+r4waCe0Fls6ewdTWCo1vyTDpV
dehq2r0pfXJ+7lEqdMM32MADliXL+XH/fLIdhYUMezOjCTg9MhCL/PzTr2+xT3yGVOljmih5hw8j
UF7HuJnD5TM0/ivkQPoiSxM4Ay0Hwrxck9PDbD3Y0d300K0ZpMl4m97SGKYUpcEBa7Hh/pDpRp2j
gRDu9Xu2WXiJCyeEqblC9CHV54ZXcSBNDipCukcf6y5ewecECYOBokK7cQ/xnzxnLpxCOHAtWzZi
PoUMqJRVBU2CrVKh46lCcMWpB4/HkQHtkocoIpf9Xdd669OxfyottP2RYjzLV+J36v2sBowFqgtM
y4ZQn29oTDD1qqRGr1wpWYAvOOWpz4kWZxNZPk3m5nhYgU+Q3CHvX9NwbXbdErhkjbnHRZqPEl18
bW6uQCZxt0/gds+q0xnx1sEdBDp4YxMIg+OoqxEwauj8MtXKb49SbXmllau3PeoZdv0T3eHfj8ns
bSYpChm42dGZ3yQgibriiedq+GPjI3Vexn/E0QjTqQIxHhvD9azq8TVnFbs8rFUWMIjGTnRryJAx
tSt7QQZgDRx1Oa9kRn5rYai5Y9eOHqEeZl6CsQa6gyxLAfDLVmVX3dH1LtjUgL5i2dGVbiWHcDPe
GDo6BWjPpiwumaOuAH7M6QbQA9BNxHx0+3EWOS1JQnA6hGXb8QaU2jJDuL5ETrhSaqReVlj2Elbe
vCWqGaxQOeg4cYJqfGAVOFIP/3qdK7pyqWB7Ekkw7LM77NszrwDvGUEBhtHHRF5BhvhKDLkStPg+
lOs26ELAIlqDhMmm5pQVljVAa1Kf4ZkCbwyqwq+zxEDRNA3NTCP+bEUsoWC41BnH9tptrYzxJCzz
H6HEJBCwD/ZJkni5rstoUnfStQgdZrRF8sq52yed8pB7iCMjh3mMqxdcySzzK0lx2udkmFZ2LCiw
glUldOSdEaD7JwCNZYJj4cpOAX+ewBT8RSyfbiIG6vG50kOMB1riL88EAD7ZrorRkVa3LlgoHWwj
yeOR61XRBQvhyIyZADB/Cfnlcn9lVqyR86VwEhKo9UXqVPC9pfMGPknjLyLaiUTVZNan5PIXX2hw
5bOonpOL/VF5xRaEhq2YQofk2yzS43zMviiTWdc7n5gz+qQJqVWbO0/uHvzFXjdwfUZcFXoHR+x7
8t+qXaKJhMixunJgz7H6C36R9HvxI7Uln4TF05WWSKWk8VjUJ4HtRKFZcCT2KiRfsamC9BqYSi/y
qo143ULk25UfUUw/4W3z7cn+TwXqcpyH1NqqHe714RR+/CIa1xyCP4s5lnU4tfGVlNXb7fVmmBbC
gGC8AQEXOvOtEtSe8AsItuaAIvKymfAGGkgpTLljzb9h3uUwUVNcFI+6eMe4G07MmAzKYA8kPb4C
wRRQX89dhwh3PlvPtnq+hP9ZVEqv2mpRd4/YC0/wBRKcH7lIR3cuNGfLYyF/5/rIYkwZY+qNLPsJ
JMsd5vZ7aa3v/MAnhNMFWfAX/+ueWmgUFjQuyHWyy95A8mO1FabO5W9uAouR8OQwfZykmak+xCXO
OlZr21/dWY7RzalffKQRnzXJ/52ru0N7aRbdRDRJSN4yy9JWP/hBJwntMbSLYbU7NTLhneSkPwVI
U1odVpT5yDU3sVP96lyTFNM8pOnwrPZAJNbQcUm83SjWsUM8joc038v+352xGQaC2UvC/PSdN71N
xUISXQVrzaufH71yLCKlb97xgnh3BmYFkxBf73/SHsccBrdNCP4bSTuXkGgXXAvchFGgsuYF8nIB
y/rCnTSWnWJYCE/p5SpQDEQ6hOyagOpeDYjIw5WtTWdzE12CZr+K31MetAekCoo6bk9TrkmG0jWL
j3AkoU6WE860ygtyUGbbfoBX8dwFetMrqNHcuz1uzLrKEMQ18hSJlNH/HXTqlYE0IxqPifph/nI1
iCt+KIc1TwavycF0AvAkUVCLA1x4p2xUNImiVh2/aeMXXIv+5NaNLILj1BMHhkVpXdapk3TX3j92
/mmmZDWVkcd5AyH3YfI1+qOknGMU66UVUPbdpie0bqvLEPyUAUnHh0tsnUO2oea4biJUVm9/heMN
XXuB864JTkRS0ll/VoErL7tomeaA/yLmAf9/tMU0CdY91sTxOvgUDxV2IxKZq5chywfrQydZ8RVt
ByQHfsc5hQdfmZi12fxCVpg0a58h4Z8WpJT4QmXJ6YGyXOwXgUTqtamQtvcseN/nhKS+wvWlqF70
K4Xchxm88pHl+mbLQdWOiQ2jmxvHAL7Nn76lQG13uocuzRlevZv9pPAjcY26dUURTziK7/3QUkWr
D+fIIm9cFFQzHkfihDEQMzygv/tj5/6BiowFXb0JOYJsJy4Eb86gSvb8I0q0eOXRCXgTT4kJ4muj
eUT/Yqt0QSuphQIJZTLk19uVLGkew8tdIv+DnJ1jtTGSbzwmsLZFe6aq1Mog/bKQE3RX6v94bTZ5
d7J+iGzWIrKvZfIYRyMK2BLiYf5s4u8/mcNm/aSBuK8+7FkAArVOfk97phw5Ra3aA1snBPjznn66
Gc8qbAcaUzsBEhWcnGd2rKczJ2WOsKGLDHje99m8N2Z5FYzutQHInPXmMie7u0YECVasX2sq9Qp3
vSU8+uHT52cKjDpmnBEubf7FE6bMBF+XMV9uNvBgMPcDR4a07mDRCXIaYzXs9vLpgSk8wtkj5mWQ
d7mu+l7oNBUCPJKsiA4yKevYlC98O0nomXB2fh1JEzrDK/BWKosPrVjcb5iCouZwh9r3HmbSjKGx
AePzTHeSrH0XS3yCplhFPM5mJgLV32d9IV9ES+VxieUrwp1COw+VUtDZwTxQaPGOvrpeN+enwK2Z
a8cPPe3Xx4tepPejW7Uye5MmzPvnJ5mHEHYwp9ShPvguITpfsw6iJzfE2EF6vlQKUqeL0ybdTqoy
uZa0epbBN8UPpSiP+Tc1/0DgR7v60W/3qaHTMY3Z++EBWSkzO73WQzjYHWwv5QBiC6f+aXxrppuU
JZG206AtWjq39LihbRENVun3begULNLBq96QZ/MthqCd6WS4afDxijkmyo2vozdJoQVbqglHT7qH
BP8Q9QlD/elGOe+BA7fbTIvTyD5iwd2lW6MzdYHUb7DDNBmWSaLUIUj1ixFSoa2K0oX+i3MgHDps
ZDItW4ZWHGflODxD99WxjeXJT3oDCh3m+PaLXQUFxwRadnpNH5Ksp3xPSx2WVzF8QqBYwdC5AdK2
rKPUYYx4zgwbw76cXxu4Zl+RaZqXFm4XjxAig8Aw57mQr76qWNv0FiPh5zUp5+IUFmWt1BwMEljQ
PrmY6xyk+74HEa1TrXD8vfaUPVkKnlr7JK25M51tMG/3U8GvMUg9GFgVpVqRZJPQD5e9yNFkCoFu
5joRdm0hVu4LHkxLpSUeXgNvkrY3H4pow99R9Ha1yZEAKOB43PWWTNWFJP92sreku7tftZyz9jdV
8bQOfIHBVX7Baj38USDqbcQnlrL2WGixUOPotZt0jxBZC3ngNAlOGZRd3Ixr9dY6pWl9EigQB+tb
f5KbKctpoOtRIWazOIxg78IO9GLl6LbcrAqJtdKjPdrV5MgK6R645Xw8sO5iMhfou4E81c9gv1tO
BmezSSgcWyIOpT9RKd/gxeYJBu+2gi0Fmazeb68aX082elOSwAEN4pgEsyr/3UnWMD9J/i4jYnc9
OFCjnx/kMCLMZoKvhn4aZFbyeJXu93mEStZBBXdAqrtcdZ3MxP99aR94HrdWFTbS/LKp7+xjbzpR
gujSAE8Qc34EssNUvhJz8JjOc8I0zqbS9qw0QcA6zX2WUX9R3xG2mOZUtqVMgLTzGYUeS+UdIEMr
j0NeYJDmuXpnh7atQh3CtO2Mf+aXfgwD4Y78KIs7Gn71P0YB2KjWzzmd3hFUBUFEQOpWkA6wU4lq
PindAZZMLKPAgoE3Y5cme3DhXNniqBB085OX0vpR502MUVGBlrxO2/HxNtHvmvwZ6O1Iht76qR2z
F6zqwBNdKQhyQDm7MfJJgOIXrmAAXleTETl1jFRD+DeDjBeTJDJyM3YZFIM+XdOU8fqKb3MgYeEo
hJy/ENvP2Xi8TXy7l01UZi3076Z6x5muzjkLh0S0/2vhErkepFK06fW1bNL+r8adPp6ZohnIddJw
/0FIQkqhT8IOAhAMl2vNXuZ1uomuRxKtKwsD/LJnxhFIy5KxRyE+TbrvHtUKMqu09ppTqI8zbebr
RoRv9BnGP/S5cYyiltVfqjroLid5aV8QR2bhamPAfBhrNwR4J5XivG57VIHa6UXT5iwT8Wq0OIBk
6kzdsSyvZyf4umMFfw5F+034+2JD8XQpEAXtA+Sf+xSWqa8v7AX1kAQKj08jebg88vAxgV7X8/wZ
FV+jaeH09kDfRO+fxg68DGgShMEt4Oqj/pGIdcIn0ANy6UDImvZAluDRLA6AP8/tHTPUffe/TtBs
X4JRznIXqBxEzjUjlPPLwl/Waq76VcjXHkLFC/SEDjzxQogh4SPTBkAJzFASOQlF0BAO8qAfWj1s
TO4/SE4kGg8s2Jt5ZuB9Oebc+gnDwrgylp1Iq0CAxsWWt6u3JSAx089IWtvvRsNF/PcS5AU4vQQI
jHAFNX0SlgKVV8gKO5BiTP5ge4fN80ugm6MnunieYyWKR5nkAv3yzClPVYzRkpTsSH8GD/bunDnL
NQugb2Aw/kWPTJS6B7mNYr8Y+wVlLWb8CPKl6Vs/nnBDl9wEV47OV/31H5gR8VCAnqmwXMUeLwDh
sWS63iIWToE19fs/bYFVdUvgb0ENcHZ3YTpd64YsY2Lmm8cucyNJFf48rL5FKJe+Dtx7iUH+WRpd
i1zzvEHmMf0fyt3VRqvnZFvX3U2NqfbwSLZHq49E3nG+p0ciBtflRXvqUTLOs8Bjh2zB37MkUnKD
UscuBL0RZJABSBxcZXQgapmvc11cwjLrr8PN6JpZZrYYNhjtXDLgrQL7Qx7Y3TAkL7Jqud4pu8Uh
NEcuq9H3aKBITPPJTEFM0IDg2Z3qE/HnMXhJLwInqV1bWSWfDX31cCbU7R5NJyyhQ2uM31IcyXA6
2Uk6j4BZcbjRqfXZ/I261gyxSwy45kLjQBWV8xBSCwIzdw1G09pHoFG09Svc3I2NqRaiDr1cnd2P
BCqzMebSdZ2OpQEgOlKU6w3MC6Ci0GI3r7+fbZUIfOWP43ojqlD0Ie9Iyhxx977OZ1r9L04VcOzj
RCbRILvFizsgP2ZVjvc/Rb6UQm9W+8iW/q/WU3dQ6XJIfDXgwnFg/0znMgdP955heriaTclAAaSV
gTt7h1W6jWWG+XchLhWrYedxQFg8hCIjOvPLar+p2075g4rSu8E9GZ+N6oPlPJfP6wGpijbx3+9C
w7/U4oeWhFzD39ZAZ/eKlGmDyzfWX0V4Z95oHrgZJ3cXd0rknwxSd08zshRrfW/v71H/CYOKlZjB
N/b03+iMBkiqztEiyTDWVe2JQOYNyvYWbayfUWzQ4FwNKaG/KKkNq4O1PchIOABvZpVF7T7G4TU/
nGQMbEB7l2AMqlMKkE+5V2J8zrzoitWVKs+dKnvcyTMplImdqmMTDNgUVwlzN1RjklHia2eYVRy/
jiWB5sugffPUwc99oPu1Jad7WpaQg+mD2hbJktqF+2CQQs9nDXcFua6fCf51fVQOAR3bQf6ZYQjA
Hxfh85lcNWD4X8Z2cCndfecbHeLdIW1qOI97BnyBnxeDRLlBJ7mv/Hql9uO0bt7YV7ZcVVBdiAok
/h0M1eJTTm9AKySmBvntfTVEmmRSI7DkyT5sCf1W/YPU5ciwiKwBXnedMwgh+1iT79jThB7ljVtb
u6t2jRLQ3lllUKP4coojR2XnObnqcz5S06EKQ0nsbsCilEAS3ry0ZrW2VjErC3pocIfypi2xP9OX
rLUXD6PwwRbeeyUdR4MDLoH6Sd51VLrqVHaaapmghDdpwrjrHBa2QjYEXEpOw0p1jgMaq7GkTxWi
yS2xEcvJoSc3Rtk0hnH/DQaDP8JBQ+L768G7VzLkzxFlbak9XI/Wa1M8inRzVHHYTOFUrIsQs9dZ
xejXcZbqzj8+mrSv02/KQsgXKG+pbM9qnTH1ZGLV6C7pILV0M3s9j8V78mlJGmhXfEKpBDsnR7UR
rF8dNM9FiYSZ/TxAzIIAskpVpAmIkmevzp2wn3ur9z3sU1OGhflqTBZO+XPedbvNP8WOAQKFFnmZ
B5nTImHkyXMhsIt8lauISNkNVYH8/aHzpgB5PPiSvG2RF8hQwKT7qk3pf+MwoqirzykEDZuNVGy1
8FMojd0QbIveZ8LJk1XDEDlrdhq8olGFT1uBUwEol9MO4xI6z8RU+QBfv42AKmvdHZOYqGK+9MSi
erEV99gVyXrkKjbVfyffeMCnC8ipOU0SaxbRytjsHSwAngM0NkoKS579yoTyymUjZnvzwFIuK5y9
ek3Elwq+y/7zdVMffTKrJyTWSBRtS8N+U/cWKfjrlZLveAR007hqsnDErkmODA1Z/Od9XtOz60q4
0y14iux8Ur7dYUjCbLkJexxcetwao8w3yj22QJ2/k/L1DWrQTzxvW1l7g6aO6NJXoHdlOLbNh53X
xTbeflhjlrusKEpY6E+JeQXFPLIvEvv29vXpYm4OVbrO9atxtkfmqxLpeIC4dCnFywbyJ0QhsVqu
MLcFmB0nP31pHvIh9r/C9Ta72/C3R6wX4rvdY9lT5NaDus9pC63MMnprQ6Tl0VJ2vCY3y043kIE2
16zyN3u5Mr/Pq1YwB8w43RFwWl93oGsqs1oGaWKWD6hTbg4U5QFkOjX+1TsXxec606n23dnz2u4X
ZmzG7S8QNGUMripwBuJLlUe7Q4UhxkqbwbYxIoglfFfaJBxJXzNzhSN5E+ELHt7We6C1g6zfO5gF
lnRF+HpI4KckaDsn+8ozZ6Th12K3H9LO8gznXqUmxn4r4LD/VDIjaMS3KQPFY68FcTCn4BZbqtoy
TGlW4I4sMXd8+bb55x5+1CSnjB3ZxrhzSfnSdpcvie3w2iJpysjC/OhyrTXcPsZDj/xS2cIM22Mm
nIWjYG5kEOi4dQa3ZSUhRS6LIbIDp3KOJvK9YkKyj0oxv011ahlNeDoHVxf2/FWLXnum4vIFTU4o
k9MGQUSTzMOrNlrZAJ3AtGzgMzXo7AcDXXDmQiyowDwAy0V8AqnwJZMn8WkRykVDVpALwYIrZ95n
ZV7SMqgKNj3FpOi9QNjfL91MoEul+7DGLo+f3QwW26cPvKbC9WXP7r2IMkZ3SxdL+LNAU+Tsb8pu
AIF1QsTbBCJINtHZjESKCM5XtjrcPHnH3KABeqad097yyK/RvvwnyHGHWf+sRIEdWCUg//DSC5LY
eLs9vvq0lXKtqqeRaKbcmwEq8I6C0DGaKwVHj/0LumqLbal7H7bC0tk+Yz4TEK76IcF/IpPYQBpy
orlfSQhUZlIBzbIrC4U/suwqZTTeIobmIUWSPFhtsqRQaBZP6I+p2NkQ9ksjzbsRBg4yAScswq1O
hy7LTJprZh1dZToPTVgj6m9deywQRlj/LsWRpzwvzcFnbB5ks82qr/KZpnqmS0OZtLfXcTS4Ap35
Zl660S6FQoBgCqHYgsp3ELp7q5hQVS0lvXpgnrJ5GXQiynJ4hvox4kMvzSEdpCL+bEiBdrWa0sTI
L0XVwiqt31KKdjBZPyiOc5A59sGEjLamADIBPFs3yAnWWITGGb8KbHmdXJQsdJv2oXPKi79p4nQp
sJPcm6ZuS3847GvQBE/Ol4B3ldPPjsNVQN/Bzh6p6b6LimuBLDBBG0AEJhmVBkRvAA/DG7EstFdo
IYcjHd/8JKahMyuwg3TYznKuwG5kENuLg+uJFQnVmqvzMkf4f/WOSXmrp83I7XP7rCjJXqD8fhkF
6PCnS/8o1yoSVqJ/STL0rdQu1jwx0QucFpH8vWBif9gfha4C6yD3CXeeqQkJ+6isNRv0BeT7wuSW
x+ya0OBTpCXXzrLpzPfFc4zq8Y+hTUloiBowNpbXBLcGyuI8MRloWJod5ShdJmBHvNi6d+RyIgqH
2RCe7UtxA3JjXKUx3/Ugp8qNh2sbc20melTwWxJP53FrpWAnlVpu/KOhG1m0BWzwV4JT2TlysAI4
HwjJwuXtQDzDIUwO7UeTjveWd/f4vJSVjC2+udIVAiQb+KjUCXabrPzeieUJOorzGdASHEWIwN2r
HLit6rge39AoU34zOpIM4qV+SvFA7KA49VDepi9XYfaWFbSXed/pRhRtcPFfg5GSCZEwP14QOJBM
n/u3u9ZE6xDOf61AheNTe4S7/nArLQcW7R1/9tlY4UzazGcTFFr4oLGUcW1rlgpIqdMqea4Xbee6
kNgFFOTkcOMeOXSYX59ygzjn0UfzGEiQW0DKpdBr8feTare067fPSvxy9BHstO5ahBrDWPtXMfj5
FBxmc0fk5CNhH2X6l5k+0aT4X9U/A2AcQmgXDvZCBopU1fv7OAIrYXtvhMHO9VW8Jo0v9oueh2YV
S7OtXp8F4SsuItBkf2q5nf9jvJKgTTzoKGB5hj1gU1cg36rZbdjjdmdW8HjyUw66B9FfNRkaOxUz
cjlRdK/03Y2FRVaLAwvC5ITp5PIr/8C0k/6DfiDoKBnlhP115GG3a1w8uOX+1RfAYCrqTcf5QsFf
MuF7IwtEBZooj14HgfDWEgaEsDL/LYjahtZ6VoUb5yRx0ZXxtfmDYX1sEMV/FSC7lS6uyjzvc4iC
S3PiHnojWO9QeUsVZCH/2je930RV8U7amwFVtNOX27XCCijxmC1a6u/+RiB/meJaSQB1lVsfRSdI
3DFIU2WzEON8SD3HfNSbM2tbXP+rIWBy2+TgyMmUr+JdD4B9EBJbPZfnj2Cf5I8TbJ5R+6sd7IQ8
YZ4UcE/vb0WHXl5zjSb1je1PnUF9OUK4PESylHecu/TSYTGrJLtpq8+f13XuHh9Jxv09ILAvtqrf
TcVTEdSy0qRld8BxBRFhnb3bZ5krSeT1Ik7N1fXZqwfp4LFN/c4SikgfGYLYz7N/4m4HcJn4QgsH
MGt2efGW67g5nTEUscQYZ0ii9DrLiBCCGyxhEIfQhVWGXgo6kUmJmGVCXoFIBcXdmr93aSOjtMFO
JGoGvsk3LZjEqNtkMuOIpyIJuc2FOcye7TUfJ1YqT3mOrWh2UwIXfpqwdpXfZgQF0GSn7zceQquO
qLGUdb/vXJJ/L7TEPNy+H3whvGQiaHCtxpNd/HZYRK6lGFPBl8l2dRPeEAyZxv7gvf9hE7IwS+Pn
bV3YH9b/IA/VALiZFML+Ftot9KkRiwNxr4O3nULkdyNvnVgPY+gRHhr7XN9n5t/+BPBl/+A4edDQ
iDlAe4seRgH7fN8h5I1McJxeisiolnGJLE4B4sIIKuoJfxk+NBkPr2aIOcEhk2CJDJqPH+NW6yvE
5cTZ6Nr2cBsLdtwK4tJD8gKmWriTo1HpOl7ZJOpEW9QfiWAKn1fCEN/cc6x2eSphAzEZHkuQaK1W
vTx3zChuU1VCLUsklTMje0uTU8R/mXdD07HzDSzPLuXNcLuE+BqXcZrlXUfO/cDwylb1Wvd+LCgw
3mWsYEAVlt40IfvhiJIne2Sz3Nz2+S7ER50lXyNTo8nx3L+bjIrVpli9p9k7+j/TS9/2JCCtRirc
Vs/t/ci41uQqLkCyY5a846PoGzUyY1miExMe6Jx0fy5hC4WTJANmV8WDh8aXVzX+ujOnKILM+WcE
UcUEcOqWzye627oKJKtlZyIJN51iboUjR0m8aGJpHDntzrGIcjGWDQ+wuVKBK4FlPwa962kvqHMq
EvZ04nkg8f7Fs1wD7ENSjLo/25HUcrDtp4h31mgXbDtxg4SPhkl/4DwaLZtGF1AV/hpbEjBRSdJN
ucT6zvyDxbKfdUqKQ2hevPOHIesuT25uTechqReOnG2qDFcLgaeYQXeaK2b1F4ERkal1h73HC6BM
12ol78SjSoQfEYvQmBY7kS5NIUiqSZwgpITtINkUPsDV4xFQwIqpFurhgtyMM4IctZeczSUUIUCm
ngB4hqpcLW45QknYxR5z7oMOlOZp7Wp4lV/4eobpllAnXzG157T/P5YzEP88LAcfZyaIomsKbDIO
TKFxqm9Q2ASAaqcMRxQxQ59xtv2IzjOVTlloT5uDQfHMShNqMXcr4c5hzj5QhFjOHydhrCzPxASK
aeLnUFl6V6sOAXq9Xsb2VP/GRUKxM4BO8/ypFGyG36yXckpLp9ENGzee+PQE7c46uz2bC+w6pHZc
gjj+gsCJr/VOByQURDL3FHhvGvvISa6GDfhLejFPSTrLVGl47yEc+b8zbedmLtVVAV+aMkfNmoEk
FE2kr8anuDxTYck/Etba/KRorjaR33iKROne24bItO0o/vAKYk3xOA+n3/9fkG/nzd6AhYbV/iw8
qquAUBwcoYkKF+AYqucBqzubWZNnk2kaPCYBB63HTEjyZA/p0hz7kyVDORmk/zXx5VuS2R5JpQTQ
iJ4HOAGOFB/LYHgEOhtx1XttocO5QLhnDhDaV6hJULZzMt1s7854kN5QkEL3y/L12MvJFwm8ETGv
H+BbY4lqNUW/HJKy1kcKXjp28qcFPs0Ud2KhD+gtW3/j0YPxMQoH2GweByEN319t6dXHClWkWW/m
l35EWG9l7u1RJzD94XIzW+jGVP+A/AqCxe/eYMDPXGphHPmK/5IWxtdwbzjmhtlx7rfRNpmLuDqZ
Mk4LXQ2mXM9iri0PAY2zPBUbhXt9VUUuEuvcVkhQ9DlaOIkM47K8akoCz5+gz+hy165yakPqbLXA
CHUSknMvBnts+Ix6p+JwvKjrLnvqobfDtJkAAg1zkfeCPCsrbx9DjzVTG7lC3WEuhMI1O7DyEt3S
ugemGg67AI/y7uhOAXPadvo3ctFgmDDEFTHpYDRsFMnRiN9K+Ctj8+4e2UkoJC+SLgSAOGvYaFF0
e0jahXL+6iT1yYeUQArARFShn2a5YaGPUms8uhQrnf9C3obPAxQus5/V8Gy8KjD48HI5RjN2s0nV
NJfMefW8tI5ZIDXUXt1mv7FXJtB9aUDGBRloj5JvvVW4zzh54rxjAK7oIK2kXLDnGbbs8XFoxdwC
tgVXAfXCqu65YmLQfN8J1XjqjmLTrAqJiYbUOFiBmsiae8jdyipKlWwUAMFDrIjPK46od3n7pb4C
T6XjkZK2jMGwH9c3Sq05a/X6PonEP9nMgtsdOglFiaWDA1z0wMefozz6Oa9R6/rj3Q7/OeE5F2VT
bot3+hhFzEfWzbnXg26mA+CNOD+n/ilFynd1r9+l+YljQe/vkg7CB0lTgCudykUw4pn5yVhAXlFf
EekC/6sfL/bJsjifAWy7cxZIEn8aoKkJSFv3/vkEWtv9s2IK1A4r0a94ShUTb+xZAlGZPF22LMXt
Hzmn8fkR7F/HXEuCYYG6OtkdNbAK4fNOT/RPHu66Idhb472euuGnu1Nm4AFRGMzQXibLOQ0/r4Bu
AuedjmFgSSpeszSRn0kYpyACj1NsmGkZ3P8Y1n80XzNUsp9USC38+QHR7WDeRG3K9bqnOud8+x5r
wCEioazPStMtZjONZskt1I90IQS83r0QOhSdPDCGTClS54X3akM0e/aLxEYcOEDAWG1HBiEGaZ8x
7on3gtocmlSFw0VzgnXb5oZqqmoj7p6xsTeKfi4IJV6sN1ar1CFmr9mVKhxomkWoZ2ITvUfH2tjS
qjw9LJTxwu//xQAQxI99xSVIxgbY0iGlA5QBrfLY8VN07m3snO0W3X+TqmWx3bCJSLapbCcrwTxC
Bz1nL4pbvZG471cGV9wC5B/9BdtQsOg7yOdhr3rSlB6h85FmknV52szl9bjZ4z5Yn1eakq24PCFc
Baqc3CJ1/qEjEhjzZR6qB2qSagC+DrUDNk6PfTrahFog8Mi2nuKnN4t36z9gimop6l2Ob2LjWDyO
wb+JT1hHuPOQA9aTE0hP91hLc+tE+NAeUeGtdEVcnc3M6935ZOTxxaUHn1k06aLGkg1aSDnkyB81
wG9JbPzBcwQcym0877vGwfco1dcwDIGgZKTVdmTcsP8hPPq58kced5Gz1WLR9g0mLBD/dImEjDsY
4u5ecmixpnPkEZIr/m6P5C+mwJ0R1IP7/vo/0L0hEJxw1fNfHmrj3Q2MZoJNenOG4x95TRPnoNu+
XAC2uGdcMIrcXmrfEPjV2mCOc+JoAFt6WkXIXD2vPk7BB7+/LZvqWYAQu2XQkfmDLOhcjtwk0Ygv
S+0CIu+A3o9trmsYUqkxPq9ZWeuqA5U9k4iNihhD4AA6oh7UfS7zftunYZTuSunolJkKqWyUYtMJ
2bEf2OjKjS8HJAgpDGSFtDP7CUDFC16Q3TXdH4Ps/w+jjkHG/zOctO7TFQMg0xHFrP34Q7Fs2k35
3refPJeSEVqst32n5RwD7mK6ydukVfDzvltwykIEmkgGlq95EZN2DlN0ec0ogijyLmkoJFQH6lmD
ZekxFiDr8VobQbn5hFc0tMh1z0cBvWMsWvT2tHEiGhkqM4PAd8kzl5ceHCiJ7WZar7Lno2+WoliM
xI4zuP4sJ+14Q66l+VoEgcLj6AXv9IxYCJj9TwnvKDXYKYMPub2UcaBJxu6CAFZWdcaSL1cw+QEe
YKs0W9DdR5HZ6Ch34bozzcMJXexcufSUBeElR3Tv/Yk22pZZvyr6P4Q0077cq0U5o4QIHYRlv0VU
P/5tdTJysMhHybb6wed+nxbZM2HVXDrnX3yVb0H9JxXm+joNZcq8rqnzyPrIY+ONiN34WmdaWwWv
UOi/LJ2RxbpuN8qhlEXTGU5tU1DNzho9fqbOc53XcPj/Hc785zY98oQQ0auJE7e5JO8eryny4KS7
CSDl7SCmMlAd2OEM5f4PL2ZhNv21TtnbxCa4DtFGgHs2ggng82pL/eOPomGZhjAnGRPD6lYMTyHb
5XVkaXeIK6V7YeasAUzwi00u9w3bulSLtO+d9yQkPbCGzyvCpf+VPcytfzYsu2Gtj42/+1XdToFY
VLzm1geHEpMMlwJKtTVzp8c6lsVtYXKomiZqrqJ3Cw8ND2BH+cS+1zXg2E7/+G0vuQUizH1xjdVs
AQUt5Tsuuo3NGc6c081+ExrPeXPS+YendZcRISngeiNbhOlg465HT0G4TysQzBf/fJ6U1uEFyAFh
FxykwUl93oy4HxHOBBWgI6dBAtZ7fovTFbKANgZXgpzT7ErRxGgkv62RbMXvgcVQhcoEQ77Pxhp9
m5nhad7NiMm1pdWx8pKTtD/z/j24P3NQfpcLkficGUNObDr4wyIE2KJkKWM/ypUZK00hy9eJ/78K
7RxPdqzPzXHIB/fC2LcLutso60XQfYvwvPiiz0QCGWULZPX2dZmNj0XcSNQ3Nwj6Q3lm80gUeGxs
VUNy/BUJm72a+7hsty3715bH9/XpKWl6f3pALCBI62gwuMTf1szruQUDmj6TulIrGFzEzf8CnBgY
gXDtiY5CcSOJXWvWbJOT9FXRJcBdIEfHi555tiNIrHXqIM3BlGwlGNQOHbi8bpgpzOp59g8QM0zd
I9PGbJcqy51tbqITdqaBysCZO7jDH4LKMZchl/1a0/6SG+O3aOyHc/uPpTJGEHk583ydZpsyI7x6
NnyJUnQNfTGlvG6fd32n8uuqcxW4sxbpm5gXy1m2XsWR6AnAEGeSdpjuULrlpULUVq4FEYtAdHv5
/sIRH4q5YwyIz7artrTQswEl8+QsrZFlZwOXxrmWKBTlOacLV1MONXXqGuxq3tY/UY4bgiUWEEqM
AbAOy+1R0UBX58mKSJkRnDHPo3ptStgABx1K+X6IgubP2o+6z3VRpOsyvlG0ptCTNx1BWQGWgHnO
U3Aro6VLBH3ZX1plsuUKDxgeVNMKO5aNo/8gkzAp7WwTaZ17znSiDhXjgFzWG41Ixka0Em+uh7OO
2d2mZT25UT1Ybt7vM703A66LZhmYiiNna8vlTcc3I1wvlI8xWygvia3jZtbh6Qu++AylM+JeG5QG
RekppvUctRS4kjvyqHGCFk+YA4pYY6Ezz++Ff+uo7rMGWG7PsVfGTYGMX64Q1TwrGkejV/RZn1h3
Qzq2ljSUStJeuC4ROajESsPMDOAT1vAp9YTm1SQdz50Pux4NCwpQf3DN6oaa0uoRo1BOIEStudwi
3u4WfEL0E/xIgZtOQxDGyMpOBz2363rZmfpeIv+fSqIcT998zNrybZD0YNao3WDYbNfcT/EMIU63
/y9UJlJLQDbDTsEzfkr1Cj5XuODdJsvhUohX2RyqUFJjiECkMXY+HlBXPJPTsESFSqG8hPJSRw/a
XOl6RQ2h+oobktvnZ8mv7usntNSAmFz6mThhLJytP4GSf8n8ArWlMjji5h95SZk18ItFIyMyUg9d
AeIZ/7z1aNqn38OrpBSVhJMwTmLtlh1Wxe0klgn9aXsg7FWxkFmz/PDKv2svls4XCOetZaHCLczG
SC99e0MClowpUDNXYMReoRk0xUZ1z119W/2G82PRIyJfpf6dinyjMoAbDcQXquGRsUm9YU4jevlG
LLM7wSncWetvjthA1fhsoPYuU0mu+hWrazMw2WeITqLeKF6DWnbqcHukBXFCSyetPCRZIzuuIuYi
EVNTBeHZfJXmMFKWIz1DWq68dKj91E4NvscRmbWa6bddzn+0WKLiv/afGBMKvUiVZ7VkZ3s5D3JH
2Z2Ku4EiSQ2Q4torNRtHFyShtI8kxRRPfeqjR6G2MYwUtZbNyn8+FDNb637GJFekmNJfDHav5so/
LwynNuxEiQK0diKJd/GnLi6FLHgdaGtBwI2WREUXEa7hXSjQfF3Ug2+V+K1efnVLHirVt/CfrqbO
5yU9Sk3ZTvbxwhAswI+d0yKFD8dkH2kev71Q20pgKfRFSVHThiOltobQDK1kHdpY75Yq1b1dBcQO
ZGHWv/uKPSk3v5RGhRsy7Jl93k7ucaUMhPqXm1yBQohhaV1OSzSP4E2+J9D0IEzHNd44aaqwntDd
wZz2y4MdSJ/gRn95kZ+gP4QEzN6gHfkxoBLW05ch0CIgcnNkYryHhvCcy0eAXZPaIyNzlPDUFD34
bQcSl8IxNE7eFGtuqud/iX/kb1JSBkP1WcbapuZrAZuBAKiJ+u7w9kwGr4tMKU65nB7BpIPEknfc
uaIYQUZjvgfR7M+EZigeUgEVM9ULR6qew1FKr5xRwyzBCWIFp6Et2lDCd7RL/Z3Htc6vHMcmp65z
8i8hb/8gCRb77nPcblDnkUTUL9DXnQMLZsCAYI9fFHXemzCVe/lgJfMm2SMj7GDelcsFwCmMSjiO
jMJ/0ROL5JvX0Jmu1HDIGEPxNxdGiXndJ1zyR14yeHlAEZ9r24sxqkJfzqlHidNyXxwUj2+HSa1A
aezD+yvAwQHuutOGhxdNEB4rMegdHvOucALEYIBawx2mFatVE1H90JERQ+ubRUw5Q4E4yih5NREM
Glxg/HjxkWb0e+duEUJaNWIPZR4klcmqQQ7clQX9ACKYXrNJ7U93/WfIlZVirABa3rdtrGWh+E8N
yyF6+ruEjFEo3lMOqO9lixzFI5+xjMMbC1ROPhAlBXCWdBUQYxKPhJU2KKWVMlAqdVzZn8AF8w6C
wLBgmO3kDClYCtWrTwlPhkRYZiv/jwawdKbUY85PIrq2oOOkVhSL+NXHVZNjbmWWc/cTfxdwKxz2
JEIobUrcE4HnBVTE6JJjqDlkv5JHC0pS/tgaqsZaYpg6nqSm3rC0vZ4tgwtlS9K2jDxbz+I3JWja
7CLW9ACByx3S1jNs4WX3m30a43AP+JNjFQWMiQ0esZuC2crOVSf64OBSlfJh6GX8NDP0dLxZ5f7V
BrS8IL1JzvrmJ0eYvfJeW+BforyA5zG0oQhU4EXzHuDeBkeB1nO+RnG2RnLrZqrV2/msF/LML9KZ
KfiirztPrGPaMezgZmx0NhYhllVMWIUcvdKObBSBFb0e2/YVYC2ieedyTDQ+sPWlLOOL/jKMX895
PH7smQnjyVXj/sg+FjhZgX8bFxdN2EITbyXN3xO0ZEwvU210FDakYLj/ZxLOHy5V+Plt6/IhOceY
/gfW33RI0zeeXdHzLu3IB1kJivd1oW0KNoGFt9dmsTwpk/+VfSK6EPv5FQ5yOnNoo4HG8AGip5hn
qXOimGcRlZvbQL1r3Usl+f2P8Da4g+5I9jsP1FP8Ikk8qNk3XVu3QnR4drsMd07b/9Odm91ZW2q5
qHfpKkugX71CcqJyIZvNzlKwVf3hvv9At6e/oWqNY0e9XhgWbR8x+APN1SotxZr02TxvCrsA4gvX
HNOUcCMvbR/oKUXTGzfKfL8xNTkHPGZpouOGvrpdhJOdl81Tx/PNg9u3Cq/pL4XFBHIVAhOGlFSF
NKr1d5kl3QU/3hWqOasOQTwTUXxpN3FiHQnN38KKeHrAjbmE5CQVR4Y+8AcYmRbCTKaSWnPzY2Bx
Zrk+Y4md+8GhUf6JujlZGarOjiHIhXBtxJV1mdF/FdqHbB+o/nUYQrEx+ELGPB6q+AuSWSsVwp61
dPP/Rnznq2h+9fS4Zu/OF4SaguwVZEWAjVbLZqZFzAUSQOZduJNS4kVFjNsSuFjvzlCr+WBxmAUW
GHg6hzgulDeMdCcdrLXJ1HBascY0BGRTKlRYE4nBLdchAQ9i+J+6fDxlaYf3pQZkkGIP3dR+qa+b
ayoiuizGiIwmtFM38AzUG8fXkLnOsYdr9sx8wcmAGw17rQhb293BHqP6VLMhrnbYAushmgPxf8gF
0mWpbid+E1KMo6tdtz7cS3nalCnrmneUO6Bx4D8v2BskhC5wLwS9QYN5fnscCz1b/OIWNacwBuwy
UbJZdV3eED/S/NWJuYcZqvBKwwxrT8+HgWlpSlQv2BP7f56P2/hv+UmRPCZtJTdSTUNxkHf4qYtB
ShTJnHzLB7BWiwoHYNYR3wL8g48UUYTIIZDxnY8uaMUQvlVzoBCHJ+P3l9TV4UgPqRsSpVDgKRRh
+RCG9yELSwsamaf1NOt7Q0vbDV/MxEXh7VncCYdrj5NehWK+8hCbtyxMWYcXmVuX8ESbH5PLiHsE
OGobhJyiOxGxKNYOgt0q2/wdLAVjM1tZPABrjkTYpXSy2pKLAlTsViLwHzOuBIs/WXts8iwziCl9
e4o/s7CaXX/OudEggZrcIZH4qk2h3yak3bQBca9IVgI3+b7pPFy5hEZ3IS2XBEYPThU0J/K+Dh53
laQ5xgcEUc/GwkND+camNDdQUwiahRKf5xGYhXaG4awm73XTQ7OuimMEMPHbEHxwiWmYZ4rASwaw
e6dVWpfbTa33LPtpsn14R7NUpIp+Rs7XKXbZEm9N5eTaCIuXVOR3gygq9lvYYZmsm7ZlgiXu/sT4
FXgddCUJnoVrcf7mYYPU7CYYYqxBKo9P/hg2PW2HPLntayGnCUgd22qj+GaoLaem0oqq55B9PBDo
jLSg03H22/HEimALlY/Or2U+MS2lOoiUhpTWHyw5g+umbqKoqtZRdyFi5ZmpHHKLmyv7/YekZqwF
67TCF0pW3Ao2eDZdaIwk5sO0NPnK/E0ORxL+1Kn3HcrfS04OL/+FPdY11BzanBJ7D018YJPSrQaN
alvzYS4EJdqoCHy4k8jgN7HOCp4CgUS49uU0oSHZaTbTXYvGcOu89Iqo9SAQlURYqfMzgPFjqXOi
7ifWBahFmpIE5/oM4liOoixHI9ttihAV1kZnFZg3jzf6Is1PIMqV6e2QoMsG4Frmm/T18AXdREkV
l/ViMFAT0JQRWy4l9GFz83UwXcBinrZuLRLvgTX9liTpZJz4UBxoycN1az0druRfwnCn4MBhH0Eh
LpnXYghYRopYLXWseNxSqzHWa+LpSbObyEBWrsqshmTftcuEM0/G+kV+kMJ6+dE5aokihlWmwnUa
m65zpOjZts7auCeGkj3yGl5y75wEtu1H+Z+RkwyCkSf16hj92OfeBkPVfYBWPxUogw9Yny1y19+v
jbalobDk9cXkMJoOutC190E9sGEbLEjZ3YR82jZ/puyp1RVQaJdNuRnSijU+t2OWNYk5hpEhJLmU
h3zu0VjpdPM2C7y6Sr8J8lW6gCcRQVqv3b0hSnouGmPY9Ye3ackgYyOuLFlKgy9PYxThRli8N7e5
E6+jM2xv5zJjnqvHZxfNlGbc51CY9sopc0O0FBenqN5TdfvTczeDSP/D6799UYyL5mqtnoVhqaJu
Ld8G16a94dVN2AE2IRVaH+d27E+R585B+Fd4wcq6TK0s9rFzI1Q+UGZZfdu9LbS79zEnAuIm29P4
FOyZe2Wv9MuOZvYmtNO1LwDebiX7PShu7nGVVLFiKjv9Ln8PvGNGTTwpjannNCnlz+5AFy7CU7xD
qRzulkfcFdeF1zZyTSySKxDBaOVVdodToJuWUOFAkplwHqF+QFIUJEDOQX071jKteBnAvZ7UKoJA
KE4C9m19KZdIl8UVzgTlWCQecYTUXyg6a+pt6zKrgpKKXcq3g63RoLxAG7E1gZZ+b0CX6R/w9mSY
RJc+EUWpgNCQ+cz9Hl8SttGaza9fluUV3TskRPm+lJnR8KyFPY/uE+o1G7GLCyoCJAS1xzClfZfb
/ZGdfCHw4vtd/erggFJumMbTCQuUQJEPEshK4NQOBA/rxdHYR4gFwr9eux2S1TyClgxztd8DrUat
YEWV5yd/0HYQWr1NLf6VuJ/s1+a9RDH3ilsb6OyLvcHK9YGl1NT6dvKpnAX+kXOAAQ0TxtKIVNup
GiUzdBJVKnMj/ycFV9eRHtP6EO7MfqYxfPImUCl6CUovMIIePO2+rBTAZ/VwKb+LcFtUSv49O3EF
6/w4bKnM2dyiaPW7F4phrgOJsYzTjdBPEjsnoYiGiFdYhsly3/NOsP/m4Dzu8iYbnLIGtfZSJE3B
otHDmNkgCwVX+iMQkiz8riqPXYZ/cVioI9c7OA4tRZFMm39V8CH2yE4cOUUESIPV7fV0TGB1qb/+
YY+oHR987H5x4HvT0opuy6Ay4IorUTZ1q1aEC0aK/7pr5XZv0hj9Q/jrcB5X66cislCSGOtLZrIU
bFCZpoQwcRs8ILb5050RwbNAZurH5Jpv6gBPgqAoS5JyvqisS0v6XulDBxPlF8lEvC2IoLZLhYPF
BCtxv1tctVAl5Vs1xt6oAy8yfMCz5dTEBHHRcoTixJ7ZPVZed7QnuvmPkKjlVbLgNm1NqqAnMc1d
Qej6xUusMs/XsWox/xzeBaw6t/EB36Uf4D1dLp3lKPMHv+iWRNZgL2mPJB7XuQHSVBaL1TLR5wK+
8859td9FkHHWxXpXbOjNXDaRAcDyLceK1SLTLsHfEnb32R5TJfUCYXVkJPnjOTrXv8lRLMsW8A//
RfEQOaJRJtUau7kt7v3a6i+1C3C0Lw7rLN/3Vm62cR9MWxAhpEJtxgZANlO7qBncjJDkPqUlxTY1
MOOvOQxyi0cScRcSGg4zT5szgcMV8sLHYcPy151ALvVAHigBpriG3zgnY/yYknLhG4VPA0zohyjn
QHsA/4E+HV2b1utn1WsVeRK59rYrm5QgJQvFm6zq4C+R0aXQBTZ+wGx9D78HEAipBvZXwQ68br1N
7EnyfwD3fKgYhSX+bTqUhcLWU5h3Cyx05AmqRXCqejvzeSsc4VtfjMcuGh2WA3bswf4u2SzkBcUk
0McLS51G/FUnnfAqZO1y/oStJRnuc9bRcHakGckpan0R4rcC8A7myhBKK1+BhvX2a0eUjqHac9aW
jQCNfWNnIJ/E61z5nShJO4rUgfW59xMRdo5lyMwper/rW/eCTs4liZhCxTSsQ55RkHSlA+V9Wmeq
wYfkyAL/HvZcgVaK3usdY8Ug/GimtR7DRJPGsdWKfGh2R7HNPeGG9Hg/jd+P9QkgJjyDPZiQnIcZ
Pk0eAF2zcXQya1/mhVmIPyzYLibOApWsdEug/xe8gPG/4kI3+M2NCs+3MPWSChLOq+23789v4DKe
1E/73pmcNqJ5yBiFY5UA11PgNsGvcLNCIpTCWvq/77ikK3A+6gKSs46HPLys4AmoM/GyuU6A/kjA
XnWVaieOEYJCeVkZ3P/3ziKuNMkqm9+XkMboWEv6NtxlPEGsanuQNAJUgka1B/2IHW3mPFrtyLC3
qqAdctF2dD8OwBULYOEnq6CAvA3N6IaWxsQOO5axMlYUH7Tm9pCSkmXBkn42fmg8bumoXAp1OUO5
SePadHwDKTbUKYax1d2H+aWoengv5eZn2KLoKRNcJZopSxM08dBEBisBrGXPnih+JP3JbbKUmn2W
Ku8P6D5wbprcMNBvalBn4cmav9lXkLyxSw1d7Cysudr4gMyBK8Rz7xAUrE8Oir9lagNGRp9rnBcr
rueHj0or5tA7nlgyqXhRg3NvzLO4Pdz8AyKBMpQNbL1c23XlwbZ/fpTM4YvtGPOdSoEt/s1AJKte
4yWAyiGAaZvP36DrKMSnsd8T/Y1aLyU/W1Ovwsy58pJvzyx+m+B2mMlQZAW3S1hUStwXuZ09jNQP
yeT3nBJsOHMorIAB5C1aqw0UULsFuw7woJQNzlo11b3ZVXbTk+Bo7f2FRu+Kf0wBcwlRJ74g3vWp
B4QHDVRG/NiYZsYWx/lAqGRBfPupVsq4SPCHbA0IuwVHBCHtaC0NkqBFD+OlVHhEtqS8Z8LmjQos
WA4lKQqYFMwyAW6QynnCscmruYDimYl2Aiv7tW2AK8vOWHVyxOhdld25eDr65624x34xP6/x6q5z
zEj85fBtgjSynj16Dw43Ajh+UzYeWb3jtBxUsi6T8hjWA1otZH8WsNVPK/Do6BqJA8HOmxOJZDb/
7v7tk4V4vyN/ibCiuAvQmZUFc0MJod3fBT7T44cR1HpPLoa0u8Y6wKy2JMjxHqXX0ny9GTATe84H
XUJO5DOkBUP4qZkTTKmB/5+qbcM8fkVZpLRenMeNATyxkqdBlJ6cLA9a9yzgiNWOY7oCxrlVMtVm
S3kBgkE/U6+fn6TQbDjGGljEYENbQ2QVEKDeJxqckFslmHsneitf1fSSXo25VFaPaqSEhtzuH4w7
zdHstiyhLZN3yeqgHXKCir25mfwtdbq+y4CcEkY/W6u/Kwzq1Z5YGECpAy0GqGsSv3oviuDIQ61C
goJGlQlKJbv7fzqdcIWTA12a46tLJArLt1T/PbW18Y+05e+ByJfgb6MLzvM4VSYR+ydmvN1KFXJX
vajvUFCIreQJ3it+9Bla4pkd/W1fCP02wwN6Gy4SdRk2WQLCZraxCrWUDDqsS3+3lRJa68qEz8tm
06XPFsZVUB7S4Rgk389dlICzbR7t0diJBrrwCYYclJ06iRMZ/5IBPnqQJ0pRU03oMUIMhD2fKmwE
3+tMiXF9sjtvhWWA2S04OIpmsiXWgfQz3ldkIbgnaDMLqNJuL2IbdVXxtLuM0mdBLC3Pz/kTdXU+
7W7+noMzEiqClFp3qAbr9KQZPmkxJuUsIpbUwOEGQ04N2RyxYO7dZI8Rip9mNLwK5QXBNYSfTgT3
I8YQM/bOUm4sVYlWNr7cDWC/3RPxk62IGMAzY6UlFoJyobYyqDVaQD/CEpWixkYqw05Mm/1DRg5L
S4+QOcWlONFygrbUBu1B1oXi8f8TW5TZmghJr639jclqJWO3XetZq+lCva2X0fqWcuT3gl8heUNl
uViiAdRDAqKwGXavsVl9/J6kpSlz9pbK+/q/AaiPY0h7EHJ0IM5i1r85VcC3seK/m6nYCoquGbR0
dj8iwg0Ki1Het7KRU9ss+DidTecfe1auzoNAVpAcMwFvBeGS0OOboUQMLqqqnifClQZliKTKHCfM
tmtvws4aGSmp8qBM5+zK5l68D20fqRbWc31L0NriNTSYwyaU6wzd2lTp92WL2+kIacUpy+zogZj7
jDVr2WDUODCgthIt3wncmi40/Qb6MnwAuuLsqEz+WxaLB7kE0d5JCrXUhGLFpmen9D/tddy82dqi
xV5rVXVA60TVxK81FvsWHWSsPvr4jHo+wrbA4pvoh7173LAynYE/6ug5olNvvZPhdVYK7sH/9sJM
eM6Nw0hHjxWTKlwCA+ALZwa2TKYnTkuxnf5QcbOJQt3rUTyuy/uTbh4et6NgBou/iEiw/ECBdHRV
KYWPTwKthd+yPyGgp9oX1t9g4xSSLcTE+Cfmbc9/ZyBmO0QJNXy1g3su7xb54oyYL8hHAE+DEJKT
JUf6t/Pk7dfeuT+St27D2WZ7AgSj3JbIqmEJkbmtWDaonY7sMRBXX14BUJGdNCTsC0BU1varAUuP
4Qs50/fLX9tGCIVtnspLpzfO21O8Nh+FLbKhVe2IGDz+9ACengmdnBcKu7B/A+M/ZDfAi5s8sDQs
8vX4OJBEzCrTVNRPctHO77LyVPaN2brQGmxMaf/ZjqbXOFXPVVxCmbVFwa7ekkBfOB3UYXSUTHnu
st9ntQtoL09bdAkk5zf99TIDE05rPNoH62VXdhjn9+D+hHVUIA1UpsL2wUFdRVqJmb4M3TCvISY8
+jOwEChyR5XFs+57T+Ww5XCtXyenzi/mrZbSz496cQdGbnbSBmZUta3n6wUaFBP/o7NjSbSdNE4d
mkOkMdM56CfE/VI8aBZuhX8NBskwXBh4DoEhP3PSfbIBJX8Hu8f40LZPY9m+AvZo+YX6S1t1iECa
kuOrtHeDDaM8O/Nuarjc4CsHXU1/DifQlYSuQJ7zRBP7BetMaDSANcXF6iX61vwfbWRoT2ZfPrti
cUJi3fYeseGAvnXHa8Vccp146uXTVq+NeYRAuytObN0JEggmVQlA68j7pFPyRYl4MtfARhPHarCj
KK8RZV6iNZ/5nxweYkfGjd8G4Rlh1YA6VcqDO3ICT7NMpVebVw15aghO9H3f172BMptwQPxt1lZ+
bv9LWvlXxHG3yc3ZTv2tHbrEQ7FXhZXNt0vN70GyyiQcewyOr0lScBlXohnZjo5HbmLoywObL55C
XYEHlAI7gHhiB4r98epvF/595a/juESxsTyuZsozeQkckk73ED6P1WzRiZ2J/k2moD3WP9CAJalo
ZnZq8hOx+yTVu5CKJCTytJXZn+0wbhIg209sFtctQHMoXF8tdYhpIkaSy5v7dF7b9oyTUUxD09W7
qpLD57ZMZBo7phIsrMYg7IkGzLkiAi2ejOHZ+jvGFj0OV2p2Udj6WZ/OzEkSHQa445aWBsuKvtYK
QpiLuioqvFEjFCSszQbibNiAcbUIW1aL4gcb/wuGSksv3zOfwSm08oQP5H8uGLtkQhVMXqaHFnfG
n4dbIlVt+97cDNwSlmkETXOe78mmX24H0tEX/BSx6gHTFMX+UjZClrxn8SPqQXD6m7Cv0x0RsYIQ
4Kul287Uoaq/P49Ol/8/6n2iQlEjQGO19v3CB1IuKGVpSliqZYizpViM3qekybTEFtJRewIDZzWO
HlvPydWWdt+IWp57WyO0tvL5nEHG2pqMrXnZHyLpW3hXtJzlB0BnZdO/hGoZq7MQJe4qzgmgrn0d
BnywPeTzWQoHtY1/DxsSq3GJB2oU5zHKYOB18DoBM2jeqibjU6N0zQ17W1NVOYpCRamy7TGpR6qP
Y7JQb6a5G3cIzjWndNy5HNC9qE78WVkMNm2VQRj3BvfPX6Vsz5Ir/DsPQFRqyEanSxqWrRW8oYNX
i7UZPFe4bZY6432wlxQLqr+I6cbqeMY7sPn//CHNZyXvH01Is4fl1jlNEuABVWR4fibsG1EM4OpA
F3n5KElofYpjn+sofqeDu/rp/vOcXBcBCpHX1brj+Gn1RoimIjMxgQnFlkoFwAdAquDKJ0DFUowO
XgrNwLPA/U/XF6ZMjhx5WtD+CBMTP6JD+F/MnEGv/oFVXMxe3j+HWEcwu2J3OAD09YGQliQuZmjI
BNzZLjEd7i92RxVvT+l755Nh8hXnS0gDhBFUT7EOIxROkeJOjfqacsw6i03+pEHM96oXefBkQxDr
urPCACZWg+8yyvgX6/jg08K9mNZjD+g9gByiorSA6PiGnNLr6tLC5ynb7y+O60BKRn3QNVk8XI0J
0i+j0Gs/DcpUdoTKp1ANItAe1bMhNjohLjti9zIS1hpCZDhtNXiuusTyiJcnvaSs0hlADzr7yswd
bNuDrBBZKOWlrdY5atDQBez07Ofoe4FxOnhLE6t2KGggSMwfrefN45TPMAI4F46mi+Hx1fTtk1gX
wbKQCGr5jV1O6hf3jVUcscSmmHuCqCP3D6P0ueox8CuPbxL2YAXDTCty1ZKPFoKGbQrvqwox6MZi
Rvh46hs4I4Ejdql2iQaxNeVjpm44lnowIm3dn2WcS4Fs0jiD+WW+eE3jeoGVqpMmGRCPGInuhy9n
CSQfDE+lKVY2I0CtYNdAgQj8jZ624jn/6d6HHJL11Xa9nBovPlM0dCY84f+uXNJnjsAOVidCQNYz
CUaTfDZdO8bCn0dcVUju2ojSEUVNkVo+aBwtXe3Ro/tpNKuTA7FS+0L/6Aas5+yp3w539nLVBvC8
cGjoAFsDeYxPAk8ntSn5G5IhtvxzPaLZPORCOwEh/zM31/J8kRv3kZSLF2wKmpHy2Xev4Lh2uc7z
h/moOzfhh43ylf99vhAiGTO/beIz9t4L2kUTqL9tjMcmTGgsllO0dKu+yQhcuf0jLLYc7AC8+wqf
OsgryyI4aSTQ8kL8+UpuUV5y6vp54FCeNwjLklMDrRiYE4wpY1bQf9O8EI5Jq7gm/VZpTgsMVZt2
n46EadtqIcIBfqCDCOSQg1faShj/D0WWJx+W9B8QHggk48xqvA5EJ5GACIB6vGJ2b1+HsRjUHP6T
R0+t7xW+l2DjBhZgj8Mz17WO33HGfigvO1po2KrP75jnwVdvDPjsuSJRAC3aaNpg9l6l0UbesLLd
98rDM2YH2PQuowKV40DuqCc67k3uU23AgKn6WFtpTuabjeh+IhAqcTErKWPzNp/Ece+Fjf4cBukY
OzIJbYYBw/Ugb/DBoHmPnTg3qrLe9WhulM9nPGP+jJ2Qqowc/JOn/kA2HgPFH9WY0RVa/70cW/vx
b0BSrGYkMeCcH5xEhcx7Ushn3Haoy90yEvs1jMTYBdiEu1kv+b+i+qVIioA9gZaLz2cOe3yi+3Wh
e1cVLj+H0loQnT/83iaY3LQnamIv4ZIROVScCy4OD811UMSqVEMez3APJYWwZqk/m09iZDBa2Khq
KrWdJSeWYM0KcHgRT2CeP8Idjt6D8tXWC6OQyWvLVH4xpJxTBO/EGTjaNCmIGbqD8A7Z23zqsTTh
ZD38psYhbw1SlrNL5utHrbsrjisdmQHE3Dfk2sCYJ6X4ElRmlwOfZRYosPNMFLXpXwKBGl6DzQ4g
qlL6hFmzpf5LsozNGhNpG1k9YvN7Ej3lrwefI4pAkGLqt0CmbtUdZoyl/Stl9uRaJ6kYJ5VqtLeB
8muiQCi99eIO1uTjYrjBZI2LNUFB6eyb9FPg4zGlMAyq76Z6KOe5w2LMqErgCzaDxSFtqhGWd36e
pGArPHP+U1C0c/27x46TL1ZhPtIPvFx3eFUkVcBcH+PnywHtNExW7xBB2k89HcYLIvXYtkDncZxw
XVF6lXnI7v0dzZFKk1iK5fCEuiinSkpktVqvuhe+eV3YVz55NOtmdyoMvHWVpLb94BGZdLv+ETp2
XQbtSxZK9XIosk3QTifnonipk3xwUyq75rmSB4ep5gHuPDkgGaWZLDgT+P5/+Gws3WkFxeDKBBTc
Lnex7VhVKGQxn9vQZ7C9T9zF1NJox4Mxs3E3pqxoydgpJWOYeGjcobAe2z1Tu5RDYTYpmDv9ixmE
Q72ZcU/9ufhjjFDo8gWeLbc0rNV6r1p0BxjgyCFhuBZ+z20kd33Yf0wSzpuiZyQ9zRLMzeX1QS13
sy52+8AA6pxMyrCAgCPiZ5Uq9/8QkL93jpZy5KklQBUiXNgDUMKe0DnZYVZ2FMjkQaLltCFhSedO
76vnAr5j21UIauZwjVOkFJDwnNlzMTbnelFP58N99CqeEhJLWG1esApAkAzJ9N0S7QtL8oh8S5oQ
dBZL563TwAwd/kaoAFXplv2kQLjunJKaIE29Knyz95/MSInXc1cRyiEvFsDD7zT41I0UqFGZfme8
RcDmyx/EWYfYNebzv0yWjQ2RMddbrA04PeeCKA8bIMME2fq96jcN83NfThVKrcrfjWrzx1jtypnF
PKBdVyvW8Q5WbSxl+k43Fnxvjnq3+fatjc4RjbNf7+eCGeoB6cRLFw90v2okejop3y59Cj90DgNX
1CHlObSRzmKiTgUfFx7S7MuVj+fg9OSlWqhsOB3vwA8WtWsRFbI7s3nijIIqWPtiSXodj3OdoUih
fIjDwEf7WJUN/wjJBsUKQ7EKYwyEfzzeObqMG6jmQuAOLnxnCU8GPz92Ure2smrFEDU3m8QvftZ8
1jGzXtGOWvhYRzO5fjDkxeSlbPUs4uJa+jyxQ8aa/RXJJtPrjW2+KtEGT+4ltnTMXxWFDDKQyORD
Nv6PXj6lQ1FQTY8UNa+Qtm+JWsyXcKtMGTo1mpCUW5JhxoUW+qTQOB10IqbCLyMAz3aOoGabZtCr
eJB0XLA/nCDWqz+9RZAXe0CEMfFrFU1u8bJQHI7/kySytYunCLE3q2Z6udaD6qEqdtTUHc5NJj+e
z5QxfzfWCLjLSVPQVYdm9SaCcQs0EoYf6+n5bb8rd0PnS7E9RcLkUvM3arP5H6x734GxIE+Q+0f7
xc72YcuIdkcmsqVDP2Yt8xxFdOyh4jep5GguHw2czklZa4+D4wMieBr2hGLTUz9WZwVORFTJzEnW
42hNjacZz7pxbt8UrRNiVTmJckg7dWtIEW71o9Khn9NPtBcZeVxZthZ3vRVd9d/JjhoJnm0MTkqI
zmYciFt1Ji2eubpHFSFv//qJvanYFt9AcSZu5fquXL76AW/g6o3bCzK6nLWgBnpC49M8igaoPHEp
ktzpQwB7it4R14iQ2/jwm6khB77f8BfWBcGz/xfbAiOsa27EQ668gpXhZ+rmt2KwskdNgUrBTpMh
2yq+4+SJk0kHfAc7aonaT/OgP1tAKaucQsjZeqhmTAv1EZKzwsfkdxnWKz3xslZ9c8nGu+MKU4c8
uatCxOfSZcdW79eWj7G2VG4f/a6Ki8OPdHjVLyFr4kKFJx3cX4JB9qR0252ZOsEjdbWkI2oGOI53
z2mTvtOsndQnumLpYyR9eVDbz2aJXAHdI+EhX0PR/15ZcJ0iNtc+WQ/mrxAIA2cs819sgt2/goEF
L9hT5JrCDuBqDFehruMdSXVOl3RGLCwVPLSY8Vqs6b0PeOm8Nfr+BBd0bbvwzVr6omtyVyqZvJaO
JZcY0k/W/q3BpFGn3NPcc9rscrj3gNVBLvpqVPLJ/K0vLEKhHoJLvjbvdb/JlFL1+o4OtAH6adru
ISUd+vGb9tz4VYGRshWiM8l28+1fMN4bLEyG8RRTL5Lgn4rTrUYsj2GgB4hpuY69olqNFh8FNjRM
Y2V6jzSSgIQj5yonp+A004X9jmzQeK6G7D9FKrbxtmvF9Ki4MQ7ttVjQgNu+LnCAGQWM/jSb+UWb
u4aFL+GpgdHDqC0yxnYcxeK7/dWaeJvN06o3o+gt2F/ZiZPnU7HXRxeOBVQfb1VUJvqwVBhqtgSu
KYIZxNicumUX9gAh9Uv8pjzml35Gp3N6BEfZm7YF4XrgHj53140kxEFrGhFdgUBzJOGUIAgnS88y
AmCQSsqVel2gxMUaWiC2F95sVhU7a+CE6tsshWUqk2XtlUQ5uuCS4scgvVr/pfu0DDGVLbIbPsfT
DPd7RcSgD1I426Zp0IBsgQ/iXcTpOD04Xu5LbadBxZfmyXLPWZMtxkj3R9/Nw8xd+uzY6aZV4kYw
sctPkUAMq8wr11J0uOlnYa1bovuw9TXTbd/xJ1vC0aABFqwKlu3RIRayzMpZqPhwjs+yFsvsKySa
RA70V/FMuQR/rBsne7GsWw41gub9jxyLgZWFVBQt4Xye/FhzaAitCk+T6du0NdzIBh1EQ+NLJ/Qn
mXfKWo4e0sIrKzRus6k6qmAjM4lLpVPxF7EF62+0It5HgX0MdKu6P/Qm+fIm+8ahd28WB+0wZfa0
R0uyQZQzmkg2b4LTqYTeHAzoVqpANh0JXE25nu4y/vxDtmMczWiZZ5y3SiA0laEtv7tRQSVe326w
RiRnnuoidk/a6LCv4Vy2Lm4FL2J3J8k2hMYatT9aC1KqZOLeHyaY8VvZZKJCBBD+FziABsQNu6jS
IOCPTyKJ1WW78HW7pokHAEWGYgSqbJWzEzsTrxcYTp5nmH85vEwqQFcgsBBGieVW/PmR9Q7gTMxi
GdFX84bDkZceCX4qir/tCl1e5eEPmfhih45kbmggU3KcPOtNHhIeoq+6c59t4Bm6yTkCNJUODgfj
jSVjcI3a+jGxerAgabkb84nOUN3jLWR14RZf1PTaxbW07PpsvzKrYgasTQcTEzur1RHboLFclccf
CF46llHEJ7tQkElhSIor+DSB2peWDpO0g6z4vNHj7PiPTdX5p3sPxbo16ITueNWVz5KepSNT+JRx
MxIFMTm/zS5hatwtEZUtJb//G06c/sORnX153r13ju9SY1qE4LBteLrTL24T9+Q1uRM1yKfnNRvr
mCbVFtBfdRHsCZMeM18+Nlg2B2QIY73Iwaimgl1XKreO/Js/yRn2owdMP8cFoUViFeIfRT8b5I/U
SbgYyXy/2AsfFjNcamMq+iZTtAuXyE4welCDM/zHEdEHFg05x6nNTndh36+QlGFq2BMvedkWsLrn
ULvckypoH8/gsSGszzOcj/RimjqS5iyZF94Dh31JFkFFSEp0CcIFWmqnqrKUJTZTTEW5Getx3BFN
SWcPbw2mfyv+7vStpzsf+iRL5Ihbhfo0W5iVs7o3P3p1QPv8oDqXOSjW4IUW5zjVlfUpJzuK3HPO
E52+kgIxN/7OhOSoHKAnipQkSCGEm7r91RcguJ5YnL66G9O8tETda6Vn0euV8zRxoZwMlEP5rojs
RX22JFnckWbOEI/OQToladI3MnzTaLF04gXf0SgapnkMXfWULTSDSs/oykIbLE9jTbsXvnmzauu8
0NfiqYbIFA67BcaSJqYNLTgiKno6lsAp/FkDx2uir0J8/tcayLIMbZ1xaBehq3r0ObDC6FkQHwXs
8L5sW5mzgt9RqBwpX4x8Zaw9s+uWJhjQcq7X2bjZz+w13eRoJmpC9LK6ZwxdOO4CVBoidvOtNPXU
CDVl+z7qc4JSnCyYPJ3Y8hotopOP9Bk693/aFugnsiFyLT3DBjPosDCLZQMDYwL4E9cVhUPsQwSP
TBwSEgMJWVSlbeUTnU+t/DX01J84nfnESa4M/p0J0tcrV4qa+wW4n8zBTYByTIeOI/CTBIiBWjqa
ugq4bjncG8wxO0x2t35w3Ikob7nWmxJGwtCjLcW7sv0VkiAIYXGxYW7MAhYJyjO8ivjqA2L2Di6Z
8avswQPSCjkz1w/lS4+0Zo9HQfuLdFJ8L4sCmOgwZ82fveF+DNCBnel4vhyhL5+UIjBIY99yc24E
hr6hOFNGSknKSvGFqxiznEmO857nkEBca5j+38ABMHSkvDhLZDCYlsXMXiGJ6Hq/0FQFY3HTbhP9
TRjSAzj5ecOeFPBwrQMVuD2UCifQ80he3aFg4CH/ocIkcnAISUQl3ZS4ctwqIHKOsODEorGMCOzN
AHiWqmjWfyea9bLmAe430UeJ8BSoKWFhESLjCGFjzqgC7GURNNaVFW2uWWLvu7NVIp8DRS9IuzGx
agW1bebl+iHgEVPQA4Q/tNEeppAMlwbTGdoMx6Kr/krbVI1vGt0rQ5eqYO7m0Ir7bq0R3cxd7L/J
7Bs7wyNO9BtFSftzxji6T2XwHxscTstuajdiNOS6p9jmv2IcoSk10vofKNK8BmOrL5kLN6tM4y+g
RhE90hWmJCogpIYPz6ru6HNcp9lb/FzUheeE8K//gGQfbpwBsxSCcIlP4wcIe66AwugPGnZ64r7h
xrC3wjI3GYG5Ky8AY5Dp8NUMng+fLAB0AIx3K+tFDILBNLj/xRmGGNVG53iMAnTzMyvQi+DV1D2G
VjjF5eraDGuIlilRdQO/fwPN+z7yr+AaEdt6WdVZjkjB4TLCNT9QI2EoyHfW+X1s0Nxibq6pnj3A
NZ0ku4emsVQ/b5gWM0vjKQs2rxoLBp0VWEbcbBzBwfflj3SckY460z2ZikvHgNaGjKD9o210hp4G
yp0HbwqfvyFrwWYBi53xycgtFBAg7Kc/qmiv7mjVoedXVSsJQ3KGULnR+/1GHM8dHSalinh00f2B
VNCjWoHtnvPhdsqncnxrT2gkbLCVLl6ocELtyHXw+WwezIiB5O0ak/UOvxlK25iSdkLclStsBvWa
QOZzuWVi59BvD6KpPgdy/bVvSJr7q28YZ18xQsKMt1nptJExDEhbvuNtqAkZxPvbs16tuyAuGrTD
xAZkzmKQGdFE26B3I1o5oZO/Y/d9StRavYuWkdrM1gvkNTUDWuF85F8eBqSpYrsPhdImfX49X71a
9s+u0D/JWMmiDp9i9zopZ4JMRV71RbfKUHMPhbmT0j9PQqXpe+OrWo4aKg/45G9Z9EKuCN4B5Jk5
Dmj98R7ZnQkv39kflheKm8dlwDQrEjefY17xcDW+Ei1SBFClidWVzhK2CenoYmyUJiuidDTbMT+A
60q5Igx9R2hvT+irUK5kgZHsZqHMTisb/ZbiZG9Q66I74kZFyV2DVd7LJPYQae9aFeUANEjn7EK+
Fnw2o6I1jKMYFRTtMbEhnkScx1DbLHIa+/v7JkzHiG1tD/oOYpJBq0XiL7VNzqsjNx3VlSiPj9x2
wOf6ngOEYo8oft2Bw45r/c8grt6s1UO2scGra4eFlRXObh4juKPNjyGaGLCF4yaqO6MojeYR8G0m
3eL8yihrwfiW+RpHj6JFLee0d7WY3IEElXjgQL/R/k/Jd7fpW+UwvWpeCpHdZdmRIDxKQk6ZGOaB
3j6lXqRJ7UT0PjqZh+bhIORXuV/2CV479z525iYk/nLpbh4j66pr4bF0wKGdORb1uisXy6go8/Jn
/bxiluuDeKh6kdeJvdRSYYi8Km0Nnslhmyyvs4aIP9eSUdwjOyFZly9D16aloRnDmM6D73SKZZj+
ks+d7LrbEyQJ8yjrcO7mdFNEwsjgkH35h5OAZJphSHsFmoC6A4K92jKac9BYHeXIO4x0sI5OwZGb
TWIh6dt3nlRTcLJb2Lqg9DpHR9hf95qDXh7fvZd9H21vaSvMamU0KFU6xdmInVTot8FL6lNdQId6
nIpZGut1J6arepSIDU/atqu22ZSesWARSbksiu0v/6Q/bJP/owg4I39gfHO0SyWROUugwA9RIVhM
liGaCZfZmjLBLTo6SuZevU/TMG0NMhaPkBtd0HiPHPw6bRW2NuVS6ZlzE8tuMS6VGz8b0/RmlS3O
Ic0e/6fDYOcqg/X3ZYD/k/ib0pWFdrHKIutqvP5s20ueKJuTGJssCZDWc4xsNa5nD+ezW2pHYLkO
3uf2/scZUamk0DoG+CfyLx6agh9nB4kOdO2OzzMGgXK8fLBKAOLlPF54fjH+4H7siE4qmDxNAYOG
NTKg6SjxemTkhRbZ2vPxrD9p78NmOeyEd6BaHHS3LMWSiXaL1HTyIaSYwC+at6w18Rf6+s4tJJNq
FGLXSkfd3o0BqhxZocM4TG2ptiqRXWSQeaLHB/cNVQzI6Kh+cIaRJXIMnTyesNfni5FYu1333hmf
zO32LiI1rj/gx4qpEE79iTGUDEu9g8YL/N7jPrMUiMy30Tx2o3fDv+9wE9QtWVkfo8XJj9RBZSZ+
HIimd9fRj+ZSHW771OEcwNlx9ItQ4yeCkT1uQxSTq5AY8VKpTecKmh7zMbwhuUcgRxdeo/SXnAo5
EIm35ABlFZ94Mn/8ctGTpmOZS6ZcEgFYFyim8TdIYE6HhLB2C+j+FC7RbuJqbr+vrGsUDduGi8/h
8M+G1xa9a94lK1Ex6n4jcnnDxTALxZGqZgVjbAEv+XnTCTV4FLIsyr0Am2UUBrI3nr93W0T1jabH
qAPm27WPV3vyJVQukoNpH6qROJq59bl6GTVF9ZFdg1prnDDqxlOveYyLz/ikfeOgGpapMGkKZEI2
4yel74nk8CftYuTr/HrocFtzJssNGMbZpgSfSfd+qzDPRLAkLfZww8+yQ7XdbG+dLebrCKbS74zP
dltNdM1bh2v32DWLKBNK/ELPl0HlkMdz8vLe11BG3ZIcgfc7GFos4NYEf9JvH7wKbIJ268MLWFly
9LNMqrJddqymNAkP0cekl/oSokoBF97DBoS4OMeMNXUVeQUqt59hhn5YvYkkj5VsEZt6ooQVUZNI
lhuukXiQNIMSLVfrDT9RGxAROgHemhpo04oqjNVdO7nHElJooCGe1DpIbxYjNjCDtxx1KUNBIAoN
jkSaNV5u3qRFAdeYX+R0X716zVgD/35yKzYDuMLo0WbXBG1+W/1811cp9OqibQbh2ZMIsRSpRUUX
xNpl6T6nHoJGk6O07w6OO4CpD/X/vWLdmpH5CuoY3VEUTkqeIqGndGqHGpPidXUkdWGuDe74BtnE
CbPuuHyLy7Xd9HD/AAmE4gV2OVxU/c7EgMiZpDiJ69M8P0PaWMUo/bkBmhUMbNIgjs8aU8kxS6NW
bL0i/odq5k+1tcPNj5+/jEZ/DWCT+kMolbcC4IdEN0I5P6tQMP/DD9hTGsKPeor8TGbs89OBGu6J
sPEQ+aTdtaJyov9S2BaxUqp0AURXD+iYiS6QsdIUExFj3bh3o2CllvV0/zh0zxSzvVv3WAQYE6Jl
ejhLgNgKmgkPFV801H8XpscnsQdQpGIdVS9xVJBngYPToROVjRyJzF2o51RZVI77JfjVNn2VO905
aitez4WwOvDaH0b1uV0W1iWr17JW0p99gGZptJhQesTbWoqBf/Qo/hlJ/qOKGeUQ1ABXGcmKpEbg
nYUhmB0tsHsG0g4p7wW4uE9HR84GHEbaRz5m9LD5Y23vFLDCB0gA+rhxea3ZC6L+0gyATUhU+Bk8
83aS0jEaIz/FFHuVZZIY2h423Cao4JrXSlFGeI9FStY6SxsOLLKY7XZd+5+Fzrv3SrylrdX/x3vv
Em5WguC0YHCfKhdhdH/vf89tpcqRejn0guz/arDQrEn1PjRYQSDmy6pHjwHFLldSOCj+8z+aDf5a
7Rudme5INpnsbq3fzzwAIPPcrewpOK8CcclCHRuq+Et6/4330r7JaebdRsBTnJQ+nf1/xZQPt7Vy
QthAunhCVdPN2veWOHYWwqXcwWaaJIqE5evXL2j3bVRNuKTx8umlIIKbypric4ynh5PZofa1LhGX
dcyr2TEpMx3llCiT5sh+/32Jy4UCSXDL8xHT/ZnroCyD6SDuJB3h41uV5V6F0XsxOiQJsel6bWh/
HQxrZCWvvJ+OmYdSzKRtsK8+ZSJCTgQMLyhKuJwgiMDGnq1BVp7j0SfmVxXMtLFlDAbuk4EB6X96
yFuhTNezUtnXyeilng6woORmEHbr5h21g5IuUFJw4PG7mT39ZFRHz/ZJ7BDES51SzWQHnTENTymB
cXyjeXHmR8lIdqO3b+YqEl+J8JXjwVx1vl/IszZUuVDDLd3+zqKT9XvmzZRgi0kRhK8xzXwH7cMo
urL4PkyYEpUiAEKTJgKWTuOkUA0YfaTroVC7pEixs34tJpxYL9P4FYValhr7nGZsvD7IXLphoE/p
wEf4S1uFtBxcK1elO5nespGqZay6gmVPK7eete4/9Bt39hV/tkaPFhImIIfLt8dUifTJwg+rL3lf
hvz+XmLztSKbOgF4v0lWTLbWls9ZzRjnXwYPNGfhl7mblcMfAFi8RiVWCXEQbmlOHTbu/18gyQrm
VEbgh7MayHaIh5DT64kN0fl6qMrhEsIg84S6y0yxyCY/tH12KExom0ZpC20abM4B41QvtHHr9JtT
vTCrn82T0qymnDTS360n0ktbCZU6hWO1bYL/rsKn9yhPPSXrE6f8j39f4cLYXzPA6YBUYqfV8KWY
nnPLgZFS6jnkP6YbDDNtTcKVpv+y3ghSc3QLcyBalSwhnzyDvhkJAyZLWrB87HRdBoO4tPOTOtpb
dWNOT+X0EIQx3PjN2d55OFz+wBu3rBHb9dyObJDhspNSS8Ck/ls3iZVl1Nko4CBZeacu1o+bkd1p
9cttoKBGsAxV9Und9MAj3TF7h5MmYXJvhV0E6vAolRQ/goiO0kf23orgqBkBiTubfr6tNfoCY/jJ
A0yRMMiIR/+k5jxrG99j6ALBG764oRJbRJfNJKLbQSSZysxAxm4noYeLBGL7teJDGCn/RaoveCSQ
q3hjNRf/uHjstXYyUD78kXGFBjTb9VPd8I/zSuSp5LaVWdUOXl+XIbd9HeO6cYHmMrI2Wy8o9FDn
4P5UZBHQD5EJwy57UzRrN5sR3qCa4w1tVcIw/YLsMu5rTA+LvYLhI2LiN8ZI5zkHSqKJO5neejBL
3414RFd997DtyRAQPmkyovVjiiDE2jx2bJly1LgLYNIHhyQEULSbh5kbwB7YQ+etLNNLtbRtt/vM
xi91LejizxWjkx7tajQfaW0fEd70P9oO7KNCfpl8bzGBDhgTWyT/Av3kza8TGTD1DrQzkfg8aMmu
WkVwaabOGJgFAJ1ynfuzYx68wl+v664eNeCLWV/eXDz2/UkkvFdxDSQSq+xDE7lOZ2V1ouwkI0r0
Pqb7iwl2jB0bwJg4J7OoaQE5PEglXURIVI7CWXhHPTk48lOSLxSa0R12QUuNMmBLHoGpZDK/vfgi
t5aZ5bwuLLT6NboLaEwsoqeM7WbOdxlYYhixNwKDkLVlemKmzSNBvTVRqIxhErP5dr2KrpvcZ4Bf
9jczKrp1iKOEBXCi+WXeXQ+l+uNAuRETcvGt7GqO7fZpN5+rXzVGJAm1D+q6krPQg9d2gnlO95k1
kaoFfTnH972QOW/za5udX/xOBKLKVAOloujlxs2dxQn5FBAs3tOJt0yxQaPM+LDAg4GAizJU4ZDC
BHpShwmnoPNYJWjO1xkNDtaTXL2QZIB29NE9hSK+jke/tomjQBoAabwulg6PWpnur6atOjuo2h25
kDrRvn9fYIjqpFiIHHpqlJQeUf4FU0ccgvLix/CE9pDsziJQtw4AtP7vQ1KVhQtqZayA7e8IE6ZQ
drEfYtwsVz5bfmL+vfvrx7catdFhw4Nv7BuISbk25mcezI0X+8u4k6oxK2m9SGeQrgesi+bf/AqU
v9eV20gc09c6vIxG2XEKoCct1pUdGOqhlGwMYVecwSJhwcrx5OzoLSClsLG1/cYtS5M+522Qzxep
df4Qcp8Z0SG4hagELo7g0zAL8/WA5yGgkv/PHmRzOi8GSCUdzDjFYXsg9J0ohffrvYGyvJ6SNoRW
SK/j/6XTfI3yj0p4n4fNkjBxsq0oMcIGQ13DNgjpG4Upx7QOBI6N5ICrFyZkprZAEA97UEYBtmyD
D9FkWZ2l1soskZ/F8jmcls/LccTpbdXZP0N8egNCcYLvPiI27WXCmxcCr7wkpSa/9FaS+P286YDD
lcd1TQXKBUq6qlrAeGqi9Av8NZtATUoUoe2gD0AhW37ZYjR7BHrFyFvF4t/PoWTxtK3xwlmGFGOk
3z/S53nIYK8rNtywj7B6MEm1Ojo7JRNI/62k7XakKyZAmQ3UA65Dfy/t2mRrPDM3XURsIU6UdG31
E1TXfXnXR45qtPhvulnlxUpSla8h85ILfysDwpcLRRFNqtGfT9VhQqVcdz4A4Ryna8xmpOKsMLoj
ZqijgXQqrExCKrssNVyJLVh4eOKrUx5GaBwZW/833swlPy63xrNjLzWKGE3G6bxUKWs7Yrlnafrq
eBp4Xj2k4J1z24Ad+9Qsz1+C6yb6OQ6MS5efBXLNN9otnoe4NwceziIR9FpjqwZ2eVr90I4oo0qe
0KAYBfL8U7G75LHaDtCc0Xms+uO4s3L/IgcL5ZqDkjwZohH3tDEl3dSWKaLixFR5TVhjXHqtPyIF
c6CFEe0i8TC6okRo5WUd/HVhfUVPoK8a0o/avSRXR5DW5WDjhx3j/Z2HHIYZoubiMiYkY38NfeJl
8b+5QAvQi4fKVSNyERtVlSgrhoD0eiCVHN8uwufEG1a6Ggn1KTml/GIKEhUIiIfNg5lvJ5hgJfM5
r1m0KqdLhO4Do6KuInSYh4MHEV8C5/9ROXrSQDG/IsC/DxI/lSQNyfGkHRzpdftPRL0vi9xjKmil
geGuZFkScKEVKbgrD11c2UxNBmTkYQaWJMLQfM1kXEEOmjLb07YJ6WeheW5E0QR3bbXCBC4Dnh+N
rc5cqKX3hbu9NvilprE3outxiircCoE5D1WJf4VnC/LnO+Y8mHE3VIgBnrnG5+SyB2hB8LRWnMk+
FM8Mb5txj/yNaUphzxw0xEjmRjNbP7LqnI6cL+u1P/75q8ZGXIpxMebQf0DUIqgzVWSVQAOhZ/cp
dUOgWC9GvPp+QjkF22q2uBUYmCHsJct13g4kvUJeiBEaeMQBwyFGIbjR/sFfw1vgs/uVon0zzyO+
i46xyekbM6/MlYUV9J+Sa4IplGnNabQky0DxI5xO/9/Yt19+a2JHiJOf3r8kW8Go/U3J/iihREzU
KXcl+zxHptQV/aO2nEiIm8nkwE2vfAqH5jyjFt3vYbM3kMTaZNZhnSzmMQQ42D7rBobda9ubWsQN
ud1lYdYCGKkpBwH5iWSfPYYA2PTAPjxb6F5NZRB5zMlyzQ6/yFpiKom5DnFOwo91EjULubf7dVtj
WNjWURsguSNwmM2pn5GPRd7BD6J2e1Q/8KAZZSc7v/K0yiBQ8j35ZJhgr6g4b03ELguqeGkjsC79
CFkWHFevd5BUAbYuDFhh1/nAOuTit400JvvSR8Pj/Gfowz+tfgRZSbjTHoirde8UXULgDrxwcoEN
SMAnNXNNlrkxJVvfjHS+QdZIpmufA3wHrwALqwoaVdMqr/gO593IocWBtUwd+qJGayRgkhldrEF1
iAqLKYv52OLk7sfeu9XI63mxJarLsV88PKJKCSxr//fxvZZ2kKNa0NV+n/BniYsrJg8BsgAiaLEx
NbcpZyv/1qr2T3xQNNi3SImzOXfH5kWUbw+whg6mjuTZq5jJtEQXJKrwqhx6nfHCf6HBZ0Z45HR4
cXpcbOiYz1JfAmFceebneHKHdkXyVvxVur4n/YTVqXBIAXaxvp3gpfevsyReTRuhVnlg73oezO9f
B50O2NIvLk4gXN6CObjuh3IBo/LA3IWLCQ4WSCrmhBUsY9YHPeJRuZ5FiHANTtB+CAYdfz/JclF+
qHGei1ZuRwZILW2EMIMcclruVBM+TZentEbzuCc3wr9ZTDG/f5fBbquWN3vQuLzYw7uw/Z0xp4e2
DHfOr3CTYaGbVbf1Buuu2ivR5tyNky4g+8W4sVlAzMXIs2WkgL6jeTGeqIrECsfNxXzzAjznigYc
7GNDi9hs6RCGTujw5GjsJDAmbJhfM7QC/wvwR4gwm0RYqPyeV8lLEPHpaxei/AVRtpTO98LJ1QqF
1qWyNEN3i3vV+4CD+nez0qOR+JCa+JHu/4c+66uVM1UdJdr8plVhCXnDFBV/chnRg4QlWwh1lgDP
xl6WQKpsd3PWiL5vlwJikcmGE0w1LmKuwUwXhImZaZ4IiLHwzVli8uZW3VW/eryctV5bEMIJpr+D
pj8PsYkdQKW105wtavGKYLOhbxDerJCnDeQbwfN8wk92DhjpXTYNTbAnl6RMkR0V88HUOmrbPjrb
Dbfwp0eKdZvCs1FuFDOb1oIlIt7FzmV2DymjRQExld1EuholozVhSQQp0j7cGh2gzyQ9JqCjoZdX
Sf4h31E6i4sdf8vKsXm0bVZZa2BLTIFB5oko0Uscg9Ct3ycvyXE0FzIilCoOZJDuwJCqdFeLGzih
Z/LCo98Vl72sJ5F+cRMZ13Qb83ZIONOxYlOtFtPTo8Q+7Jt+SZaHms7dRh1mFVVLcPajYHKbStKk
r2ICHQEs4JzI4OyipTGztLiapP1pIlKNIYcSTaG/QgmORR120AhAQ3sutQ5/9bHvBV5T9PFMlUNK
oBHIAYuh7gtebzb7aCOzpnS4wIFEsqTt66fKv0afkBUFaM41qdSqV/BBSovT43kj/6fD+HB0v96P
k1ZTic6VLmxRzqFOollS0RRctgjiWJTfnyNt2ET2P1OKct23X3JLvSilTeSDlx1IsjIDbLsmbgM9
062xvKtntHiW+FgknpwNgAnLhW0MEdIYodXENRBOrZTWxBkw8wv59oIywX3ml4guqmYj1Q57uLfw
0U0ZlW3bJ0utlhV1kfknRlU0/SZeVxJkuq/ctxvo+6v7L07EUyEz45b2ytkPN/Agr4DxcD0iv63v
BLfg2fnxd+r2CIuqKQ2BQlDnuNxtnnywnmerxPypKQR+m8BfgwfK0c7AwEI1sQd9l2sY4yHSN0ae
1HFP38o5R3l9HoNGWCuPyDE33r2ERMcqLKI490bw69DGVReXg+qrDV+M7Df15Ib9FaIr1u2MrHjz
UykoU6kL2bb6M4CjddPGhqio4AbQK9Io2roMXPLBqTQeU7OpSmDvItaDWU4dliD2gSzsV4Yb8eno
tazg/MtrkVw/80E1mDFD1h0ecauiUloN0cY2hhweBDr63PvqzmHjV8AnOtNc3PuHLkZ+N3se2p0R
VCJvjT+bz3N0wbONR8T9dPFblwoD2KLTsNLA2rAu+D4Z0ft8KjsRTKViZZGgUDPwsj1+h05C9kIS
TzBQYnP8po0NF5H9tAtp4gRGfUyFo04rtb53RrsOIu7syYlyU3gQyQTueio5AOJlK0cT7RelXTo8
iSudbqtoAn0F7lGrMEAXqYPEMs9mgh2ZPF1ZJD2+5ji48nJZYYWgglgrmV5CCosEzLKqjxfWXO+h
BdqY9NOVOZnmzlZNKD4EN3l+2+C1MQBb/EPqOxaH3tQYvFXdXn9otEHyaayZHI4gvQvCGV/owmwg
1qH8kdCiceMXVq5MU0gmHbRJmNgOdeUcTj94LXEd3I5IbHZOU/sHE+wIGXk02HRHP3gUtVLk2tbE
eIJd9ccT4HgVVYHVB0mq7NBagrO/DvYSdeo17pEfhBaco4NBfKHVQqsRF/+nvof85FdV9veIYCS5
zFgQXX2CzL2ofxsLwtJkzrAgu8lyG5GRKFebTO8oWfEhrZnPakT44q8Le9/YLiD0z7sxY0Nz06Ex
Ncj42pw+Igf4BKZHwqdkRFr9wc5uXzvjdUROmUpG0SbO1NNtKWTkdnSELJT7aJ+AMqRQowxViubd
gkPiwHJwwc7aUvOmwrEE4D9y9Fk+e3lU7NJwHAdHFBNvYk6pH9mwjHp7GxVfZX2t/QdE+nm0m+hz
lFfKYk0VKASnLSR4Tgj43TgYdiJRjVWdrMsRgg1bJGt+khOqCaxGiZQJXgvfOvUc5GRhBqYfgkxm
7L4fNVvo7R2qpS9sDd8FsOXYESY/FriCVRpDXNk7fG8aZpuJJIAUGzJfFmPeZTfJ4j7KtaF/CMvx
2eilvH6CB8yq4EltmF752h7G7EIFrf+UZOgfE+R1yk3BKGCoVbhwpqkNOrQN3f0tiDGnMqDxG6Yo
K2qW4UKk9b7RlLHzR1pIHqfsjcEOQOKtt4c2mgyxqeU7mO+/UZl1ncaJjGhUZHXxwzHAcE2DA3DS
DnPKH0duMST5YQb8cBPb7ftE/iKkfJNMGNfcVVnPHMh18aQGVGi3aTjuG/mUzAtfMWvUVVa5GUPE
0dzY3ZbqcGjxbDa2Sxqc1YYm6lUGaXEjhKjQ74TJMT7U0BQnNBjhZCtZFjTRTMeCKsRlJ7aozUwh
jRWNZGYIdp8Wd0B3yZWodqkVJrYTXQP0aZI4TZcGhtP82IjgJNR1r5aeO1w16xxGANrilAQ8QsV/
Vlw/B5+bn4QA7Leuo2HfNx+P/yW3IxD1x7f5D7FJ5ZahXui0WIXKSraIdl88lg019YEwZ5QPFP8P
JSp6e9wzUeUcAAT1eXKzOQLwQiNQ2AJUWxN28oXGX/0cqRMapEX1kEnAmV4gKijbHnmYocBf4Pc9
X2sV0LsOOgICdWbuVSG2T69Wa9Yx4zTbMTHuURSMZYP0BwhqiVemnF3/rUz7OtfXPbeJivH+eEDt
6tWGvbR45yTRbAxojBw3eay325Ujjwz8OBnpFDeNXQLxMqF6qUsTTVDpPwo4vqwDtHS7V6qRorn+
cHsz9R9FfPiE32VdNSssWL9Hv893MTk9lq1abQ54zpQdC218NvTpEp5BeLk4XhGjKpmp0EaojUIb
55YJdDwcMPX1S1hwqyBXPz9iPaMPVTVK2yu3INv7n8qqXfcxaVPyFi0AfAus2TfnSVNvJDj59d9e
mOEt568P+LHXMzf3wGmrU5NIYdLLS0V4Gg6bMzPb30Zf4cwfUTvqyCCdj3Gw4YH96wblMeC8PrqQ
JFlshGTg8+nKqDQqaKvj6sE2glzP2HVl/TbsgJlQ79IN+GzHKL1MBUEO9Ux0VgBDHMks1F/ygQui
GfRXL6d/1iwqS+F8dFqKTezsYJITrWKxP8JUSz98ZlywhZ9RpKPbQOVH9bP5qUSzI2vBtJEvRbFs
yYwHMjotV892XixFIVczbCh7eqDX/KXHzhJxZpzjWqOI66pKyjV62dHouhx86CHSRnXdlmo0E4rW
f835X+T89Z9oLfF72O/55SKYBZ7yEYQMIICoKk1OCKSvyqH8UIPe4hR+E4tk6dm45wn5IMThEzxj
I0hKVIY+aAhquDxVvXH+3WWWYoT+rMfUmgjGf83Sypl0xw6lo+wcKDinfRDcG1eHkoo2MTy4kr4W
FywHuh+kB+4kHuqjhTt2oH//mLG2XHO8OCuOXUqDL6tasw9cwjULFtdACYMLS6n6eZPzwia7F8dS
KOctLC9mZ5rvwdXOn6BExAGMqhzeFmt7+/stxMiaPc9Md0bcXEmvY7WKgadnFenM/CwWG2Ssd3pu
AGMg+OR/oGg52yBBiqOthrq1yUilv0CYsvQ49mbXhDYTlPPOJoZ1K2Le1a9kAJ0aZtLy9IMfbTAZ
0upgqMRyiSymVkzPJh4Jr+0fCw14+QuDdcPToXFAHR4ZplDpj8In7WNPPtTK9HLc0TRBqkcSarfa
uNxEhidxpemWB3nFmd0u5YJz/YD5pRvR8vDDr2+FA/3byoem1K3NflIsChipJuvPfPOSHvN0E7qt
T95VZoD9HQDH9fkRpZyV+F63VlZvVoNBBvncA9EFrXVpuOF/f7RYXeqsc6AbLLO7FAEqhxp8WfGf
GOGI4JV4qwLEfykUnm2L6RsKXz8HI/k5u1Lnu5ttW3ysBGPPrVEblE3uO0LLjJAzn/JXERKeBF8v
P36srtpAVhmc6rPy0Mc9ZGBGkHb9pFhCReuOp4zXBUyG2UllH9Xavhug9FIfmHzqjcXy+a6Wpo9V
kB865OAGDJVwAF/PDLE0yU6WTWsA9Ce/TCTwNn4lXPFx0V7LInLQWpdpd1XowNsOaet8scT/2lsT
Y+V2YQcsbrDeHdAe7cwdGkFaSAM40neaDAPQ1mS3f+4eRNG5u3yGatF7R1tUCg+mIIWHCzRnqMPU
itFUVwC2mPFAm0FeZUCMgK3kndQHUzNxbrnGG1gGLOAmHEIKVBDN1imumO9awlwYQhdewNVjk8lq
nQYrobfe8yZ54Iofh5zDtRYucOLdwWmGCh9zqI3lOfuFR9X9esTZm40iryIpRBQQcZVqzfBZVps1
caFpkwBBWVmMyRJr99H2ubiipFp4uw9CWcRQ0Y2g4b1Z/6xV2DLqKsDzbfqywsx05rEicvh/8m1u
21NKVrLB8OkKGrik5dFDSuEUSypngFe5YZK0fPFlEMVoYxmnyIOG/nWPOwqghoimEWDfkznNtLZc
7pTEFo0Cnd8hwNozakTgfHsBJr5Tkw8EcYYJzjt8BKhHc+sBcUzddKto07eUNRELHkPhgKqk789A
3xEshWU0nlzhVAq+vYuVvPjsrjtDHJAGBl/1y6xEM/OeYSB1b0ugUwTXOYD3eXlk2Xheioso72IX
XzXI9G9WWNPUQe5TJ+na7yEav2XPqLStZQde/5AKFMl+zOBo9qMVy+gQujvOcXaHZrIAqnD8JC5e
0905CNWSaFNNMwDHyKK3qczs8XTkVCU1ZP3HPYIR4toTFEgmnUZViwZTxPNlLLP/RM54GYbITYtk
AC31+h8rJZVgC9d9blCG+3CK1sP5S7Gn8ih6NhlPk3iPbc/Lr8gcoSxCHzTl7o/ZwuJQHUgOfiki
6LCP7TEUA0igpOIi+2jzpKRtHWHzfXvbb0PkhbAdSubzdjiF5TnwKY13+/Kg1H4hFhQG+IjekgNf
JLe+a5/uZNewuINLjw4fOQ2zznkZAeboltnOm4ZDM01hfpuwO3tL2MPPtrv5fdVq7KqwPl9dXdIw
c+VEZCJxf+6ScMNrcvT4y1n6+OkZDnrf6A6O/QchmZABO/jzLGyJZOfS5r4mX4e+GPnT/o0Q07SV
Jf5duy4q8oCoRgPLQYjadjB9hpsC3cMJTcx7QiFiqTQEZqvfPbI7gL5jAWwy/GfHNl4fiq7bx2Dx
3iTT55Oiz8ic/ndqPeuMNtSC4UFFRVGT+cscTGcmuAjy3e3YuUZ4G4wlzgY3gw40BU5H2DMmzyZA
/6sRElj5qq+9jvz9ZKmt3AViOB4IbLbG9NqomUEjl4Ug0YbBKz+mXXJ5Jv2kwEL+5wqjBU1g1asf
K7z+k69nVW5GllZ1pN6Z7rpxg6reFChpbtNHhgJqhQUYlPqDngd6jKhD9kD0tS5+Ef9xm2Mna3NY
sh+CrmRvV0qG9pbzfd/EWhXjm/6HdMNgFAkzSPV3uOweHha4oOHRX9Es0oqBOvTtjyRPl5nUvvz1
cfvDCugJAqq34FeiXNRLhVQ+XRlSXNW56GmY4kQwLUNOvuNUv3S6ZqQReOxW8UKxa+2TUXhMf4ua
TWaUs65crjZO8UUYuO9uZYLPsgDGm9aWEhvH0hC49lD5W1PyTaBaOITgEsp64ciKwXiqc6cayGxT
CLwQgvkCCqt+MCVzKkwN3N85XqzvNKtR0qDZT8iXsxy7wq9t9s9pzhxkXE3vBGV1M2XErOlsgU8S
qHpGFbGZ9d5i+xnj8kTW4TOIKMcaB9q/v0q7gKVfaAVAlSXacdXJg10fKtAXtNAuhMNDgaOB2rWT
FN49KAge7uL76oPnL3VTrzn0f4I/hnmxxcOy/ebQDO3K1t/xJETt8XVXEjh+2nrjSwJPPmHn+oG2
r1yokqlabszrvgHJnJy0Jp6W4IUuap5TVsgXOO+6HFAL98cf8F/Gayl2+e+L26BN9AngI1YJMNd4
RPVSGvKOpA5GM1Tn7bSxp9W9klPHclml3vnlWhpeyhXoDEOjC59DMvv3G/O3ho2+E61upOxrGO3u
weDzQsRVPv2m9pt/QT2pWXn3Qf+c1ujicVyzmZbe/u/eZGq85BUGvZ4i0RujH+AUq0k2pUjqe6jp
kmjbM7wyYCDGUbTQ1P9Ec7+LbhQLlVZSD/2LFUDsoJfuT5DdyWsGnV+0S7EiJ5Q1GrflvEBH15Y7
UXEAPtLpZZIZWrrpmabU9794zxnMGJPbOyEy6Yv6XeNQCyxY4Z/iBOwwm/ObxCM+ZUvitN3EBdzG
Nri6DF9fNb8gvjCnShrkqJfy4NrC/XbjuWm1T5SlyWQa5BbHNeiozRN+MbrGK9bflg8AIPfT6w5P
Ae+BvLtZAOWSwPpdlHOLXe1ZP8FqF8wDWz6kGRyLUUDsGAUq1fwg0UIqKaWzXnW3eOE0ub1YRijW
/6fmms5i9e+0k5bRQ5o1A6PhXRtX8LlRoLEZJVi3n8iIZIM44ITdZCWFxEp0BTTuDf3yQ6ElgWPV
ATv0GK1IqeSr9wthzr+ckixPZHWozTpMgd8GXxD1crCCYuUsL4cgSon46L20pw96PxHB9ctiMuP4
OvbdBJ3lJu/4dllCctsNvSTZfnx0YHKYIhgfO7vWUYHHf9EqA3vf7Z4oJJ74N3nfZJ9Pmj52fF/P
PeHkEbvEhyGdNASHqlaKrqMNyA6Kz6FQjB+ULLu0JdRiOfGf8vlhZYrp31YlNeg23J0O/XAlHH14
T78ZqG0f8U04H91wSNfzVGvkhC5eLmmrsOxryad1+LBZDDLCWEWau2HckauKR9bWJtUsplA8h+SM
Av5fq2oJlIq8shcj4nPAROqD1M9UYKF1x0lgo5zv9RPAkRsvngFwnL/8OcOfL6aPpCPBZ3wscP69
iyeF+IN2lMCxScHvRZn8yyE1yxtygq5rJo2JopQ1PD/JPxOypn5qrEweuhFark7bpccHR+na8dzz
hOxxoaX7o1E2Ey9DVIZ3UZ0dv30tdahKPV5uJR3LhTy5+qjFGTr+l+uxI/Zl+hEjNJwsaHMLhUKc
H5FbJ6i0BPYjT9rhYTtiqmZZgaQ+crZFaG2E9kumrinuFD22VqPrbh5HrGqfb1PFuCsQtradl00f
pSS3vs30OBIvRu13KlWI0wO9SnKhdMUTIWR5qLD74Z0v1IlCSI1r0t4c58vUszl/ku14FrpQrtko
rmKom6bgcwy+i7h60bx5cwMGjebZCDPnLGuJbREVxQ8e2yKo1StrzAdePfaGTWXzsikQ9wEUK+Rf
lybFgWTA8jyp/vze6eVVbdy3ySlHCOVj07Ui+54bVH2Si4G/OmcMBOhqT6DPguJWKcWYQPzoSRPw
t2eiYMTnzhh3A4c2IXuESYIdOQw+kQeRRCfETr5map0WG3DVvePZMTPJffiHXE7YmV1eOdrGld+p
Oeh58zTb/0VDZVHyExOVDPKOQqTTzwtRVU1fLIydH0oaNrmxNyNxv84gWGmy+p53FmgKPuDNEMjg
GJPJPzsd0kqC0Yu7ssTco9bY/1f7dYBV2K7/f46AQDiv4I/XzzFQnNdeVoeigqM2kR6lcG1w/pqU
YWS70ymyyfutbSLv+WgK402drhBDZTJpTqio1rmcSB7YLY7koAhA/tRxqMw22gfUcZfvxq3DKQDE
IDZeaVCO68FIzGT7KBQRI6NSCLiKUJnoM1dA11P172ap0aLs/LZn1eaRDXATIQPHg/Btb6+iuJB3
dpMZJ3My1nJnizhB7MoR59Xys03uulqrr0p6E8O+wyoS6VO8Yes+c30J6tQI1fWbnsGQQ5PgwCE3
tOuLNLF8B7y8xw2RueZVVWBDWBH7saeR0MaK7MgZJ8MAhH6M6pA5ptZK05T64mBhyAQPDDFgEd4x
OdG5PL/5Lp8gxCNZKeW6d4q9Bbl7BBt2hJPt6q0OJs7XAVGNFs6b1HJJdRex9skLDSAdzXHocWX1
xYRICbbA2Pn3nXwW3CNp4A4Hn1ZGxyftVwvBVXjFfInItWYfZ2oo+E2Prug3Fj9zc6WyxxJ9WDod
WSZ0FOb7aXFHZ5knzFH8J13KRk55qdiSbd0xSKDCubZKXy2okwDuwUJv9dkKNAiwW2PGG9RDSz3y
p/1ntwPQuXhriroQamvpfsiFoxrubrHHSqmION/QzSspS0rHwZZyN3ymEMaBZBakN99fTV3JHmU6
7YmN/CkHQNNfcz8AlUJYCrgaAyzbRwmOcKbFRC7jZQcdaUmYvCx0cUZNpWMkTxAA+/apf1MdEDIT
QnGn9tNCg9h3pYDWMf5c5dQPM+OBI1uJYy6KgnxtWFS3f6FaPQxFQod3L0OUcqjmmwKo3BKaKofI
D33ZQC1cVXK4OKALBTKq4Lnj8qAd3UgOgFRQZl42TUTI/fst+TIedUoyquVEHzouMbAXJSxNIQb+
693WEuYps/oqAqiahnv6WGg70NoO+ZfbfeJJPSE7pFp0nxP9FgVToWAOm6LpIx4ZHOoiNflLbV9V
4zkP9BP+wHbtHT9LfHQ9otUV+B72N2QW8WduX0Y9eD+HyjYsPiik6rB9EBgFjQibyuc5h8Ttk1pC
cMDjeg/l1aCOihjZN4dmvqeULICykTcmLtT+rPUWQLNyNnG6+cPrOFE+Rmp7qNFrHmPQe7yOEFS0
NeCEOrsaD6TFX0t8hrvOvP0ps8h7HLXqSWsDG4yprYMi9Y9VPDRsDFHZZ8YbjHpmodd/jyiDTctZ
GkZqzyYMtX9vQ/dljveCjDaDSr8vLGEfWG2Px1a9V73ImxZ5Rg1ZMf0SWwFA178OiX1g+241LLQ1
Qonbb9X7JgQU50uL+WjUBJpzxEMO5F4LSBR0bMjfjG8TcCs4GpD2+iMttPiHp6PGhN0K8bRTgMy3
SjBsScuyM07z3/eqFEVFbUPYVhraJmgiLyA/L/+sUbAQikDjC7WKKNsrd/tVEbSNSiEUfLrzxX9b
D4EEF0JBGoDqRPRWKtztsuI056e8gBrxfHrSwrVASH8KratFnpKUCMw0886+lZmxYeRrVTHn9Oov
Oir9X9rPwU0mJD2Rf99UnOuPL9/aqq1s3Kpd4NFKYQW+9/0u3uxr66HkAZOUj9witzKO+C51z0kd
FOFkuPYM9Rz624aaj8A9aqCzkmQZ3IVM+9ZHQktrcTOI6dS7MqHOSGDfHY5AZBcOMOaHUd1ISABf
KLVK9LUYxNZyu5MbNjgE3Ahj0fIVsHJQoTCfrbipVgupKSJ4mLVYFS6+Jo2hjHvmNe49yZ/ahAgQ
ZaTdqrvqpnnhKZl2uRZ0AALPpbT+kycGbtGRCDxW5LlOUbIAImjS1W23iZg4M0FYVROBJmmfpWqt
SMnQhBGQTtDu6TgecG5QVyifORamh8tbTdaMnsgGfeW4CDIGBwFBhIasgbxq0MDTr66rOTMjA3D/
0oLflHKVOvZqmS4E3CCsXTe4CsDou5YAZx5FC0UZIIOdvPXqRR6NmXzrE2dtegtgTShJ1qwvOX+/
biP3qH/Qu1xc//PsD+ckXnMuH7ifqzXFIkqzzh2ESuD9xjw2RE1Yidw1A9UTqcz6BdT+wNf/yoIC
CeBSYRDyA8RPAY1RB3zbJH6z4qbV+8PKZaahET2rOmgaWLn5s7l/ZOHPOujH31LkgzcbAKI5r4V+
Zkf3E9W37vRwt5k/+3SwTTbrF8eZAWUBxsxUADgErikfz9FmIb/cyTZD43CdRcjSWOCRbHlPItYi
4tt04JWDhSnL24/dFYo9jyUM2zZQt8rIOGMa16HcY3QX2AH3IQqgK0HzTm62tW+V4YKzx/ajkJ2b
vcWxiKjQGkFdmfnUTZXhpghwhRmW0umeCeIue7MgaVmsGUTpiXvFVKviUZifw/etUZlVFhfGjU8H
XY3XYuYvhrKeR5KVUK+hMSxdJj5z0UZxGTqFWB3uf1AFbdg+Xj+ZhkArS5RLw/RPRCcVYzEdhGMI
Onmf0fdbUg72GARkCtJqn9qyjFQNIaRT7yJx1saMBwBLDGZd9SxCPVtd0tGdXYZZouu9IeiW+749
FFy4oYi+bXPt+BAkFofUGe4zJIh29AQH2c/DsoIrCVHSCDRwhQDLAhGDz8OUFPtOwDSPqQIXFZht
onTI6QAxeTZdqjUgChwipPxaMg2KoghLOUCtozKNcDzjXO+cicgxGCmHIShCu7uSuKD+HPfw/7Cy
ObFvDuKuCXkQF1b6Wkrcn7j5EHz8JgeONVONHXf16Nuut/5DHDn9DIiFulS8BSFPr3cTXP81hlJZ
q8IJWjg5c152uC1UKnPm2US+zDTiOPNnGBH2Xjv+pntO2rr21Ft/iGPsnwFZvTlSzg+yYOkzKur4
+jxnCzc96zHEC0KaEK4AuuK5Iv8psJRjDzy5BdPUUFKhK2/InCfMCnxSZlklY+Dmk4DY8QQnni3S
8Req+W8vtlKuSfrbNiWWjgv3us+w1zEd9FwdiZihRApBGhUSVmFcF2cY14kYOXGRKBUsgEHrCVNG
P4RWH1gFzbaPaVVWfjcFlEWyGmvCPYIrLnZbxcmBPuGglHZ6xY0isLpTyrZOT7uT5haqE2SUiEl5
8oH/Tb1CcjaXhDijYEuPfEnuu+xsQX6Og4txJJPRh1w2BxfY2vLJWSTGgeKi3jEZDORvdt5/5XuQ
Mg3a3IuYmt6Gv6RPHG6Af5FB4p856WkznaS2GzCF5ahMk96IA6YCOdykp10r7NyH3V4OqQ1ED5Ir
7pZOrmkEgGbVaQOwMlVhZ5NgFJqW2DiARfvb0oEdf54bzu4y4T6Q+jBWWxjI2V5vn06Jv0f5PVMS
gP+jW/pj4dDK7lM1V4e7tEF/qzaroZGR9q5ZV1mUCkVVsdu/XkytuZIgRo6ANTZjChOmgJ1HhTXm
LmApHWn/R/sqp6sBDbO82TF3lNinYwl8ry17+AcsbeceBBgzWMxJumBObzvDlEea96cRbVyx/Peb
lDRWUJLUeovczSkAtMuniVkBgSu+S9dhIrynoDZrvE5bsAVLKIsccPiMeq9R+hLV6Hc/7MCqqpu6
n0UWf1OFF2onc0XfQD50J6bkaLn1TizukmMXaIxbaf4P+fJB6qdEjbwpH723ujd3u514X7EtqoHl
Kjn+wfFfcQnHBGRPqBh3Kt+PHKbASHZHCap7ADqqOXB8eXAdcnrOZR1qr9tURWVYinpECgHcPFMq
gnCNq1CqpgP2RARd+hOnK52unZCF15hfJLjt3/kODywfTXgpqe5hN0AjScTHv0Tk02XgVZ6PbLOk
HQtvCjUnLLIxG0kXRMQTGXA55v6tZNxXumhiKZA8LYF+3EJrXudBdzGwzAVDAnfQYEApkLaWbo6x
K35MJ7DdmAoU6OY60FhP1xtmf0xgtFn6F8jlTtUQy286YOAqnz3raE2duUDMk2zLwTB6nGpi9Wmy
L+gIYzARtIjJwBzM+pqsaJWfYKRIyEBeHvLAPiqXRMrkUoKYOO0NxcgGI4Z7dlOBAa5LVn+a/1fp
122UBmOlXASgR+SQWSiESAJGarwoDky48vIyGZiK5uBHnGT/E6NaooaqzVHCh78H/8LU+Dip1Rv8
Ml+fmYUEJmMGh2getovrBeQUs/AJlOzsbGyRiLY9TQ4MsO3uz+qPjXQflNZ0sJvFRtL/u503N6Aa
npZNJcB+4EdjDQX/5SC6i77Yu8oUy+580thGM1ibhD48X4g5M1DMfDm6rWRx5p8Ud55bPkBa+j74
qYC2VWKe1NorHKbM3139/4RfJN9qlEvOmZ8FCW8sLxLmNdCAy9MwIjLlekwdrAJj/ybR+sGFJmXt
T+sQG9aWQ+nvM1GHvLrVL8jiNSRVhHgX+GPiGE9i/jSn3nFu+gzc5u6/HTyxaCOGbXw6ZD2wise1
j5LDxCpbQOjuyP3HsUW6PSQoa1n68Lj7vWPh/LBASKwlsoGZylP0vIJrBrWrEykaWcg4/Ofo9zyy
sIMC9St2qzrrGM3EJ0T1nPaP3D9Y4ijQG9Oc6Aa7RKbUmba95WW99e7FLFZQNSo2pcu1gdXyN8qh
OULaSHNSmaCjXJtDyHZ5KyFCDa8T+hZ5TqD+5Z71WFR/8WVR4cZGfMD7UpDYHYD1XVLXYjJr248Y
76yAGdhqdzFOArQb9FAORMqNOV7d6F6+aHWhFMCCQJZhGD8YfjnJ9Js86LN6y47PfQsq8dMb+Ph8
H8fLxSREVPDFdCxe/Uv9zjoJjOwDXpBCT7YKL3kgTh2I83zfzC/95BNcb0vTh/GUIo5Hb/FTfnwO
etex4g+XNGa5Eehz1T+IBp2zjkbkvNGDbwDsujcsbZWf5q0ihFssqnmo3d+7DhTnwL3Niq8TMjAI
gLj9FkkbEIKJUE4d3/xtqK/MMauCzdubFAfJ0199wSHZVlgSHMUdVvOHlKMzoT1tz2u7houUoUlh
BymFjb8ayR1rY0J+ZgGtQzei5DHTgJeNu0Vx630VLj28T5C9n3dpEgOmiTf5+142JJ0CicX51POf
7Hx5wFIibyBoW9+guhorplpmFMT+dyFykt5mxIZ3leQ1cyFmEdWyl772Nzq1Nsg+wiSEeje3tdaI
0fjcn/W4WtCjVQeXb7gH5mJw46/vjfv5qrvQP/8gJ68sg82K81vGSIudek91g+jdS8526devnk8l
JeMntXu4+8cyIOSJgrUmDpLwnkvuTnSt7WPWIfLqeqOHK7M2yaasKb2+/KM10BU3BeVxmIVQQSj4
nej5UxhZo912DlwmQnkNOUrr85gzy7jiH3UIDmr2Faw5nToQpuSE2CWP34WLWE53dR/wLrDImRtR
JO4f7k1r2wprio1pyMk1CqdZVwiy4pBgJf6wfK2huRb8FdcjNKpf//7X5uEQANYEMesx+pfwZd5v
F4XJSuGkDfQW7gtnEhMKEiIpnwxMXMinIuzEqqR4bxS/0SkvX/gTUINAsu0git3hBvFLJx4YhSYd
swL4uRONDInDjGe1HR/X+HDM9wnxIMv5ThZ+2tkPtMRnoWDGDelfcdROCkd999vwg3GVF5phqwbm
h7Ku+M718tL7OSIhhb/zRKErg8aXssGtkkTBswM5Kq9U12lrD0bIdOm9W8Pedi5Ry6U/TNWjPmhr
LixaFPyVOkJv/F5AbbivDXOKdH7HJ9PB5eE9lZsq0SXhqaaViiySRGk/1Nzhxq1cL3Qrbgd9p+CC
Ww5aeTOp30ozVpBon9Dt/35YaOyjjev2l6F2IhRW0XX6dz6fE8Fg9sH4gg1E2JBivzc+AoszyJQi
mo7ltQnYO251Y68shfMtN34rVPQMjl8m542NRMMHn+zokaxat6nAqj97bqogON2emOjk31fsegZ6
tF1jORDuVVIZDgH5FtIja2FPCn7p46fdW5F1xQeVxNx14zkXksqcbP8e/S1jpRSbbGq6Gp3dT/Go
iSDxMbXkrEHdBsduXv2GIB4z5PTMzcifr4Gm+0Zf90ebHZQrV0QwhuMDu3kW0OmhBi++1pt8mZ73
ns86JuIpfBT3r6MjhfMT3F3+nDiJaBpFmw0wfftOCOvKuY2ilTSzsChk5vJwvnIS+YbOaWPW3+lC
H85FbRchfrpUB+fQQ8bNHzlYv2t39vB/WnaaaaDQluQNDr0vgmMd9WiVUsLlc8ol5KCS9wSTrR/E
Hk+rao1Kiyu4sZT0ML/TWkbJmLpRplSQl7iDFNVzQqC1rZ1l9Nphq0B5ytAz9mZHZWyXzoDPr+oa
o3wk/AN4DXPorbtscgKGfvgsotGmvL3wBv5BGZV9tWE3fMD4m7jjHh2sjj3IonIsNkcmffukXULB
xq5cgdBmb2Wv6mvZofMhI2nhE+IO+2EemeBfh5WbMFYPdX04805GY84vI24pMuPu/7DT2HqWFG5x
bHmsbHX8yR4Ypqya1+dgmupU5i//uOQ178GEQwThxfKWt55grJSzHQrw0VcA2N1L20q8yQfVLLg7
kIwCKuzvhdhRKuN67E43CUO8COgkcp46fwwr2r/06SgcNzKm+7+D0ZD9kbvovdE+dg1+7djRFCFW
COfOQoy/eGUzyYU1gx0Ac7unLLeCleFJmErLTRkY1v7dkWC6qTrp9+sjd2C44/nWlQoeD9Vq3Lar
3n4Ul9jLtlyRdghAefi+3hksKgsfN8ZdDiR5ruVnqbpxLTiI97oTrkGkpWwPcHQ191/XvxEZpKGD
iFLaaD6HEPKmF4h6JH4OEyzFTV7Ef0TTV0oE0b5YWFwGhg6mMZgSYFRWkc3htLt7eC5aLf0J2GVQ
GFiNNs13HJHcSZEuFPFkgirKwDqqGnejVf5Tb9aamlam4IOo3euTv4n1wwFRj+QDuJ678FXw62WZ
hAw8/J0Htr4DI3aYDzDYtq6SsQjk1NBSdfGZjcu/Sw6QNx08x9s/Gt0+jwat0wU4hARWOc/64x7K
WmHkN57NHi6rSn+7mR0RPzxZlbmqK4K39WcZ5jE/V2hZBkIMnN4hsto4WSDl5RmO+9kEXbOSR+bS
8sT8MxGBafuJPRvo0pfxWimjjfeHMjdNMNmf8ngD1+npatEnevkcYludNKwglzN/gAQ1jKuGjaMd
Cy8xRLjjNk23bGOF/Ntlm8QjVNCQW8Gu2PvUX3uW31uHgQ4H65ipBnYx5bDhhajGEBVVFN/FURjE
p4y4GvrY3ykM6YZC5VCI85LvKSXWI51C1hvc4j1/koOOYUtc4HdjloL0gXOlamCopRT/SzZRhSKa
lkfxQl5T4gJ1O2xQl7KB1n5DDrZL8TF2VPxYYha9t2aS2YB7syTNmcR5TdilC14caKHrT0vLG56A
2lH7w2Q9LLAyhUza3+l829kzU+IzyLCZDEdGaVvUkDYenFwa6gS9wtuqd7LiRnrHK/yPOPSWX7dk
WrIhpW70c5PeJdYMf77s2NsrruDitJC0/ajL0NYNa57/fQcvrDaB9Hlho9qAMy2xzBh6Mr9Uxvtd
pbbIqygaAose/9W9wfm1kzjvPj1aiT/plDlCt4BsNZpmYUNuwZXUFHKrttcXH+byajh+o4jRnKue
N9P4u2snpb0nrNpdSAeLk1HqoLce4JqPVoM+p0Ng1GUYRCQDo5BktNGTv/5pN9ufNoBlid/Wsky4
1GYrPCRWzLJ24cKCfVYOZPSkQnIXEXE4xWafYmQddrrCCyNK0qQ/ghuG2kH/LftO/qznnVtqPYRx
23t9+wK/cqGYhSVm03PJZLscGWSdMPZ8ks7LYysUz0t2O1cSiuOBXmAj82PIOsCxCP0/ROlYM/Vl
WYNugULygo+vdmWisiaYIFz2icCOdE7yCwQ5Wi5f+q4fEq5h6GOztoKnCrru8K0yAAF07Y5pjtmx
BvdddnEngEXwjC/uGPT9ib8xZJSyaJiaoWcn4YzviQUfOJ134k52mIq4vksTrIoD7wZEplkM5Pjo
w55fPH2s6hDGcF+TwcTT1gGoqlw7XHZZnggVW+bfEOdZ7h0vqi6MFXuhUJ+jGPtxl0aLEi4FT5ZA
5jdm/zHIL8NQUF4EhvGosOhw/9cjF/fpHge2FoiaXuApccpASl44QIVsvO+eL7CS+QgEWr+C+Rgf
bJIpjT42meRxEJwpTiGUE1czq7K0ITbziwLzzc55gp7FhRByXPuwDJmt2NYTfGX4IBbMHAgdqGcY
ZsvPT+IP3UsG0Q0WlLhkpZyxhYKksKwkuasT16xbXoLaNW4D/pdfBft32xILX5yp9k7wcy49ghGH
LyIYrKR3aN8j7svttybEeEkjfZQsIBxlCcHTNQifUA+Wz+vtxlPgvjWZKk9od+t80pVVTMdM7H1Y
FlEOP0VEP+b5A0kd3pE5Fl01IMagEdEKGhp9AxIA1aQX0aQTXNc3y07BREiWdkE6MQUpotv7s1uA
hGjIdhbm/+XPsY01apZUTGgnIbS8hdDOl+WAhgY/99JM+8pIHKi00YFTVmuFJhdcnmIo2uT8/mwG
+zEfJU7YRUMLH3irG1GOjQ9Oi8cVmN5F6cr9tnjT5ds1EvrdNw+s7FSO10MOKbGOwFzoi++QSfU6
rebzrBD6TuebMsENTrEgS132cXvcoQ9+IcHzh0RWIXkq0K9INV6oF0Fvu7eWHyQjFqvXHi5f+3im
wH5oexpszpERew8VtX6vFcxq5KAiIxvUuNKUgHV5tlS0xFQNI3luGkqBAncED/18jJ8gLvODnKII
bSvSQRNet8+QWri6KHc7JyH9enetkCQ8t1UTqsrN/wzs4PqzprOZl4kZ+EWwCoiYpwUFKYBzK0oM
Ur90LxCLmP4RBoGHLOuLffff9tniQG4aRm6Tu7j15PdpNaJu353mV26MD03kHLVaO+argQ3RTxVT
nnO6mcHkTU69qncEISm8hpLVYN5QSpoIDTNaH0/SgrkP4H/i+K0MqEDTUSNT+9k0X+GafmU7IRTT
kMAcw6xqsjtnagREXDCI3oFZ/2DUlgSwll7q4mK1A5VITReisE8l9zAp9955eiXXuiOAadNITHGB
usaiP1xgJXtnUPP8FXlohgAfoaS1rteIgnZtg2oyuVrLvEvbiTL/9ZSZT1+xf5meb62DaQTJMPnW
QFH501o4C62D6t1VT7evI28+wI2OWbjlsxy+KosEfROcVsaljFCnqQe3VTU2dotvVmUXbj3bN101
AcbYNa7F0djr9P4hx0qh4z8qoJEUtNgExpfR6+h0V70kKJnW+eWg+oLjrygbLK72KfOp1XkVu4Vy
QbtpC6fsxshOIXdtr4ck3DOrYLaJq6Fp3D3QNrXXk0DuN6Gqq6R5J+o4Eians46DJAK9wDizf+Ap
C+kCUkbcPo/kRxHNloOPbzMN/E24OnZoY9zUdgtsWIqpqbdq/iLFbY1U5SOT/mWAEIdCgVmyqoCW
6UjSXeB4XEZsP3yX25IhZu6wcaEU1nhnthGtqhGChQ8nfmGXG1mXTOclVTTgQ1DAsn9xnitYT8+q
zY/OKgYg62blLDN/HSNKM+U59xb0z4ltKLOk5rgqPd/XVcUeK3DaX+MNbbGspXyuIC9dT5beSTUd
VWU/8j2NQHhPn4kr0JO1UUzFrZAXv4ebstjYIR31F0yPf6y1X9iiHIrKzRBvJBvxUSWdjQDFD11Q
urxLqYvoIDyhLxBjl1TYrJv2+jIAJx4c9cxowDElfCeWWotfF1graPiHHiz8/8B5hNGaEK8sW0ZF
2qbob+QzpvnWHxQAG5JhS/V/PGQw6mexO2iLY0Vyz52DurZXJnNlN9mZyEvOGh4G+Qm5rCnFYueh
p5frIsbVrvRx7O4u8RHymvBxOA0wrPUTQKOwFJi1CNpAXOnb1sDPA9Smbsde7q5hIECOrWcI8iGH
/K/zibfXwPcARHVxcM8AbPBemJgcNWxWqRW1gn22LgsLmfbStu9hhQCeQNVKIec3mJQqTdsOEcle
uS90eX4i+VItnV20kyM4GAjO9WrudzelbW10GDPuM9XtWqz3xu3U6xiVOoQfsnZCxzxgLRogUFtU
62CD7ddGOtHQq2DYA8IFlUR3QHk7a2xBgB3W5mz2cq4rkCRHWXE11EGkTMzetN5ZIj8SAMG5mbiu
8cwIUHHY3Uj1jGPEYJJMOGgwvYHFqzy9z7DAowNXDOCdJ+bdTAcubgib+Boq50+V3fhTEvngjHoo
Tlne5yCesrDXLslu4ClYVW8iy1E/bNGzz0VB3mLvk/QIaPlrPoHGAzZAOCICvVWHEDb6hPw4a9e0
O1biYUBXH8caBcfRnqJydQ7mgMZLZNL0wpjcg2ineGIkt7ltJOz8DsCHNQgFkZIxxijwWSSPsuMX
Se1NkqNmP7S5X0dSFLI7mcgW8dAzTG8VFucT6qYs+X1c+qtmbYWJEYCg6z0pd+0RLxfv4eh+FsnZ
6cwDJ7spL7QRtmSa8mmBdAj4fju3INIxDzIAOorG6MyEJlReZOCk2pLNrK4WItZRf51hl+/s/oTf
1QDCGBed+xPB3Nr9aUyHw/ujD75wVIKxpQc7vWZZTRAb1DWO6Ooq9+pSulSQZRuHkedloOWjRgb9
jYtftSZx+hvcUucr8FSFFPJQnbSIh2DhGSA9U7tWHJQUJZSaI6Qxw5xnK3DSidzS/18riW1Q20Yz
tAEfQWr7DLkKtO1TKzfihSkm+LVeKuQ8+gI7coDGzxFUSAZakSKzeLgeVjyxv7TXE7PEUEvs6BtN
5m0tP2X7HZoxNEc6hSWh4qO7iHUPhv4P+G8YHQIxQ+aVoJCqFZKOzNu8MW+xhxfHMU1+jHUqTZwt
WVZCvpNLjnYNM5v0f0zBqcYDUmuQy+25qOhHHiwLpue0/nvll/e6kyfpnfsfFyoGHpUCyhexK4kD
c7fmoubxtGTuIOUuPhcc2uJkB51V06BVM6S05jKZO2FLf2qq6+qtHcHK1nqcMmB+jRuFAYrL4se5
h6aSWrLM+Cqj0hS/3JrJ9BhLzs7nddebSxz0zdC3aM6YZOnMOgsIAHABbgS8WtKNtVsiv4D6RC2T
2mTh3EQrqtKVshzkHaxwCAj0PZe4znb7QeiSmrEGxG6XGsUOrtbhjRVoPluu+nGrRIZ6zF2RaaRB
T5LPGTttlQHEd2vO+g4KwmU+vNdKCYtON5IKGSnn6c3hIpsA/W641G8vWxwdB+v2upnkCdgPK91p
iznsameOl28O/0oYNJrXkerdDhj/xwg/X4Zf5q0uXwaSz28BW+qI2BoFA4i/esOWaIfSAghM/OdX
ZSCQRMVJqDhg0QuLSsK46IC//svUDx3JL3Z5oz7mdrN12jp1UKemsMhIPBwNlXIiiRuX5mcu6+RE
mZF8KqlSEIyvLkga7p7euYxBkekjjpwhdtPU8SMoCChZQ8cYgDDzJDYQosO3k1FfpMcF+DeeX3Ya
MM7gXuj3SsKENIxLgs5scqDl/sNGPPa+i9tVGdLkgMaTq8Ym3lCPitnr+kw4jA3Dtts7q7IHVrBQ
DFHsFo4C7RgYJC1Rba0ic6/Wk6PFtPh4OMKWFkoMOP2CrRqfg0BN6E4YYZbM0aH21xoeSABP+oGW
B7q1YZvQuaBqcl5YNqUVT5Vj8H/8frcGT3mXchMmpXpQaxjh4GrpGbOJc3ETCyw3BYpqovm6cTzX
Rzil3uCzt+ONCvuzCdCI7rPjfpcZYErfw++tLrQk/RypwAaWvc7VIQ2nEz4XhoFCQfKlsPbqHOvD
Iw7euwxud6OgK4AkhYOT2f9Rd9lg0GdWgHKIpHRmMlAW2knwuUip62iu7/ffdLWId/5y4kMxhK+J
soeh5LsuNcqHhyNA5FBgIkLhWww9ZNVjXcBkgTJl1ud5qKtv+QjYKfedFwG/xD3Est9eIMqeZ9Lz
gi6bYYUbzCnxyuiWj79NhbkM3WUWub13CcB063jWs2Y6P5FQrj0nyAlOKyAgjr/f8tam7WUd58LC
ldyQVvrzffS8noXnFcGfQPepWo+Fv/tKd+P7n35TjpRgcvXpsn3A6GQGcPq2HHqE4qj+cyRhvlGB
p5LGdt4yh5Krx5/SARMxpRkK0nncLnUrx3UiFjY1oezSpWiUp2XD52Pg0jeAU/vMS2nZlzfrbmJz
O8yTQtatHr6U4U8CJCsmxmBjIrKdzyLyzYLRiR7DVO7YlhG3ZfwUycr7ievM6fFRr+o15Mkmokah
02TOIw+dMl+QXNLoCIP+KVMRqcnxseBPBam/2f4CSdxRCBfWXfIwD7IDfwZ0eMPHKEEztt1TBVGK
2E4Dy6sTtVqCV7xmo5pAkimWUrwCYXBfzwOcD7CgqO1z88jLhmhih0qveGIySQDRIXBpxN2rCW+G
TgMSJr7fGwxU3NZgmvtemTDYAH1EoC4eJ3pg3JipzT/LzktP6V6wjHZhWwcJ0CALWrK+uYlTGagt
8MDvAPZe+ZPBsde+U64bQ+Og7DDC6wpHWwqzKMKPYkHysTi2Thwa4tWhRu/Tanx33CbuMD5O7Gsb
L3mk6KxX0RTlkGpA9n/W8ty+DFrf1RT6O5X6phJddNFICxR68jQxnTdpzMSHGJ063Jvic7vOzw7L
9mU5G3KslYbeLlFlMZ3fhq9OGk232UVn3zFY+tqTc3UOiNjChC54sssMPLgKehJ8IFTkWSKyZk3S
k/2xn3C96cT+6CGNbPkc51F1mk5suFoZVFWqDY/QQZqs/TNci3WhKU4uJnscgpYxlvo98vQFxrLd
PeCG5y9sLTU9iuGGZp1uPNJCrWA2DzyH+6UaOz2qXCwnBHcW04vF6MrD0Hyup3Om99Rq1DRAMUwJ
TyP4XYlwfcjks9aq1ElM6um+dOI8Wkqa4aLV6aHIz4WBGMo4wDkHkPcvYMkGeyOctnaaU9fXdfzi
IGZFT2QXL5vo+4tb++ixyjguTNVtxKQk3p7nERPqBGssTKNTU2jvpqIIXOtlTR4K0apg/Tu12hLM
R2ub+S860D3WS8gjkCqui8tpUMAKLBMB69+1R2W7JuDhZFczLh/pYmZ3AMRFSg2Se4O5ZHWcFsIF
ht3Hp2m1GYjyBSsZHLOgyKG719SFP/18BvTKS1zkyjuqm/BtM2pEE0ZfBrGkkg7OcpsiqwlEfUTX
IX0r/oDL87yEn9+C5PLYZJfBN1GQZJfb+QSosjds+tQXdTk3KAm2M4uH4JCyYPW3nCqGdv03scOd
7KOeCmpzztyLHNBlkbqcA0LZp9CIvR4y+luzENR4tdDheDY1OxW7JMKktYHfHE9WLmEJb2uRXK5B
zn6zj6/zGwHQ8haEAKznl17txW0uWI/U+g+avccTuprcGn83pIb6+s4vH1eo5H++7MruTLkTEdkB
UFQWMUxu/PKLaC2ug9J8QCokimHzah9ya1JNFjQxNuCDNcCdeFydTkKzmJIroSY4EABZ+hRtPolg
YsOKup+GZGrmGY9yR/a9rJeajGSDZh/R8wf/zrVbk+cem2uFL7wDqgsXBpCkWkeCLljGu2j3twsi
Z4idkpf8HYtbFIv8JCLtoYMX+ptZAYl80mg9fvBt+LvAvpkzUd26vnosY4b4JISCnDnXkql7iBRK
IbK5VauGaZ3JZZYNphKs9cHBayjY8oWJxmqrQuWUGP2N7B4X+mgB2CdihVIv1kis3tqe4xHudr+h
S2MRkROxTwS7Z6fUi5EmgdbTBs5oNSFQol3Olx3qU/e+ECr8F+L85QDMKteaqFB/j5RYwNIZpn+2
5qIly0xEjFd14AnIVfgAmQwdrHVkEFiRzwGZkAyLqN3X4qIzcGSbPVBrGoOYn7hL8xEe/hzOrJdR
+9t+IUC/oAsacB/6qpUTVB6y0u1s7kce/Tb+GkNLBIJ2Rh2+uZNiISiXZXyd1Mxq32vsZiXoXeoH
c2quhIuDhsARFPqpy2JdXCeAfMJYW4Oyu6b1ObKGOP4BREIKEQ7NzzX8b2IcGSY5LlgTcOYUAOGi
aftgWkT4KNKd7CPm2cRIHU2Bzzr/xNkqHM5MvEWDX7LBVqC/CRwsyDXrIPYYbTmtA7obc9wp5i4i
enXd6M3w95ATkvFWXoG2uNea2PRdSqdp0XyJ/GEQz3Hve+S1h1ONVfwLDfubm2rkqvGToQVL2wMA
lz0G092M6sPWNJ12vpKIFHL9PhZhjUOeoGtYmpWLOGZP6cqN4YEPVVMUdgsXGXX86jxRobniivxw
QCLXyQQZsxRBYALlvdlD4kAFWEsE9qjk6i9tht8i8s8B92iKvMH5UuKRgXsYDrUKjschsGcE9tZX
dWdiSLZ7KOxWGv4fpMPAdQ97Dk9l/9EWvAifZOv9Kl/U2wxiRCxKTjXGiEgKlJJmIqVVqb3kjkcE
MVitAlpkSy96JelbV9BG+swS/1lKMKqbC4vVb50ZcqLZ1hiAJa1RhoxybvRBHiWG3Z4sw4tC9K8d
qkPhpyTiWQ/092sKEVQoTwrQ93Ty7b304VDFCoJkVpiO7pRlt2zcgKyKfFHplIsIWOJlELJRsTFL
VYrUQVR+j2LICDuGf+w+EmtvGNhBr0JO/w4A36NNakpqJ0WIhh7EykRAK5uTquE4MUCpwhozsxBx
PxbiuMYCcGTHx9l73/O8on3gZ4JOfuG7SlcQWl17FAECgEe8/PCy9IdZvg99hNPRzHM7LeAM2hP4
cmBqodUFK6I1VSAbUm87dY9J1W1W2ZkmjrgWxX+wYEXi3DLo7GGt6vqHIY5emsTjM4uJ5luwi+9V
FiwrW6uxOmPXzTgeJBJaZcX07XtUGkt/hVmlUM+9S0rC5HyfvHAJf8uuEtDGSCVUPB/NQi7dXFK2
OoWfsbap2TW+zvgOEoPXjbnJoWpTu/ngYGyJZvOKbGm4Vktw6uom8KM1JsTiepEBfSiM2KqtrFXv
B/xt08HY6WmfNQ6EXeZ1w7kNlYOr/kmQcTzMeTNX3Rm194pAaw7t28X/BvCaueHulqwDPVt1xJEc
xVzI2GaMKHkrggIJbPUL5svKGRFn9dGaB5H9LkkN5LOsLxl8YLNdX3f22FbYI1BiQggHBL8yxKbs
dx9zZdoIf9SCL/lQqiIBvtSNPdGVdEjXSdYHP9BX4nT+UNb0gYbs9ofADHGE4MMLJDwpppCFIkKs
02yGPUQelbleo1wzA0AUHxqGFsc3NksYyibVJVra1IOYb3r716t4umw9Bt2uASQLhXwMRtlN9wAS
kD9U5xKUy8xJZei0iGv33KzN9W3cZkgP7y0u/SO7cULczJfijqYhrvi5RBxG70Aa1kEnWq+NVaAO
FaVoGJ3KXd7X6vAjFXY9fz+04w+sVgVcrDdZoI1X03ohe4Fwli6PDst67tQDe0E1XKRO9LxWEC+K
/emLtZuOqNBHPUxL1xMEDRmc1fTIZ/kMf5wDVcyC2xVXiHTY8ydZBniE1IRbspyDqNNTJ8VYosPM
GlGJiXNMT0HZxDghr6hqGnoxtDXWt4FM8fYkXrbznsweJ0xdSKgaBu12//kXE07NTVYXr3q1eosR
3PYZ4OWf0WX05/8Y/9LxYHX9O6sMmPscuEWS2Va3cou5Ao72iLAmZurQgL6aEhWBloKZLH+QX5mC
NyqRBB6N0jTAz2aS4xQUsWsR8S7cI/WH7RP8GEwyA8JNoCAVWZ1qxSgKO6gDkVoLCeToin2xTHcP
9YNcYYXzHf9ACS8QoC3q9lm7S4pfvGeERbCAkCbkZ1pEcGc+V/R6sfUJ+jVfvoUtatBsrdQ4zQ4E
lQCWsHHPJFkTreXrxhmO0LiHxYGZ8pAoTLfomOkIA5FN5xpwoE+zoSLf4zj7yDdInXoWtEOInrRH
d2C/BkSrZh05NLai6X182+UBQsrVvXHUnFXkllzpTlwYyw0SPIh5UoqVBOhXj9DbUQs2jsEU0lgU
3h/lL7dHow0zQmEcefR0qUo9K3QOm/DUXle4zNJFJWaNu/dbaMEYCW7Ji+gW2HrzEN+RLwe+gsja
J8L6WsLoaTqrf+bD3ekAhbe/k9kazXoHrQcUERMqGW+0/uB0shhXrd+r4NlUDcuOwIhPL5WNGNCV
JMw9WPArB9652DNZxsAxLYfVg6nkFfqwM24FRZjV0Cersh2fTqFkTwWk49fqWnqKfiUtRpzSBNCB
NMQgzjvS7X+u3QFhqXgxkwHFXNUBP0GJ89jSzjvpBWxj/n30REZsvVDUdwMgw8mKPk5Qx9k1cybR
x5aia56YK4CUianSjGST0HOG/EJ8ajyacJdV+8eivHoVV0ZOBVuvc91pl+L0m/Bkv/f6oW6/NAIu
A+rKD5UZKSe1cWD/wnhMVbhasqwnPReUjYOergtzQ+UJ8oUEUfc87/IHAO++GPjGqstlJRSVivuJ
HnxIB5CVm1MTFR40pbemcvYi0Clsbzx3NAmPRE/zPkYLHRhmdZJDZOk2FvonubeLoBc3lmOl+X3U
Qlvw6jd/RshV0C1SSw7zHgCO5sIUc22iGn62899dwApnQExgBrGz9YQTaJMrXMAbM5ms1Yge2X1X
7rB+SjyuZfQX7fM59HUeaizzJlbwRR2FlVJdy8IzzuAw9sg2QbBDcNobB7A/4/OslOL7rpf788ek
j7D8uEcR17GJG+pGtNVP2FTwUgHXaq07ZI7FVQioZTL9+ZIPL8XgwZ/ud8GJRV+G4V5HYLMIA8KX
4OjuYoE/EfqHR2nDMhKnzS4uLl1aRgnIjDHvza4vqzngtQb3eJ6L5AdFtw0cvbHc5wxevzGcO7MB
VtBEwzwTtKfQ1eePDNEWx4h0dj0YbRIslt5iWIMIEKgZVLuFyEgDHKVskQSqRmAW/LNP+VX0O33a
L74MZo9CThJTn9sa19TwTJE4GdrZYigvj9eLVK5XpACQ7QrN5BrpT9lhXUqmdW3nm+Ppsbob9lIq
4CZhdCm7tfw91Gy8JKCFunHGVmXBFored1Hx3z8Bgwiyi5g4YxCeIbRpfXBw3UkgZRhT7di1IinV
ysHc2ddpuSLIfiqPrhETRhGnn5S+oE3JyTCjloHXiy6TJlimFzvy1cDQ/qkjZaa/mrGEv6TkuLTb
XcVuqRgyDzeCHSpPu9aho+l5sGAlr36/Jf554W2GC9DyoKa0CTY+2dpjDEz8a3lqL/ks4L+9BD+7
x/5C/6zUcs8sIj7qpiwMS6+N/rhoKzQcrGx0H1nab2W1FNbikzwt6SRe4RpMm+pS72ljw5Rd9IzG
JMmihTLt2/+rYucujHkrZzzRb0jvElJDWAzx67KeaPJtfyEOZIDtuvV0dWwpcZtj2WV4fYxL+aGg
vuqh8nqrSfrNRZTCm4RYG70Drj5lPzvQWk19HlpqhB7CqyeB5h1xgPIih54O81tVeUu7EtFtHDln
BTIA/cefeC49UQve64ZJMbSJ4NxmoSmkCGKKsK/yFvDw0M8wEjIVQzwt/rH4O2W2xdqxD4QICSpA
nrtiSYyrn2Vhk+ok3F/VeiXcZTePyVTPtVFA+iF3/lJnXlzg+jEzIxs1E9JnnXxrhMVmYpRe01u5
LknjmjpQmAKst2/2n7Ffkb/Ew1Ailt3eGHRV10N91Au7yMBm7Pn9ih6EWQ2dU5JIkGl54d7lXl/Y
tHxSaeJLAAEnjQfdw5NDERDTchiMXurwuKB9PjAFjcTkdOZi9bxUDIe1+kPV7s6B/dbVVo1tHd3/
OvRRKPMsTOPk8UaZohUNA9IV5qgKSFnyVSqtc3A0zNiTMYRHOdBG5wt0AqhjDu8OGhP7+7jbPukD
Krf9BaxNxeTLOlXG/0983p4GbZ7F7Kocjwpyk0oPcEchRgP+9sRX6UA2bfV36RccfD8iTfqrXnqx
zml7BxlomYnjepuff+inFIiiF1MBADWx0o8872CbdpgDcyQqGtkXEP7FJ2vlS6RPO9WrDNWKO8hi
rg1Rh8nIqqzMqvFR+V1GkHHuYcCba0FyJh8W7nh39MS2AxcPUCYv1Ypqv2mfSBPa5J9Oa6cRxU+X
BTfI+huQ50wsi0KqkxbyDnNnEWA7tbPfS+EnDwYy6gXbGIf0r2UTakojUC/UhJLULYnXqBRzZ2GQ
njBJkH++avvqRAxEsjDIDtjWgYjLjejgugmVBiRht/iLO2y5zcWHHIQ0jpejsNYUDHanRKQrPs1l
0WLSGi79pe2aSGwrIdAwOZfLTgREentivwDvAD3G3BPl5rGvuk0soTD2fIcArLcuRB+Mbz230WKV
bWFmeEGHX7btBQDXa0IBH/RtPjp1qbdVCruA6YKVr/xEHhMv7Sn4rMjBcVN0fuIJSjfPQff0GcTh
s2HIaU8UDfRORvjwk+3Puv5OWptL99liYZaZN5lxn63WN1u+6+KMtmILa2yNFJ3SiL1CXYhNZTiE
96XPXd2IHVcT4k1AdL1WkLuiHAW38L+jE6WCNob+m4yPjJUZ+uKaOL6P6Dim5MJxq9hUK71jXoWU
EE89R36aoKqszxlk+U736J3Avl9JAG7Qm9Yx1X6faQ4R61RTaGZtnELbicoeE1JfcYj3q2s/CFwj
FYTp2A4HSQlwVLc866UXjfgNn2qhHoVdKrZprI615qWS8s93RlSqDWSWiReSZDsKS8E677GTLY++
ILy0Y29MFQn9h2wX/tOjIDOxUyjVV0XvfB/KI8lBOxD3ouIP8K5JT72yzoq3iU5oAXztWoTOodxQ
9uYkXwdevIYAteTN7+J47Oy5nhannpWAZ24X1qHJjo7+vX8CcG6tIqbi5+D5ZcD19kJOaCJGMubE
6fGF73mhsEfROr5mjssD//nj6ApEBnYeRXIoSlStFQ3Jf041USrh6fgy5F2FjoZF1gLG/NdBIHoW
BjGYjLFUY8BDhUzFjdCuUSl2xbyRhPnpQnsuV4KKMFUGwvrGccymXR+1nk8i3mAxkmuT+dNalf8b
S6En50WUAP6Dcyu4Zx+7saIRfiPsa4hi56aOqybaVrO2pPU4b4ZHYsUhvWvhrPC915dQRrUDGdYg
xQ8BhO04KPkzeCsYXC8g72PfePrvbgI9YMXZ0hq5K6u6j6lphM3eABOtQbUbPgFpYs3hkLZ/tbtM
+SoRv7t+pO7RTKXxqsm6vxtWlL/nLY3KiiSvrbawpuae9tmtFHGmWnSEsz1WxQHNeNMBjZJddo6L
Gxx/Fyw+6SnzT+k7RMaJNoJGR08UaeCpGJGurG/yUPwbIvGKyqSMuAQQ/emTs4/xZ6f80xro0aua
97HaLcBLMYBmmxr+w3SPSkoYKB0C6ZG45P1l7hVmbLN7lPRfuIrsaIjtUk2bYu65v4nERO85B0rP
/AvwLC/SUrlg7M7wMdqtpmDM8+aoBV0m7uYj5BmbQOH5ar4vTIPHCfie6iCz0ugTEC4EyOuOcVgz
NkWoX0ol1Uu1raTeGV/qSqNTsQOWXGXASmsdQgpaoBo9nFgfUNDHDAoAI32viBNqhGkWPibH79WL
a837l5Sl0H1AulhvID1qq01D2HShaBliVBo2PA2ctdmAfsenwuh7g4F//oH7azvbT/iR8anC/MEg
r9h8yit6Mek3tPJhv5VqA1/syA1IsBhu98hDGQCVnkosUdQ/czVj/s1p7kxgInXRGzcnT4Co3bbk
dB1BuQciFwCZlIjnNyvH2zZ/TN7fsWajCaZL8hGU82qh3ZDO9kEecbHdvLAKPv2tXCNaJgGWZbPs
ggh4qMni1jykSw0/6mGxi6wf6ghW2RX54WMbQaXkCDcPPQvWuzm8PHeBLd2tt1PmmLJJ7ADDOJX2
4REeobhwxFTUz3hFlW1ukiQyyvCKSsqRmjXVg2lT1t5Pip9PF+tepUpxYNjKiIT3ZWC8O82LEUWh
XeYB1VOGpokC8N9Oh9qR5PyPXJEvnpt1WkYQUPb729EYxQ68kzs+UATaTmdK3BtaGpWdUctpCuj1
0raZ49KYRtQtuSAOGwvYMogVlzgwyHKQCgyCCklgislIzKewMrZwf6Yzkw5pLib472Nhpe/35wlQ
9wvueYJFnrHp8B1FgpBctaIYZOsCU9B2eZfWdKCrhI66sFi9wY7rbxX+KN0N0BC732+G4G53o+gC
lycLEG0p2MtjglN65iqbLk09emoauQTvlk51nnYuOyIfnQ6wKgeSyu05I0n0PdjoxwN9Bajn2ZL0
kqXikmJ8E0O9i/7p0KGGtODLPm/BpHVxdNLr7cMSzHth57BWNJIuxrEW7PAMQ6V03GFTtet+jYM8
ZKj8WFh1nA354CapYgwNW5lkdC/ihiTrupXCchrtFXkv83xY3KgD8j11lZ3RmxU5sLwaNxev/3U6
LojDRYLp165GeVxx5aoAoynuW4tmTy3vdLK5xExs/7ZUEnA+4HdZUp0x7r/Df+FwMLAAB4LDj7y/
bhr4WEmHdIWthvPas8y/4ZJjnCjq78mJ1/x/RIahQ2zUmixuojvCCduqW3Dhhfw+RFiWy+y5UrPT
1jCkAFPP2b2f/Du32ssUA5aCHlo6LzCbwvrV10ARzLhozhpSt7Y3y7XOwJj6eiJOr//WgE9Hr62q
TJbYj8P/4ObrW0Px19wZ4ZCfjRfqruePQT+58itTrwOpnld32H0V4Z+JJSR2h9YIR06HSvWi+dD+
VxQRykX16kTwspj5HNc3AVkETkFY632xmBCeYX1omW+tN2hR+By1VuyLS6ar/CWjXbpQBF53Prbq
76lXnJgUyMjKLfNzV1KQYIW5LIc7+NZ3R/5YnE2B30ZjBcaR2pDRuFO+RClXms5pKDR62dSGTyYD
IRNDTweZ3QTalDGVPrSs5vCPaWdxpBC7oZor0CT5QGTlB3NhiVrpWQioT/qMmwLOKnA0yt/FZDRQ
cnsaf+dcFqImHMchRh5rGOlAbnkbzWM7pJg4u7SLFNG1CMoYHzfo04bOnf8MepjVCZakiloGm8g7
Po2NuN4E+z0H4dRQBLqqc8YgPtmGC+mXlP6OyHvXElINOrnkYvDcrtjR9gRuBbOH/mOcMYRBUwfM
1duoXxhmmugg7MB9UBzl/TJSqfCIQY0tauVAcraZ641JYWWM1t/DWDF4lauka6jiK61/BUUc9fQG
+ZEi2JdPLBdRYg5PlK5nyzB6CFfvqkAWe08VG6XXJXkPXLvJUjNqH9rcyccs3vjH3k5sROobNnEl
dhIHup/maQB6CFl2laRMk+ym7T1zW3wnifoxxeUOEQpuEiiQYdiYpbMz4svq33S0FzgFp9mOu2Zz
OBCmroaCHQGu4+p3L0QB+5g+5absRjBo2/WveTynkxJ51mJjZy/m9a8w/irKyzHgoaiMQmiVtzkh
7o/bVwHuM1ZU0BPcNuu26ONHKvxv9UCGuVxukOz2Eg87AxLrBDBoaeULp38YcOPqgERxxZuIe530
tCOiv/h3wv21RqOkg+Li8Smi1KMui33PKZs4UeAMnKhrI/Q0tAOd/J1Ixo+Kv3dXSP/cQTxs39TQ
K3YG7wMGZ2JcebywMHNT05DVFjSFN/G5vBDylIDmGFDn8gknAW51kmRPEBPNRW6qEz55InkjWoam
URU7Gwu+hFTkgxJgyZqMvPD3icjAPNKRjknznyRzKvQCuSzxSSSxxRyUyaZOD77nWAQPlK+/l7E7
Xq12wqPevXh+qXArUKDFKPK+kWP8MxNjnQdouknOJRhfCwv7MdTDIMq/rYqS7BHRuISMI/f6oK+t
g4lXe3IRONTKI3LrJOGnc2ZkFiehFVO8+wgCNwyrHtEZYa3BRS4EoO8uOZj/8ZsEjOWRBshTrzSp
H6UlukjSDQjFAHkBDjS+venouLiPS7JKpn+KRt7FLYEzr0CbwNeTmMQwSSSkrQrOnGF46GCR/4q+
3fSKYAiqDxXvE3ELrQ646jObs5BLJcZJl78WMFH2PYBWKYf7AHz+R3H2qsiwLPztZCNHDtkdY4uB
cHmNAO3buquQ83Q2XBCjryyJe/dMjYoMGqOY2P08HoOlhlUn415wngcCUoJrDRFYyeUolwcow3UB
j6qrTLGF1xp5h78nEA52YZCnbYmkfESoPW+j6VbKXz6BcoDZ2wicw9SDf55BK3jzCtG/3znpSwoA
TVJoPWud4jVXlSWLaxMFscr1l6AAyB3r6arDBK+mVXFGXfHfcDwWY+NlGWdgKe5Ow9294/3FWRAa
T0ecFrVD44VbSJ3XmtluB+3aeWSDG73J+LYanyWwEzWr59vthIp5LXL0ax2l4FxTGEpaUtEcLzI+
U9PnG3lOsH6sMc53G/sNcPJWShjAnMveifV5KAfYxQunMh9gYjE4fphfio7pMV7Zk/arha8LhRPp
ArNnpxrWYy6ovlT61pWNf56W+lIcIGZfZqQRlJO5GC8dxxN8rpSRLIscFSGg+MTUh1Qp6B1sXcGA
5IjIglegrrjdorSymUhLrPshcIBzkyhy2BZ81tclN6C4HaFUmbv9gIZnztFiR1rixlcm3z6Ge3Ja
elK0dUlTW6d2+vlZFh1nlVnzq37bSguhfIbjBmJROe9SL/SrCnLBlXz8RVYlJXCZI2BT4n7eVYHv
Ir25LkBarb1oxIIChgg3MycqDo0rJulaKsmuPx/dSeG4g6puLtMoX4RBAtiAEgT0PcVzn5Fn+URO
fJEDRYXgR1eQGW77zF+MkRNXyLPaq6MQBhkkWHuL6Bj2caPJ7GRizn9giAbA4jVbNTa8tXWMDBqY
uLMqdFS6eS9NjKfDiby0WnMAR3Aw+QtcYKM1C5ltg5O0vu4aSbZt0KI4XnjFSyEoklTKGpHsn01Q
3a4hJSSxhrVAlc2Ra1+5bedRyMtU7fmk3LkJBwJxf1HFFQb4rfeB24+piKLPeNV1kstZdqeLoiS+
LMeYSqmQMoYGf8WxLdjQk3HQZgklzddr9Lh0GzaJb+j7Pl7AdRBjXS5bXTTH7BlJnNloC4TS3KyM
KtLJ0dmm93xWiZhC7UJKjr3BKGfDKstWfMnosFyJN9aoqFDZKYnVYc9kZi8hc3wCMqLo4pgTy5nD
xlOLwzZeT2HB7OoSS68s8/VBIB/1Qoc+XVTy0iez20ghz9Qu/GBKuRZQlG1LUrPA9NaTPVaHuJTc
JV5ls+yiMPHOYnlk14mP2eHdOZhY99IJ1Ez/aT0gk/4wWkW8TjXUG+7G8/Z6tIUjss/onLwWKAhR
bmLKDXHOV6ySq3XE63yG0aoSdjPoctnARYi4aHzQ3MuHWrT+QJDzU6lNOe5cqRLZnw8BTDYyWzXc
x6M8PkPkT8I6QIED9ZUa6FbLAturUpuCTXAMzSvJHuO3mi+nWnJ8MpRTuAVJfSXIfxL1nzR5Sm+b
l2puONmj5wGB8f57/NIaYoQLljyfjv7ZXvfX4D2oK1sGijhWdTD4w8wz2OhymFg/M6yUdJ8J9h/8
Odmpu4CScpYmFhqto6uWq51MHdgBPJlcUv+0S8330gf9UCQ/tCsdruze6OsT+sQ/8aev5YKGvNsJ
mRA0j2OzMYDhcyeRHKClsIk8ZEdWF6fdXfhO0snnEpAMhMD1XeIQKxjQTEaMb/CSWZ1eOPPNwLig
/ByJ5MbgdXWXT9qQdUrANc7PrAHgKJRMxmSB9l4Re2pABCNwKJ2gD+Xr4f8lPT+VH+FZUvXBxoJD
scnvK7SmFbmTzHi6jR147E4s/maEGQrBDXYbGf4hGiq3K6KUG4lyLb8vbUglvoGmFw31hXXb5vcy
JNSU0Lm97uIbTPMA7wkpOLHTjdZOF7EB332NnUUHLMQA3X59WqAw1PFMIX89NAVJPLSy5srAU7Ft
V3LCFND7HUXkHNen+EYel8nV4KPa1d9+5wbpl8zNfJXXec/5tpg/GqVuQ/o+MT4yrIK3nnDi/7rP
aQCKe5hz4h+Z+kmAd4ssQtehCmi/5FPoeHvE40eXJh6J9earyE8xVxOMMtPAzmp4sNjQvomAfGVP
WGj5kCQdrBcIlw9qpYKxEtvZh/ZOgzN3omFBBUXNU9t0qEkM54kbf00c+Wa1B5GsOklz7u8xHmq/
pWJWDNbdZoSNQk9P+8BvbGMq5MfcqJdKXRLY19rEb5Y/rdlhRtihlU56wAzc2ThSw1Zjlfcs4oUQ
WsCXz4K8pVV8D8OcJnOLT8Gi4fj0ArLAZ2vLmnTJXN2UAVvnsWIO/uwcaeFUnRbabbjTQvD+aL6b
wtxYHSjETLn3Q7HTcFdZnpFuID5y+QK0Z4oraRqYN/Qs13RmY13cbtX67ANQdJuG1kYXN8ZemXEm
F3Q4MixOW2BKa9erHKTDl7kpIXIrU49AWYGf8gCjdzYI24ihACMT5WmqDzaF3V2I+aCSkgxEhxcM
OLHbvD0re57Cg03aWzxHFUZWQeYqnbB16K0uiANCYd3oXrSoT3JtdsOHD2reRZrS2HdaCVZ67DrN
k4VAvzfyA2D+pfzGj8dFX65eZyb7W5p44UpoZqbHopSiCP24ZKoEH+uzun6QvLvhPMfU9U2Cd0Ws
cHnN46WtmrACT+92T4rZyIocOCnACaSFaXXor3KGFg3ylwlGk8zVRfWMvHk5JwolQ17Zh7rxgiCt
bIwDFIEoVT+y2SyO1R4uw/S6g2QkT2jMSII8GO/LgPL+y//oh7g8Rm2FGQ0J1mAWuNkieIGV0OyV
W8k7WPzOhWT+wJgqb6JRL7wG6zD2kUP/CTBVOeZSiAnJ6J9TeTclZedYf9OuNKT7agXBJtLf/zRZ
J0QvdCI/Ucyn+j2d2ISraZejcKS/+FisOHOh08g0VhyKzIbKLDCX48XDtXXOUIF0ttgI3pe9ICIz
xs1mgyGk0cDGZwwqyhQazDyyAmoAYGH6sdYbcZgRcz4VV7OiXf6Baqi493jvjvVTtR4Av5WRpNB+
JOnmTW4edESGcbmdFRaBElo60jr9J4vOE9avCPJk3/qFbKbIsAq9NBJIOD1sRhc6aINM5Cyq6tFG
WY8AX8lQH6q327TvalRCLx9qiqEhh2m4suBSKeSwFVky2W06/6wWsch62putrvLTs3v64TvFlu52
SvHNoOKiLP9fMN7bhi7qmCP5yq61LUIpuxmTNYBs5CDFdYWwP1SMM29zE61qJ1SwRtlIch37BDOZ
0vlfDracCtDOl4vX67PVadC6m8RPa4s46dQS/HCsI9J/9scKFjqDnhn7+tXDTaUVELDY5Fy7bFXd
CS44dMVCbDIxERuIcBTTiKVDYKsiClHzSsadBvyH2abs0pTyYbpNYcy76LSgwm/M0ZZoExb/x4b9
5EeAVzpKojJ2celNIa8aPCrOLsE7a6chDzm+yISZ9k1+T/e+Y3r/ucVZBlJH7ZVZYilt+kHFz/Bu
+P7rN42tbMtExQ85b6vVtGijzz+nCdIw7k1X/DL8dve+ybmdNNmZj972S7nV8RfeM6bH4WBSuTuK
cO/bb4TVGDkCB6jDVIYwhGMd+pCewMDPuy7DPtDsYZSJsnqSEJ/omRw3/20M54yKGIQa0S1tJB+Y
BcDQFZs1esHisgPUBHk4uaYGjesESdNXep+v0ZmgIHygsenjO62VzMfXMFi8g62luLNW51r2+Td0
+FKx2rQOMkbLa/yZ0ptMEsNA/OThVslBxx4qKArnJeZh7Aq5KlWDxP/j0gRosfsFlmPTEvY4gzFM
w+Su1rBs9Hwi+KobCV3c3+gX7BWeBhia3fv8Riu6UMohUq6vtCAxhEbhSGXc+rq1fXk/H+sDeJuI
hUOxkVTaebP+BZW0QJo5y/82OXHpJs2Dp9uIlpkJRVaDfp4y34qolXjbxdR873KaC/orMW4W66Xv
ScB3uJspzKrB2AmFkUHFZqbTbknipfKa4Vj7fbtK4yNPcaUrYkQMAqCU0CvCfEQhkPZ3C3S9beFQ
TNdCVbSZS/s6CWaoFrabpr39qa/dFBynB/evFuW/Z56rb2g8ZcDYmc+XHyQ7q3J8vM6CCxdHqE9j
VCZz+F571IC3cpLW2a+JJXTZX19WTouX7SlKYspELqh6+klkXgC+XHY5g0nLU0ilAaNHtsOE8dTP
RgZn/x9ttwFmUvepZ6qlLemybRXYKRWYvWB6LnPofwHSwXYwU5u2wi2lMfs+QmVZENxsPkJlB+eb
rQ28Dcb/QK1cvXNsTQ69GesDusM11mwEwi6loHvvrBsPLihcY8YDvKvDbaJbYAlRBiYZdup8pmkF
mf8v+O4hfPJepdMVKtTwqzKNA9bxxs14p5b1vkk5b49EbYjXRkFGOcneNk5BmsOVwIgI/h6FON/F
jF4ga2Hjdr0iGWwss5pWWpv8itu83Yd33JJTe3GzIdgiqUtR0vktoAV0cp5pdwElR6jl9G47sgOs
G/Rb0UHD9Yv7wBFMu4icSmtnH1LQ0KcjzMozF0l1SoZ7hqZ4cTNZQ/X/tqDjciPP3zWkK5wkYGKp
T2Fx1s44YXuYSgt4pw4ERHIu86o8iR7Zz3ZDI/Mp7xzNeZ/KrBNPq/CK+Awt/dZRwsU116jT304A
lYXJANpjaSyMq3i0LpaWbDV1MNrSS2bOwUNHNnktcKLprmctbceRp4U7W8mMmkK3VWoqESfxrZgy
XZC4MsLrWtRhBt2wcLy4kPi6D0UEBSzwcAoAALRAqjGY+9xQ4OjOU7QJ55DnT4/dDhbmerx/LFG6
S90jDH0M3YJPzteo2YVcGbrqIWwFw3Q+NWEx3qexKfJsb/3YYfmo0jea8/NzNZipAhN5Me0uAjR2
uCOVsnECDpzSWoNVwfNuF6P3rCQ/kE44azoOwLVw0WqqN8YNdzc5Harb1i73nq8TX7p2wN//Ald5
SDzItI4PqlSXa51KhGAnyVVqTR5Gn2nD5KsripGM9GSdjeBZswvKT34A6bhDlsU492CDXbO5/UvU
joMQF+5skhQTBziIltqHIOEvH8J0+Y+lzM6j16tV8slnPBi/YbyfLA4dp4zuvhOfBYRDuWfssR0l
hRcSx/6au5vT0Bo5zA+l0vVdN/WSBenM29BeKuMQU4HlHm8ctR0mBgtjS8mPtYdNu0oYYKTreOKe
vWqsV6fflB8e4ljZQmsergiAEFn/aCiAPTLtk8s99wNqVhqXQw5dnbu8lL5i+c9gp8684VahN7HH
2+uA5xZq6FT/TQ22RKILdJsH+hGe0E9Cij5jt3qb6FvezqmVKAkBR/Q1SvKOzwqkpsR2gNNqJTZT
Z10zMtOWXXQD7ewTZgMLIB385zVICbetMqZu1DTUgVMnCpkuRaRfIqArUZ16/fPWKMKluGTKjLiL
vby6hVugfevoOrhL3PkpcqjTrskvBaLAsZGqPQw8IHJoFSokG1y0/EFsIlQ4b04dzW1iQSlURyUb
eJ8hL0AynfqfIWzMxLSCceZVG/dZKpSd5JMl5o/6Po+tVleo40vv8xM4x+edvNoHDKv/NjpgfOin
VK8BZ+kY91C01JqjlxngbR6gT7UO8r3SZPz1Kg7MjKkJnC8Bsiwe+kWI+gclajgNgvHI3lLwDIDv
LEReB8MApakqeC5P48FuW606/hQ0jhaNvoitTDO2aBEWVUN96M3xe+Stfp9cxBiDHwqaquJNh205
5W02NGb/qPdOkA6J2Is6XZyPRTUUTR1XHsR/X6JXXL720L6xtfMp/sr6tfgz71lVGdoXeM7ZS/zz
VgYhfbHHJDaFBd14zkuoV5n+GW6TJwwK+XuxFJMpSt/Id0ZROnGxZBNQ4qelcuMTfnvroDEIRfC1
ebE56kI6mgTgbMST65MpVMCzSG7gJB19QPePKD0oA/beHkSUEPAdj4NgI/OKiQtI7elVHTxtFkkO
tGJdMw+AsTo1yrTJ9KrjbgzaQchOEWrD+Std/M2g/xMES6s13+24aVcy7Lv/u7yDk3/X1fHLzVUw
FQmHM6+LBHJ18Z8Db/u83Qp4H6kfSmAhp5UvuSPOcdWABzAjbJwwgQsBF6fbj8GUKCoMB/VEp4Ps
rpLwK5MXPn4+LbKpWsikqX8qU2Un6s+hwNa16KZZzHcHtm8USg5J4oYf4n34jodSMj6NDG9MZX/Q
i3zBhdUb10NU4KVT9p/Hs/Un8bFXq0AAfwu3a24IR+09xap5aPSVOo3MqBalwcOep9W5rLFjBldy
Hp+OPTNevYaehSyzIECLXI60LW6JSxmdiq/oZ2vw/Z8WLLcNCLe3f1zLPwZBBDk5tOjbTgzDLoK2
NHJ1qbyTePKLMElCEo8rfr/69sbYtK4KUeBrqICwuVtrUdLaownr2crXu2ZE63yvEb+3lN1IjNUL
/PtApb+kJRDa6wSyiGpjZFivXrNlBr8GnErrlYNwkNOXz+JlK7bS7zFUTPWaAGKBObq83ZkH6hUk
KCQ9Nh+xAlGQpjUNmc7R6aSEti315Xq5u9BzJVJwikEHoZf89VjIT8e9uYx4+6VvM/lBCqqEi2uD
BSdsV2zGLhve8kzOdfjZhc9EY7g+0kX6YT22dLtvZ42TRGKX6869ZV0KT9MGDSYdS+uOPHi+SY1S
Js9K4CaWyYDwjx/2eybsiie2j6MGMulxitih5W+fOOw1vdJc0AwJpODIQrMkKH+3LrP3J6M+msTi
rg1zvq4biboBfRA5UEXjzrE7LjbA5FpZKM4ZPklwtNzhSv+38nKvunxZi0DXxVATawTiyt0XD0tZ
ODSAfW603MBJUtfK5W/8ymmjtKwW6Amg9Goy1IxWRe1qowGMePJhnhf53+skenenYoPFALJsq90n
Ur5oBEfcqR/iuDkfBXYBGnmIDX+l+sYBSyYUFBHVQnKZ8hPYEPh2p0lzU2qGZmqm870v43SUxc5K
uJ4dfy/H7ylim2uewLu4gjpqVZY7HEZySTwJCzkPR6vmB94m5ohLPk52ca6w+ZzTFTt3W6rlkwaa
+QinwN7bS5tw3Vuk48rXib98ACSKYd8AcUHVNsCBl/FlTc01zrjDJAXvXydvLpnDFE/w793EKi+G
XmX/O3mGO5knvJYiO4D/REajBSTVm9cJdZnNkWr76gcd9uryMLh7Myn6DfZdbWWFgtaTBSPC/sT/
lvBjKcf0q795hc2BLN6wfj0KCErJXYbwreAjwr3sxx2PXtAY9JelvxDUwBU/Pdx+dUtQA6eofrJv
Z6xJJON11kfizLSuS5SV35kb8jE1znafEwHLoRsBhfU0NuVwpJbjyeWugm/pwBInaQlHbzsnpsC6
cwLRBQ+bpo37xYNEAWtBvr+MGkLZ+1VfdSA6Ltzj9gdFHR3s4RtB+KhGmV/b++bX1NcnQQqW33iP
1DcNr44wNdTRWdQC0fudpxeSu0fo/g03s2QS5iDZ3laHCiHMvtBiaryLRv01SkkojpwzipvC6UWJ
KhIV88vLc0CG5mqCiSNmFz4Pec3Veyk2Sm3j9ULiFHyn9x14CLIeo4JIycm+uGcuzW/IiUzKGckC
svB/biqILsx5wVoIoTi8+wVl1tZhU6sPJT/diPIZZWH4ZA/344nhLMoMJah+9Nj5bG0HaBJN869k
sXNVD7fzMYD66AbVPT3BpDT7pgQUcamYaPK7VxrNriipe2CQeJG/fW5lTMSMODoLlSzR2iDG+Fl2
UIkAPZnegBU0ZmS4ON2zJ4SnA4Hl8l8N4Plik9vQgkX+MA9bAAE/xPUFmhVprYqmLatNfIyPylKz
6kPNovWd1NMfbIiXAuXFlz6/ArY06SpUsuOhRjTrDy5FZUbb+uWj+42sxgJ2rAZh84W6gqcEKGnx
weaNJgJMWPEG/veNbvTLnpGkYQ9WN44snwG65sLBh2mQjm9iv2+D2XxPrx8XJBViZeZ+HatnYBvS
eompm/y+GeF4E2Y8K1xelPuxzvRKKak77GT+o3CDweqliK8zZKvfG1gIgoIf70OPo5kdkOB51qGy
QZuQGsvwOog+kpqDqa86FPfFK4Mk68l2p2ui72Hh7/CY57+mz46wyM4wMoE7S7/R5QNU3jEQiwTk
1KTw0plT9FgMKhxrn3BgPAoJLdfisFW5XUJbuqO3324yjxsVH2TRtqJnA56+q6Z9m1CegLDyvNRN
fqUivV4GODIMgL9Nl3qybwUoAVfcV7uTGBHmMXP89SnMLthyfGLtV/LM9A1RdOCkW/JP8sHViS4i
qvTxSx1hZqm/bcu73BYDLyxcYRbZ1qMWc3BkMJhmEn5ZdBw4Niubk9+rDrWOuXP8Dkt/ad9c5xxF
rrUSE8nAYhPTRbIoX+i8CoW08y3AljKzLUpD9/ClqF4FrdUuxDfiFc/lmCSJNhd4vxwxTEIVt6NE
ZhFoElo2yWHXeNLxJfkaM83yRE8vCO2U7v1hnyn0gEI+RVN4UmG78AvA+5Ln1QhiXV6EKw5tvcgi
0Id6ndbhsKLJpXkjv4XIbcqdz3dKr1UTuFa2YKbACkQRDxH1d02lyMaF+d2YeBiGfWav8KYBTwnZ
ZFq34OZ7CWr8ogcNo5fsJVc8726vCgSdNs5Tl5J1xGNqRZDli5Hz3mFnaxWLvqGcfVYW5azsgU1E
Icin17wUSvx4TC2LLjWTgMpwKJYAddtlAA6fM7sQ7E/ryI6DC/6LuMvbgQz9UYk4t59ON+fbLTTj
LLvbTm8VuXkr+PPzklSptvBdcnVVxo4ePhY1rMPRQpgu+iAbbfdHVR3ylWmh3jkw/Y+yj239MFjK
FY+PAQEZ4lxfIfENx5FnD5vt2riks2JAZ93W/Go5Ib7rblwsBNwJ3IUmJCmbKEZpmR0oo4hXE4AF
r2P0VZ4QNnKIBUeR8YiE2u6KtYDJg656iFPzUbDv3KxRFMpYVFBGONPwmqm58PHmpbEBZCF1BexO
2Ux6jBhDn38tCWlG7gMan+HqWpa3pCEZr/p4Y2v88O5Tx+qu+lzHQKa4hFxvNsrz95MHTJJMZ5C5
mourdE+tyYJA5ORXrQ1oINAPKfoVav3DkHhU/YIIDe6jlidTZShtUDDUQzhvuIKGGHaBN64L67ld
foPgjEqY2phiedxCbNQhA59zdkKfAVMP/NGAgwQjR5dk83jAnREuL2EmQGtNfMQY6vF7r7BSWpUf
ityp6PgY5DXS1a3zauUm/iuafl9eueTNOdjJj5IA8vMWU1km+neQRaz2crGbGiXySrJM/o1dv0Bp
/w1GrMT77BjUJ0wLuHx1PcnaVbvhmK30b66RJCTY8i1rHLRh4JhC/i71z/S1q/40ET3b8113zcQe
UBvMUMgVrahNTu/q+bM9E1sKkw6NeyQO9jEcFJV5j2fpuFsi1uZ5B0CJsiF/YJAHxEfHZLqpEaEL
tlslbLZAszaegKRmp55KG0cXRwmPaMW61WpKwafhuOD8PZQsSXSdhmihmDKiF8VA+VdMI/qhKDdn
2ItnrCgXQpk4hN826Mh4LzUMJWsN0/Rlj0g/P84CCpgB0TYOIb6AGyMmaV19hZrNnJVY23gwwr9R
6A9WHFaIcSyNnklUrUnRtgMgJftFQeuoJVBr66nmJHe/istuB0qmrvWOAc1xwV++fTPsIVGSJrI+
iHgctDZrC0WDk+ouWaRyHUOomCnlLm9IG9DU2yOsT7zjKEU4+iyPq4pkmHud0SCi6k6/MdEO5f+l
wokmaK8YvQpLO8PyLup7DZgd4tL7UthatPktojJbRjVYznxz0uzIgsSb00erOtLaXOw1ruIvEYj0
52YM7EiYDD28WaOsgA5rRVCk5dOWsiNn+K62lB6szRRzyBNoO0ZlB/NhTjB9pQmlKm0tqtuwqen9
0QwQVH61qypJjJGclrHSwedv28boyRZ/njZoUfkNJIjzMyy4of4nrG1NEVR2FucjKYbX5P9SYH/g
8L2p2KMMS/fiTzoUA6jlMHJ/wN7j1II+sJNdHkmgQhLyoE6LDI3jFVJZODd2GuWv4HHCqefuRg2U
OL+PN9s2QgsSaGLX+4N4RIEckTBo/ucFwpeqSQMHVWb1/cXpZ/E1HvvpXlBs/415l9mh6WBTuTEB
8FOMagrKuzaCb4dBsh94UgTRYh4aMK0eYaIP9pdQ2URadS6QB/3XZTIjn7nhiY2LzP6E1wvXC1vZ
CHhNk4Qy5VZGdF01z+YukG87MXCgUoEFU7zCeD82F1EtVIauOSL5vyTu+uPMFhgTnej3b2xK+vsB
sdL4bcgqcMPu0If5qJWsEx7JLWYGUuFp609PUkPtnhed910D7MOEfHpNTWXrUw5N1IxCC0pFxjNO
gdUA9Cqe+L5TXORXmPzDagLLP9VGQ3dp5WNWaZmz2dFnLSeP81y7vFesy2Q1+bU7fBmEMBWHMUJ8
30Vtrhj7NymYRdfaQifSL0eCKXvCErpEb2Ot0mRT3E+mPOcCd0y/X2XoPegD5o2H3BfPFfOEMsrp
xo4sfIADIa+qOuNSBcxsfuHkgIeQcH+9d5Ql7CGOsMzEAH2q8T6fgIyBaM/KiLmpsroZEmoM82KG
1mTI4PJditA5kdVYaHCRrchRhaH2KXjWyZXzm9OryaRoptZBreg5Ag/rvO8Sve8N+4lGqIrENdkZ
aJAT3Yo2XDivndVA5Fkbeu4ADyQLyV9SnRq01I6pEphx3Y9e4i78k1ExzofiHfQfphz7O914K9Er
Jp5ZiZlQsIS4yigzfk4nvhShTJ7MVh+QPFTbhlWIQ7SQArudw9gPm+k93gLh0aiU+T5E/7WiVSTs
4SYOLVAbt8EZ5syYdfy+53asxiGjN262nJ6qsorBm7T6TRjKuk/fokFJNWBi1XPAng8xae8clrL7
PVIJwJO1Kw5azwOCPVAysgM17dNP/NlciMS5DXgz7OwSd7IHtDl/EQRIkWrCFddlgT39qjr91vJG
s4okrJtEdKTAVDiWpRLln24w+y55Ef+Y5ckSKWIfrKvRICQbpbCpwXe3GHto9+WCMpzFg2jmB1i9
S7M09LGeHHVrk4NsXwGqBpFAYTEP6qzCsHCe8wxnS2k2TKh2KIER9eJoommqXHX6Y/WK6fFDIU3Q
FQ2sgi2Puj8sXbnnxVXxriekkjQg5C07m8/Yzh9/ffNp1qoV587rp+6FW+0126kQlVREEEPo1TPJ
Efeasliee9gImvZDWASB/xPbThOVLtSySrf9NWsDVhEPtqwmEVedVj7YrxGR1NWq9VcKhQx5/s3u
cKfF/kQ1CHzsOlkAtHqgXeckxKtLEkbGZS1l3/E0GscB5KdRi3OGn92ZhTqK2XrokTZawWS9r86o
WF37qIC4Z/JxnomEypSdfjcoBarVvpny8GdOeFt6O1eL80QR/xdbeT4/nn+qS0eK+dLdSL5h79Bi
lIq1O5PRGSP+UvzP6yzrshiu5Bq+1+h/nydWbGXxz+L5pZbPdGlYXQ8YJ1xNdekxWsPlfVrdtkbx
/MtkZNsDtiPvJsXI7gfIVP44/pFXjThTOQ8aD6am04Vetr98IbV6h7QyUuFkmvDrDC2FojqobDBb
t7fA7O63T3z9o3hJX2RSsfHnPBU3RcquCtYCc28w7q2Q6xTKaM6wcMXThgSOnUes+z/41WOmJa9r
OmuG4vDoOPXn+o5Ptmy3/bodotFwCh64rGZp1utgkxWZy8CH2g1/UMf2R1x6z2Bjs84p+hbxMHoZ
my1tex/nNQtp3Z5TeG3BI7nSD1mZZQ4Me10fvXu5LvmH7nQXWNjief9jE9qBDu3rzj/5FMUdHrR1
vD6MhBS2rd/OUqbDBOdxFiW/9uER9lSeMFgdIIfpQSo9IH1I5EEI7cc7k/ceiabo1V9lgV0Tk0p6
WRmVkSCBuStOUog7XnXfLSdzS1WqPRkGKNo/2OyBFqYI9J9Jn61z92/o24OTiNieMlM36dYZ3NhM
9Y/aWxYmfd+Yt0PaVzq4xPADtARLq00yNn8mVKthj3M/VMB24snqo1lyMdmc2qsGT0srqtgcuA50
GlRmAaJ3fecv2qaH/1oKkQQmBJT45438RyOUhHWHers5pm1SsUmsCfb6zWwGV1FHQ1/5lp6vV1e6
3XA7Zq7Mt+jTdYlStbaddDBObp/vqs285WwuHtYA22afGTDjEQ8xsDkYeQ9z/W/T0y9WG373i9I4
6XBPogc1NB3sih56g3+Ne0QTiJSQB9aHmRkMz1pcuacxsehb1T7bm05cQIZfgr+pl+QgCsfMOyk9
7Grpf/JloVL3z6w3sY3R58awWK1rtJBn2XtREH/oakEFX1Dh+LRcdHVbgxmfEVRKE++4fbZnPw5b
qQZrli+bOFcfJHNoQPdbpaxalIs4cJMW1xVLRKq5OcwRkAF0V1UNIxf1adP6UYN8Ez/ZbOMG+hks
KhM3D70tH4oatbmnf6Sfaj27EwGub2mx4zCLWTD4Gk7oVcBBKJWVWdPsSTaDCNngSYtenilSC+9b
BSg2Gv9jUIjdsvxpJk1VVsps3cZXaRYyM2kd4vHB9CWJY8rcmZ2SvekW91bWcq2HAImeRk4j9sZH
8KPgiuHNV5qC2qCDLNzldCNtKVqTFP0MgUad2UKv0nFbFO8NuYGly9N6dN4f25wh8AzYswR6dbMB
epyCXsBC4FLOOfJurtRb/pmgVEIznkHqc7xoLoVBrUMbxVluii7hMBWoN6HG+mvZXbXT2A1WazuZ
gWKH1bSup4byXWHpE0MOQsxUkD+fmE0rc5pryto2AARxkKKRkqDJA87H+B0uWHKXMcCKHt5iTqX0
2+7YQ2AC2kg6gplODnsY2EYuPaDrSpz6jQ4AgWQ20ZZ3H++60T1pAem9VBkPVL5Qch129hA1NOOo
FNd3cnkC+tWoBlJ64SpLO6xfdjeyBe+kjGlfWhkiq4oOOpnD8wzXXrPFiLzaWCRZEq39QggXB+G0
eo0xl/YND3q8Q8tYUTN1yVHQYqZgDe6Pc7TuQPpeoumSTW8JpGqGh1paeTzQ1nq+Su8rOG/MQ7la
Xd4Kxltsn4JkWHBt32u3uzbxF/UJzjEC09Dc21+ObNgLfXwnf53Lr785nHVSXVTFdMECxr40ZFTN
VT1BdLLCLycWejE1yWVYebkiN5DkDO1UC99ld2yw6lTGANw0hZA+IQZT3mlXVaA8SAnxCnIYzNKN
Wsp0r2XtsY58f8mW/y5UYB9x//4E+G45nvWVS8jE7tFRbdQClNO5pdJsC2kQu+xQdDNsnj1lMTAa
9qTKXy+to8OK/xyIRs8w1WX6M5nDgPKaPBI/t1fYtMPP/b2ULwrHNRZKdF2ts6GGgxGWJgIjhIrF
P0Fja0MuZBH8H9JcXGpS28ViHRE3/1Mc9KPCg/tEW+ZIo+GmzDPbaXLXInQMQCiWZnwjFlMA7gOz
V3XlA13/kuN5zwafyNBycXebK19RjNGFmYymmiu7iZ8Fno1kfiKjvZ8VNZcNs3yR4X/VnmAiqUey
hmVv/QFs5lvRYRRomV98Xomy2OBuMobfKMcYEo9E/CwW6eETpdkJTBh+OWUMJT2EUrvQ2X1crZNn
vK+O+gWG7/VTVzplQP0BjcwKdMupJ6HdoFVG+c/5Vl5ANZHumWYVXajRnXk91HCOgmCE3qS/Jlow
6f8swihAjDxnoDFtLhllMzvUCKlzIo5stoDKzmQuVVcXtCmvOOEpejm1YDeD0Pa/drw0Z7LHIUsb
LgZTkG2oTGZedsCuNH1tCoDHPQhex/hlaGvzwJRXrGW+BZIiRw22TU+pHN70juHNJfVT1QOUNvz4
Rrz1/cKGzIE2ymjcEWFG2Jh4uOlXqGxWjHAM9WPMvO7pjnlBUpob3XQ7WUzfW70fD59dVw6IarGO
Idxozce5FaUa3Ee/lL+dEzEC+IEiyOCYBlUDUOU/CgsvrKx1ema8GsT1bU6oAereh4fqUVEO2wM1
f7UhcQHz5PWjl2x4UsB53QhEjJNrZfkk/0bl/AhK+PK1xgWLtdN6p77gNJjM7bifwGB92YzBOOlW
EvMFt200c7+pSHM9RvykortMUTsOx6nbtTKNMDuiGBVQwtQXS6OiH8/+BOl93Zo3ArLf31mxAePN
6nP83x2d15tAqCo8Z1ZVmP4xl1hexakflfjcsYlfdb9uPl6mM2Qsw89LtHbyOKNtACM9K3aBzdOp
zZuoicQdwiufeHzU1hDpj+G3Db+2o0oXVx88gnUQiAmgi8Lcn6hi1zKMP/WNBftEmoVKeo6YG3Xc
JTMATMr8ahNNd5Dfr2LjIuX1KRjan2nbShnADB0pRE+D7vCsTQxLMhQE7N29g/bGPZsWbYvQ3D0Y
J3S0mh2JE04Rc04S1g6gruaE4zs603vqXNPJbKhQq4FCrwGbNw9/XORdPqocKjJdh+cnFewjmEMQ
05s5ltGJ64IY10oSzRSvRdDg8lS9CdCoEBJhErSef32o9rjADn9yXN3xi+DKwLZf1XU+jHAuVKUM
Wy2dAtDYRemmJZ5nHKZUbLUzllM9mxEKP+e+AxUtWS4h/C0cJhla71CWwjbFKYoxSYD1IcSABl4U
Zn/92uHX3CVzys1o2zgX/udBMwyZoeqgq6iDtwRrUE0/0MnspDRRmbR7AwYyltLHXyQ1I9mBJ7KD
uouKDiYwviFz/WxgQfpUND6GN6MtHTPA0BSPV7YW1Pz1GGStRE1E9FSorqyH45XNUkswcpTklECA
4JSu6fhQKrGd90r/zEStACKAiHZK1RntGaYhMoRV8T7ShWlsq4nWiNdbol6DEG8oJvtS3wDOUSBa
+AjiPQRwH22oDMoBjrCGDQXNc1/8IzPse8BESV8fVgf0Q4eWEcdj18RhUgGY5KBxp1GjQFDMnMZS
+InHrB6DZz3rnE33kfhioxf/2DFx1OqNEVzhXCOEwx+zReafHTc7Z/HMPTe0O7TwsOmsKwya7PLV
rRjcT8LTVJZaErgKaCCddmAjVgJ8g1T7XV8PVw5IwB4N7zf+dYBp4wKHv2ysZispyaMVCsD2+naF
uxcbDbK74uBG4a8dqwGTBLplzhLCIxlN2uAMbmFZowlL7H5UFzEiDnIYx8OBlwWwCSQqLKXZu7q9
2ArnCMylDZZAb0cCex/gC13WSZ9f8dkMZC1QQrcMx9p7mUmPTxnF+utxbf9Y7emToYuxEJ2Sh+p8
WljtaJ57ozqyg+jJeR/oIsTdCsKmCszNj5iYHVuPGdvX7RUBtFtbu3jzTU026wEho5si6a3h6Uia
oe3ByGrjZJ/YOAtGN4Lr76rlXJhv/KLelSXNkheXOLcsCrz75soYMn1GvRLRsJU+1/hLQ6PPh2Ku
5VGbNcLj3logqtlM94faOIAM2UH2Pev5ZlXJrno3vqdcpdaCtNRx1Z6HruOHC2xEuM16XFthW5zy
2H+161ExeQqrH3N1Ik6WeuD5lughFoTKROBPgNcPFGwTLOpZcIDzSFFQ8Nf55R7YkXXTJPVAXGny
yQsMg+8ln3TYa5lkiZqPfmlTFJegt4Fc99WIaSvbkRMJFc0/HPjwVNjblqvwg3rJfHI29IuApKC9
Qxz3LALYxxGbkymY+VQNlJZyBItA6SGK5HhNUFzWYg0l755J80gOLXYBcwIOc1B9Fvpkt4EWFX4B
oh0CLp964KEuZvVHLl5sM+Nk5uh4IDeH/rrcq5c5LuED3oEMJeoiJKMddIsXEMpE9HAsDzcg39xw
I6MyA7eBUXBrUGuiGnUlTt9aLQ0Xh8/6RTOVQskqCnPOyUiGmyTlhwZkrnsh5wXXYsYZOOoWEY73
XliK09eoMp+0RHsjVK2oPBJGXtiyGNT41dM8jcR3GP+Qs2euYgyJx2PseZAjHRbvX9K1TGLAUHBE
3jYqRshOK0lB42BGwtcLaGeX+YsH0+XnTTMUz8p1y43MiaUrtq7X+0qJuG+KZihDtbqPoGh50IWM
QIw2o47hdNoA3JcGE2JCLCs06ifyg5ZL3cbU7M0RjCiXFlQDWJJJDuVpmOC+2VS/Fw5SWDEjicHk
NcgIFdznvCiUgl+HD6dGBhNIGlEGFETpqadTV5HmUUvxQHQJxYOxSgzNH7faaIw/yK/VhOX8p0Pj
MBn2znMnFL9fJ87kScwYCJnroD3IYnDPHrSl9danJEQsKlCqrZdak+5TmBLOHKyw48U/UhJTb5/g
T8ayO3SRDyL5WTd3U7Skm9u7aM6hYIgHTNSbr+VjFEYINnI35pFfP2GrFGMasHPmzBJp8Kn+q4FS
K3Ufzztrcb+NesdAcIU4JpRQUvVIdQIBahrYWhfaMNkJ7Jm2k+OE9qjpLMI4Ts4wwSor2RWPF1NT
u3J5Z1c1BC424icf8Yjyu1x8L+9PPNtDGrU5XoiA+ze8L0qG31Zq7ngHR7/HDNL1+8IbnzbZvfA7
K1zlVlI1MElm851sSC9F1Ci1gOTQQiNF29Xmx0mU5DigdG353zaBC6dmGCUgQFuW/qfYNdsBrGS2
w1RZUq7eSVrPL07JKPLc+J3XvJev3RgADESbg7lgsk8mxfxcPVFm6cHxWsuwF0Yl8ltnUgCP8AKx
EOATS5Sr7KXFewvbJ56evsUqKo3H+bcSYdL50ZbHMnBuYuqxZoqfXkP9kOFKMLIiM/7r3QJGp22f
ENnkrd8XMqiAPaOfdCXdr4tMsLXtL35/wxJsVZm+jO78X8J1WhCDNljeESWcpeWAx1JSiVhdO3LM
WFE3+e5pv1T0VnjG9Ahn1YBr/LdrDRGL2gaoEvDgzqkoHLabG/nxLk5992Nddrym2OFnLYkgwkq9
PtMeYPCQxnNP8f+0pGLFhNFyqS5inlNKxbAS066jBJ1AuIGPtBot9EKFqfR1uwar1k1P+W4AJw++
N5amSJozPG0T5Yran5I0fJclfbHPswXaI6EI4vzwtFk1QAfl6WBEX0xufcHVPlSr5yrV7qRH3z3D
U/IT9OIM7wC/R29vmD/eRNH0S5g9hvwELjasGFvTPq+pxYE+JlBHM8aMFz/gVtgkes0+CTT2WehP
9XP2ryIRtwdXYkbHPeasVs6L8rji2qH0b7W/MJ8c0UfSA7W465Irq6xB7AiZ7KCfSA509gDuARJY
Jx5RgsJCyKS5flqd0hLkwRCHlkhbu6S5yaJVbVDJ8oRROY40ZPPUcF4PuqXj2YBvkorVTPVKGQYw
6mDr/7SuVyi4stSWgi5s9tuJhQztb+VmRJNgkWGbR5T3owE1fFYSLJOiKZXy2Dx7HuUNhyyVUNpV
ERKg/wBzdMnqyxtTF/QBEJJ5Ys8sITlB6m+vuVb9bSNwivRUHSuBlp0AkdU9A1Z8TKbbGwVs0hvt
Neb56lPy4Wmhq9iDzuFSINivAuc+d9bTvFKhJhBV/jEm/yD3pubA1TYk9Y/oBYBmPg5RAim33tqg
XHwT9SyDGGTs6xj3dY6pEXc5McMVeKYaZyQVAq4o2DyjR3dN8AxlgFehklpuo7ByDXtuhFG22VDG
98HeuZUxqoNXr0IsPbMvihIHzrt4Iz0ot4dsm1IbpZkpBQ44pqtLz8jyEdVoWE4R0P3hhA/vCeCK
qi5InEWV0C0xZiJhhZOCwfLtRMcdvCVQ/xqvGdm7uVbQjULuBeYNSYm0DMn7ZHCC/1hVifJbFMAo
ry4WJte7tKIFyCiFlwhyhVizrGnUzGy5etQ0nrIKmB8QLikpj/6MeDwq3VjQdKtneGUwTHMRn6g9
A3W25ZDX5NPK5s+vckMstE3eCoezdIYYGez0+e46pzfvjsCQvEB4wIfecZp7zMCF0yD+9JTwyFeY
OsSO/iVN+sGzWEO/NWnUndttQljbNuDv/BXKTmZm9UJuI5I9Q+f6/y3yuySpnBKU5N9g+aW1AAYK
14hQQIqIkFUGdGXj5bONw3fdzpa9afhzw2wd82M1V52WKaI2L23UbMUoVz+Guha0XG64TM1+OGmj
F4IDZTS4uLJdAuIcmASeKOU/PBoatRpbVzykSuaGh3GUmjOeYGsWc0eWeOhnJDR/cJctQsh6DzXZ
Ep8D/nMmFfW4E0zTBbHSG6b6dB41yIoa/GCvZyYV2FeI76SdGDP7rg5lwsDI6E74+i0NfkNv6GxE
6mEFDKqkDMucmKX2PA6UnflobzDMBuMGqNhZs7URnsWTAEBQ8rLlQO0QTyHN+aLI324LkIOEcV4T
Ua4fK9EUDtLOqcyB2V/4sreTny9an5BnE8aREBFAS2O8QgKKG34sckFzUR282NRkmCbBwg/zLoRu
cB2ZI7j0AFt128yk8H46sTLaUlr9lg80KpDDfPKDlKPgrply07QkGDjGBx1ml6k5gHkvJUO7gyYc
zvS8XcpE9UM6J0jPUp3HPVYQP8JkCYiiiXv3X2ZHca2ZB3NhGbNy0fESrtlIsjWo4nvcvF4C8PZi
9G69IclLBR89s4UOvWfRHbGaNXFnrtUvNk8ncj3TK15LW4ka1mSy5K1Y1VZ5xyLle0M5bu9Af3Bi
m5vNnxWI+hjkWLgjg5G9tkqavzWx0Bec5S0ionX7gc4/eQ7jTZ6WlWqbvmIfMTEbKTtOMNi1Udth
K1vHHt6gpTnBsj4K/ZLSDdZyRzhc1xhOdMURdTZC3a8Bv9Q1E4rONPk+VX6e5DIeQOdmngyrB+wY
+ng2iO6kyufF7Jue4ANIIOoZYK8LjvKA1NcNJAx8FXhxbYG2hh1CQe9vbaUsHbFwS15LEQ6b83In
g7S9dRiFoFj95F9HFMZmGAfpWs0RhRzUGm1E9626mHfsWqa7rBA2V4Ai/C8rxax0L0l9whw4W0l1
NcgwACW2gENy1ruuwM1DGjV+5NPLqVX7SbdXM5ht35LppUy708sTEaivD3ic0PMcF/Ir/5ad4iGj
Ue3PSxpE/6aowibLjHWwc6HCkHOf2Y0pB7JmjTAmjxEVLiJn4and/qMImALlgypAQqbPSy4pJiH+
hfH5mlxuoB5kqV3W9k6K9wBseV/6t7teq8BcEh8FmoViw1qmC95a4hIgYWI71TN/T0mIHDwIlfBE
3/FEipi3aMDZ0EwHsg5Y536jcgGCvWYSOTGu1v2CIS5wBd0msMcPXCXD0gFl4RHYzZSml0p86+PH
kNUZpP49l5FhVg4RPHYwoju2Z9mzwljEIUEsubV3O/y4kcGe+5MxyaHYltRY5lx5yCyWvq234ari
/jTm28yJXu/nq6Tj34SD6yazvsa4GoybjiQezQjix2/XmrC2q4iqx+s2W2FDe1F4JeF9KW4ArfVS
AYBCFzZcONu0IU6Lx0r9ZJFRTfXuQRpoGC1B4D4OTT5uN3EVY7qOfadRW2D1kttIcg7rRMmeM30C
9P82FSBRW6U1u3XgnGbzrOQr/+uKpnxLKg4VKpSGY5xlFQN7YykBsioFqmOTrudu/D96AigRb1Wx
Pxv7UNKxrBMiX9UcRoEj8f1cTf3OePTNCCXkz+mwrUpN/luoXMRcZ8U5HO3/OM6ojd5MiyKUhPJW
Zt9zzOySJmmoIn2An5RwG7StOdoRST3t4v9W2My5W7dVKPJlYU18g4peMsaBL3ttRCm2Q0osERDK
AfsvtqIKDLBhfTX1Pox90vg08tBZ7pcCFidpX6JUTcX2L+CRF7ryb1xbVSwDeraCSwBHnsTSXS7+
gJN5TMS5fxyAsnBhUZjS4hASoWQIFkn90SnjlxLqjeqz2yl0BQbk5jSE8d0w/t3p5HPBMNDBr/6k
ScWPhzuR5PaO3BFUSl29KEusKLPvi6bHu5Cv0gLka8GINvPyKbW6CtwQ68YqRs4if7ATHCH25pgJ
iD1sLMsmw20pZ6fsiPTM+SCKjyg2uGVLKzX3PJ1gcQK+/8ULgsWHEsMjjjypIKSTxOhxSpGpgmdm
m0D8mSVQmfMJYOAQPOD9rH/sHtLIXq3dFY7cWcVJRQZnKPJtEmC0eckn75vkEq04JtEX4TNBJBzA
7MeEB0UYwPa+EngfJW2QnnyLdoFph3hedG8vvxMT8hlM4anic9py32qrF74jqbMzU7p7d2KiG+/t
6M8BAVPpgABAw8kgNuQyDMkq8L7nBMLpkC3lTn5IAjccastSy7zQGozrws2bAKEBy8xMcifD3qhA
yZZ8lTAa2bhLvfYKEcdNYjohIOgsRFXN7IkX6LfSpQHgu8TWpV4oBBRerOVzBrTWUl9fOwuSMRfb
0+b7/RnF/N/AQDDcQ4o6AlBTiwjQ3QCDwdpj1y5eGdbkih2B+/3yitcSDFZItNr8Iiasd6VCyIC4
Jtte4EEd63j62yjXUd7ot+iw7Fyv/WTOyASsTBYbkmy1Dj6ONmyeqSaZUITWwPW7O0lZPGv/Fyan
279gawfDJVK5NV2WAREnv1kgCyQPqIk0wY1OG4bMrrxKmOrxf3K1m1v3HhKPnPLGblRiuR48MeB6
QfzbYyupSE+Nh5MbStSWAmvWdpiKHVwVnMZEqNB8mNesVu3Mmi9cM1xJ33Jw1jsf1NyucVp4eLQe
NtUg5DKIQa6x57rg/+KV4Y/lg/fcf6vMLbyhSvVWN9Dt3wKPnJlxbSNdO/ArL1LDWbqQ0HsrpCGv
fob/705+vdXiK0PySASoJTWMNeoIkS7OJAcBiwl4w5xv9Aulstt8HmHZqI5OD9NfoNryFAKHWK71
ZDfnIXnE8Ky2VyToCcp2yWsYnHxaE/7mNhLFRS70wBBfwDMKYmaKh+H7MieLlSskdZp7oYh8VVEq
/Al2xAFyY4QCC9cHKBKuzoEvuUfbSbYKydDwYe8RK2aLP853z8jQlM7OInCEP6V0B32GNYlT4aGj
N603lGtdmG5BzxqXPJDuFSPq+bWAvdEVkFej3GXafsMghBPzhV/SirFcn/8TVz3j3rWNNV86qbbn
xS6D+QTG1a9kQUv/iDeWvNK2kQwkCL6cBsXeXcQp9ZUaD+bZ1S3XfgKCvwyv70VDqU7NLAlEXP5u
e1V8xCxDbLhOeufSyYSxUUgvyZ0s1FLTih8JYCs46ypj5rV9xnpJZZCLo6a0vPK42P76RKkr0OUv
b1WbsKVX+1DPkL5L7ZrmKTqzwJpK+dGFgmOxqKKYx+MFSb+18XAfv2RQB/cPn8NTa7F6DYkCt1xJ
fKSIAF6q4dCQzazwQagTUahDaVCgrBLTwkvZ1FfdszLFve2rqP8VzHbKVI0IhgzyCfU0VbtEg2NY
96/3/rwtrmwXnemxH0kVDkyf4qNOwll4PEsSBYVFmAGJuPZCtvlSHcp+hsCwAJHriFsQ7T9zXzsd
A7ayotvdaihiZdisMOCSWLhCUEx65uKJFchh1tk42oPjsu+BIQsI096ckyr0A4KvPVZz3AVvKOR5
JaxZ64z9cqo+2iIClbKHhMSMN47XGCJR4ZWncU8Qh6npH2Cd+/bV1mgpc2wf2SqqRknh5JdUDv/K
YCWKMiOUPZQPgJP2hp2A0VyhwNPXvtopvaJpHTtgSoY8mOwkKUUekLnYQthnyRX0C+68UojIGoz3
0MseEE2/oQDUyRiKS1CMfn/aR+VWPX7kjuA9oO5ZxXf3OyMNi8ddWShvAiBxqBALSZTCNTQ2QHW9
RDd+v0/eHUgYKX1k09dZK3q950m7icdc3y+GzKjbetiDb63BOKiTl5aCB2obUZPyDrZX2G5XwWVH
E3I2fs5E8zDDVGSXN1tCTA516c7NF8juUGLcuu8XPAiyCx8A9hcmkTumXnTfWr4pSAsADPVif24I
eBlJDfqtSxysCDvurc9VhSSYCvyiHqUDr5ShuXwqtmmDQ/J8cWj3kaSwYSU/1c1OxP5FTdsODE0R
8rvfS7ZHxh3uGAZzU1HbZbXARNtaC8MkZNnDX1xg44NR3rUSwl+P7eJ4JtOkNVIF70mOziAwS1TS
jQPqcjI6JuD1uDkYdw+N9BUza6WxznY+LfXUV2fUxXPU88Y8xmm6JCjXFoBlHhFMw5rBOUZIBWbG
+dairCPKCrKGg7ZUXpaewG3iE/n3P0iEb3L0B38+KL9iITxrV5OB7Wwx6aDVzDCz15SzSOJftFVh
jAaG7Fqy4m9kOVPaM0vbztdymBhG/bkPLxOleNH4lytaNQvASbe0GMwdICxnJuOvgo616GPR0gr7
CgeFrfFrepTn+lB5Zr7PdATjiPqmU1ovXs+gtdnBBHn1wE9FT2Xzzn+zdK1ZuwxGKDN1rfpIRFcE
+6vawB9w5Oc1SFJ2SsuHJWW3oYQGZPu/6QQIelJxLGNwB418oEfKqpvkTUahqTyglDcOyCIH7ZNq
hYDi1pcURoxR53XNQFc5qy7T9qXq2aPDixu1COXAWyh4BkISr0zYobNllTWqDGlE7GMG+DJpX6Lo
7I8rL1iSBjX+ONCEmDKmODMm6rktcxhNjlJTIyNSh3AA7/MJj3zcpTju/Kzhnz2Ij/0IfVEHFwiE
DE455l8qAs8EqVUVhhI/rxaLnc4ZrY/yJbTUDmnCpmUZ8cpiArkOo15X9T4rPYed7lWFtS6aov1k
ndqZZYsrlcklgyDiko2FFE0K2lfELLndNBaUGDJg2yn0NFdapsfMz8/arcYtqI+leCXWGjJMAsr4
vQ2eVEZZwLD+7OdVmfdUKRwz/p5mywzJ18KAPmblCHPl7qdvcJ5APWNKeMw1BMWo26LG2BZqKJOJ
SbbtWDWa6FKjQHSh5pPHyoSS/M6yi7xaYwk+we0sUy1tGNG2jHqbEv4pmGgaNQecTKtdqAr0E4BA
FqSD3wWexFszopgx085Jt3dW9/PLSsPNQ80VlUhPph6xPWKgeaxw1ZDHCXGnn7QSRHG0wQx0DV+/
w79tOxoDAlxRjWsCBtn6AXrvo1nTDCKIg2cjjKakLUlbW0xy+j4BMgbAfDmRpnTRhQL5q3oaCBhp
NHVQF72c9RL7EYTTEFBc1Sp3NXOa76sQuEDntbB7aYzJYe/Gl/B2NDM7dtOUDfU4vCyAvvwtdSYk
Kg/ZmxBhZqzLy7tP2IkP1cliOjrX7r758OCes3Jxn5U8q2pMqcBK76d8yKryL4ed6chHtDwm7pxg
vx6+MgGmUt0Tx6B33d1QOP9CVKy2urhzOA6j9K+PnoeCsLKJcdoq7EyWmRdoqI5Pl8M8F0xd0f+r
tgK08bcV6FHTnIWfQqEXQ9tgDFD9+FlAMitcM23xoZE3LO7oGh+u8lQDfR07gc+HR3vz4d0X2RUO
+4Gp6OctxrirVNjyHZ8YJc6kQMm7M/WS+qJBIJ5yhr3SAK4Gpx/caVTcUb759uQFR+hnqaU5ApC/
eAE0zRbOiS775TPWhjUKm0dggQ85onm37JKGXuBV9Ks9Z2emqPjR8MQ4fto5fUL/sly6OJF1ZNWL
u96GQsbD27ykMYVS7w/ZZS4ofj+NGhbCL+SYbAhmsWO+hxuRe2Fn17K4Kdt6lViBikp24bpkZQUT
3lKs1kFyQxEt8Lv6Tcq3zWMclj+yA045qW3y0RCLe2Ze6ejx/ldWJYt6p3Pu7RbCeU/TIvv7/EYv
aV2ce9OLN0+bHkCFDBkRkarSH6ESZ1Er5d1fsXXLdQAzIt3h0kN3+J7S1a+IeF5//6aZJepjS+zp
RAVTy6Q6eXLc5LnJY6tLAL4y0RpFWCTLqWzELGaDGtJG151exSOikC989uEWIQ/vrJs2y3K6p8da
+GIU+i3lUBpWq6rsfoLO/ek6F5Y3UYD1oI01/NCk3vlJMPIpuXIu+PQ1SLaX8PREeUPtxk6OqSD+
uxXOEQO1gfjVXmGbUgpFOEoGsTgnHt19MbGvfvaR2tYNf8zZvqo6I4FFIoUPcIPO2OKxEqpXN2Tg
7k4rHtptm0zlpqb/rLNH5z0Wy71vDhAIkNOpxf+infeFUBd2S4/ncHaVjeAAz2xk9ISYlk+75fN/
hNTx+LUcMMS6qYFLTchk9Ffdjf4kZKa3dDPivbd334Hm6swQL8ZQNyMOBo3S59iQa/curfyVTPyz
ixFtB/QePLqnNnYWESOLVRmXEASuH3Hz4bOK7R3FP+A+3RU61jGvvhu1Gk9ZjRlsRRHMa7BGrF/a
Iq6Bn3HPgksWEh4Wdr06g8riZJxqM8K1EZ4VUi+T0UhHlmGvi5VdCt4k7GnyENjst+TPVyGUOdc8
UFoskUgO6D1j6sOdgy5hRvaMJAL1R02q5Sa4L2SuzmvaRjVDv0D2arCMqcMROIdTBheJ9KQaUBrd
faxpXuzGIOCjWZgG3ANCjelOU9ECeNu7bGr37mPRzqjv8Cr+m/o65XhD6zETmQhuggt10ZRZIw/q
MASZlhSUnDiYQU8Eu6VUuUl3xRNm9mDS3cW6zWCksc59U4y/WLmYi2/BW62zHAOUkAfHpLsDSoyy
zd6YN9Z9uo8JCpHAfX57gAmGoWPh7619tvftWI+b+tR/n/qxBmE3Qzuztz+PPra7ULzo2fEhGB/H
MSUiAgHnfqTb/vCmDkgrTSfRrFY5ezALgiv7dIBdEgcj8XZIpK3Lye4zfXEUSYfKZW05VLvYC/G/
ArQ5HphUrRgDIG8BRA3ODnWm4KcTEXvrmYAkLAU/uw7hjsqDYTzbVY+X2ZmGaMQZmAlsj9TbeIVd
FWwv838H5pbm6TKECVy9aF/GYpETSDvS8fTXrUHxND0MMFev4GK3eKgrko/bRn0QA5LKRgrYrEUa
ETd9wq7YeEDF/Dc9HG4ik5A0jmFGzVR3TceYb1otnUENZAGyGeaWHRDwL/fwWk1cGKH7RxYMS1Rw
OkVtxXNVZo9/9jCm5RHvCJlyDaAxZECwu1TRG/o4NY+RKk8YFo19XWo9jmUb5SOrS4UpgTY8n/hq
HAkk+rpYutUo3jGqzC8ijSCZHDBWn3IJyrKUzt9q/XFUE8FBacYFjTUmOz7fZmlSAE0+bX7ofDUA
QXizLTsCQXg+fZ0qGeNE8/9mP0NTMijBcCICddUWu4q//2moVCQ6ox9JeywF7waweWpikEhaa4rL
2V8DSNX20DNhowcMQj5zWN7knIEgx5ensNWMZ4QFgihzO9YaSIutBtOLxblT6vWN/awpC9JfroK1
p3rwAXPK2Doa3cn1KdEDR4BGQFzMSDi+mqq/SIm8SRqX/+/039wzoYPVYFZrqfKdYIX3hayo0war
z78oAvZ+82vnPI5SyFMIUKQ0/NmJgWfF4FjDy5q1S21GA2pTTcbHY6hT08ogPn6RuSNrMTNNF2Iq
HSiX9QMXQWe+xwgBa/1ELnW604qUsvKTUzyMPZ9pNTUk++qyG+CHTv3tLBFzX1mTEgIQH8fR1Y9B
dWYiEBBgdGRmmQsrOsG4/HkYCpRMY/oYvGrohQEy5/yV4jk8oCr0U+I/odZLgzJ+TNmyfv4HEEQE
JYEYZpYvn9xPqLKPr0JFX/B1JjVJ2/RSZtICcHeKJw4VCDfi3SWzLnvvWldXQxFwXrCjSelHUsxF
KnMJdV8o46/S6tE3cjDaT8ocVucyq4KbH/7TKrZgBj1pbDc4KnerReW6pfPKj33wxLVoY93hiwx/
qt/4JTf+SiHswl/QsNjYmDMkKQLWq2louMOCswI5oMs747msdYEicnYmy8A36IMgd/vPbgcEV6TX
mieobu+8kWnVs9zaLG354yRgeySfMLLPRbDADfdk4MoVhLBicnC8dlG76ZII2vvdbZf0bOyFkezN
tPbUAWze6jhn0E6TxIVQhyKFfWuD+gmcuGZuZUaxrBJY2rX8hKuu112s1zDOwqZ3714G22vogPiI
ureH2+LklVb8HmWggZXKxyJXDEpJmVT/5pgbG3eoRXkPip9eX6IsZlbcq+wMzJprz0oPYvXiIIq4
4najVYtmSDCDTkf2Hzv+G2O1adxFjX6Q6oR4LTE97zMOH5WOG+IQzZUQwwR3Da+uxGSbmqJFS59O
T3tqE51hPHKlQNo8z/CbwWdH4aDmkEC8okMqMrvIMx1IrfhrxPczLxSDyhZFvXhH0S5BS2LqdRpK
RD+zWza4QDK2nH9OpUFSZHD0bLTbCqe4+nyHywYZ0tkQNGigkOQaeRtIff8Swaqem3IeolisiA5H
NbdpK3lVe/ZaY49g+BqHPsmKoDNUM+xWA85JffLEG0zm6RYfTDGRWGJyd0aw3fxbBzBoWwlwYbTR
rcyawZRm4YMGcJ981CXS5djooDghpxgIn4aya2QT6Phrc18ViNY5RoxelJfv+BO7RBrnxwGneS4H
fyIpiVn8BW3Ui1WEZOSSJSLND1+T/ttf1SstttTICFIsxhphv5sY2zsZZFeq9ql5BUvYY0+dDe9t
WUG0tByMkhTJigYsQJw4bm9rBW7e24VYo0paNqAdcFusG3cqWmfNwZljh29vNvhV2tZtNA1AEJ5o
+w54HyajrjHD8olejnJdP+jzi/9lJ+EX1qBPeXLUOOXV0ngFNdBiAdTBoYiKxd6/jgVxffnoE9dP
ZeHyZSTHertkQ18SJ3YT0LMztG/Vdiel9co1+UOOH6pRCJZeKjjhwZq1BmaGUQHjfoJn2/nix1wh
IW2GlBdR02ReXwdnMDidcSjUvrqQiQZULo84ADblwqfyJpBd6jyrzazdXWnN/9pXQ7xIW1rqQPcf
fr9sxABcdsIU0E965c2OH9cXSUluBUv3ncPVWu9FO4rpLZReSJNNnBBTEOu6O/Io3eRdWU5jJHOX
9fPpTh1U/B+uYII3seLXDMNI+qIXLbcBarUZ0JZjfNnFRH4wATcTHF65pInKvFh+jblgjKKbPXm/
fVzLogm0WcGu0KRjpTFby2m4IIlvIWqmRD0vj0A/r5Imh3yyyiQU7CfKhJTu2CD9mU9WBOnXLOZM
XzbXVwuIeUi5iaaiye2HGBBDLi4hhmlT6S9dOJJxmP8Q153gX1SM2X0B4bLU/S5QgEpcqA6Y9ikC
/Dxc0G6wXHCl3kzA/21ETOfrOk3HLgvorbLi9p8enpnskIzzj5BJeDNR2Jm62XNParKxub2tfyVQ
oJfnIEPzI8HBlvPBEph4TvM3gd5PiOTstQhcAPssJ+PUndyjeHICKgkvnPs3h0QiiwLpNrfJOh0G
U4KV6/y+U+G0+GfSD1p3TNdrXVtvRen7EAMebZTq3jER1dYPgZ26lcs3ME+A2GmtkB9grW/d+tJA
czq3y7UQPCrdE6FfRPEuv37moZ22bGC6Avp2zCtrExY9ksdYUvkjp5tfzbgORdEVMfK/izVGKzhr
UTi2Cy72uBzy4mX10Muq+60TrJBA9/KeVd+kO7dDb9UDmkpQKv5t62GipCkwFGudivVncjBK94xi
qMLAgVov98Bm4XlyEKyN4oFl+1ZtDhLhaLgnJsJCxBjaP242dfGktbhqfuNXtJo5oG62MtonFMID
BrD4cxmqugG3N+RReJv6rpwqpH4FL6h6kOcqnaoorrbLOEwIBKk20AUQkCCbO8lKDjHl+PKiW9YC
yR7S3XOlhcop2jZkrkHZ3+3bXLdEtRMt5DGFnmp9B/mq2+6B/SvbHx0SnPz3/MA33MA+eQ8o/249
Dsp2y79z5ko2Laf/70xcflLDocx0QIhiZDoNRvLICQMhOZd/TyiomOq9v/w5zzIuey5zH3jtCAge
kmkYNBQyhe8DT8D/SUZTxPqsfyHr+AjKNyrWs2AA00JEQ/YSAvh3rV1/pAnSFRz6gTSj1O/0a1zF
mwiPdcRK1vfi+cZ1/pxGoDFxfVSxulsWz9MX0BkiGQNHSkm5I2U2Bg6s9ud2ieRk8g+VsCQq9MHt
dw7VAO4ZVfJeBpzw2R1+V+Od7ZP2qpzydHqDUauv5YQIWwJhzY6QzvxiwHk1EIO1asp38yvuMOKj
f5R2a8o264Dj15km8O31qutKF13aVs1F4dvsr+8NCQ3qsR/nzmRttiHV9YocSE1EaOvCSjgqFedS
J6CZeE/rH9SRrXh1ANN9zhDSfBWPOjnNkJbbxZw8XY81MMZ771lM4bbSArq7ciCwmldR5J/VvQTP
NPsk948aPHmgCbOiqt1M0Mgcc0oycOsPM9vks9PF0F4IsBUX0mZl0esm0SocpcoXC87EnMnJsbvY
jl/+RYDiUjYas7XmqWyLHDMd95qemaEdJfiMhkw65t4d8uQHj05o+TN4D8uUc3A+taqDQWnd6vO3
E6zqswCxC5QdnzKj7xQdl+gvOhWjgnzEBLP11wAjph8FOp7S0l63lcxgo+GJQok+KWGvepFbqPSF
O0diqoTEzrnNc4d9xfJCdgRtEtb497TLmL2ePeuHWsbptjJjEmQ88biOeKYfw5QOgm9at5AJOVFZ
n0PBkFY+typ39UkYs3+k8PssZnysnlfjkM1wB2GO8XDud+nAheys/ueJCnLhN8WE6938e2f0pBVE
lacbBujOO0kvsV9DbDBrJTgXOk915ipAUzNJQNy6H67nzPD/q5HrrX2o5fKaYDzOytwkbpjr18oD
J5IHqr59c7YdY86glR/kRjvXR9K0CP0eF4tUuHSehM98DeCG3uTx7TYBjwDhKcykXVmt9PBj0XOE
00k94qENoM2jfC8tEonoAFF4sdSDYUtgzO6pM36YeQorNkSOBbEGxzjeLU0swWWNP9bHt+WCqxhp
Z2sX2eWc1oJKjI/wlGb6hE6mi/4yRL3Vo9GeKAFptkqQrCeIV6oAoJoBRENomvBvBPJxVjqLUkNC
p7wwIwmHmo2okg6lMIEEQPtbZWMWubWjkDixT2PsvWLs3KlWnvRnWP5Rj1X0GcCySma8hctRyOSU
dqx6B0T7ax2q/FOG6IrU9Np15r6SCjQx1lVTorK/FJtGq/KwNmVvqtv/wF8ysSiVxNQMGRkbaRYl
0agbCznbMR083dQQxPlqk3qQTeAj9wdacaoEniZMUqbyXfuUKPXBwMkwOoMNACAQk/4zeqt0slNJ
i+cinXSoLB7a2zfUnvKmxr4L+I0WM2gLeUD7NEUdq9H21JX0jjSc7Wah1zaXx9hg5/dGFs8ziE+9
F7wYYd0th5JNtMDA5dj2g6vgB8mJq7WVllBk4ImOw/ADoxTMHevQ+BI1+HG0TG2rdr1K5+DgzR5f
Fs1MphGyneGkGPjUBoFo+BPiTZ3YjTwsgiEjC9BZEA7H99rpO0iAwBkMeJoeGJi1OlGM6fNA5nEb
AP/+0r/K/4TuO6zux5AeAPAjooA8c1Zbasc+fXt1Jmem33/yJvuMbIFUqBu15aaxMeaXgW+p++cT
WyN/FiJFjTXIGxU7zv3SOGENx6WRf4wysnHyto3GmOqyS9wywDKyTOdKCqlvHNV7iAh6iuh/HgNs
pRVjvxkvKPjQFVOcp5yf3qo1fosMbABb+gnhKhKBqr9/u7h3r2Ye6t8+nOZPT/fpCuuWoxwDdNoF
uwVnojkxCLfXaaeQ0otpeG/ELYvTjqKKTi1K76t8Kd9EIQfRTh0rCEKabNXm5MWyELXOFR7ANaNE
TyurTqZUxHeJBFKhziND6CKhpC1CUowC64m4qDhM0rZV7GqIm02nGbXdHZYnM6U7ESEOPGb9NTPs
QoYFl6jliZGs/1yOiJQHILyzzUoBoviSsmNj6QR8DeLRPVn1JJyKZAWDZ4HCrH2S0MDNhiq7NRmn
fBYvg+8nyXshkPA/6pehk+gx4MNEVlbX1iVoGIzQVl0LknJTYa6NPmG6Vf3cLWp2sJgaL+Sx9lfr
DKC7TP9WLBRKNC0ZUt/Wrz0eLiMcQGHnb8esjavWMZ3izts1NBPUPXd1ucCToQKSJfluyQ4NTcTH
KUTFRoflukO1+cjOfShCQ0FKqGJLzUubqbeAZ6ITrsS5QyaOyjQdz2gxHEeJV/bPetytAtCPAt8W
eCXcs0aRaJFGMuqvdiN87ol3q5PQ3n5ndNVcFkh+5H8J0OH2cg7fXu5+TIca4aRxqlnISVOPP1Fv
dOZikK1wyOzyeUIaOnCKz3z0ah2QUeabcESlbPKRITXDCdHf33pxLLfhoY2oPh0tZ4//5n1gh6ok
dfTVuJca9R/qNx3cice0V4b6QjA3QiPIxXhgB4OdgPDDp0cj1uNXovmvQuB1FJiP1sNxMOeWK2JS
wRSlAUKwEKlG8lohHwNC6C1wqcxv3NGDbAUTlJaGHonkSGdWKQsAjdcOoV7NK63aMMHUMPw1oVfV
LX/Pndg2VFGE3D1hj8FTOSqYkRuw/n7a9KJbud1qZLXlU0Zw7wGvwxJcg28mq2xHPr3yDl+ouLMv
V3HkDzQXWk2J8112xhf6QJaGMkoD0+Gvwo1yACUm9er74xg2499ahjQNeJsQ8r2M7Zbf00FisVAa
czLG+vUR13o4mKS+0Rgpy02m9r07e6lDMF9g1aXL3vrk5pG5IciAogJ/ZA/u4XhaIartOdPnkgp/
mix95Z4xE1UeJbf6VB47/wh8INlA7vRiXAdDiwo5rTEuvSPs3AYK6Xxed0s5rjjJYEgdIgzFuAMZ
WvAjUBxsBamBjI0uAQi08bi1waq2XElxnTN/QbWwgD/SazzGRzaTDGpV9ZDIkNbaq335ll+Oz0IA
KUov5pvzORgXskM74sVbnzzPg6OdnppgF8B7gnEQFEL2RcwqXbjpqlCcnUcJzsubYAAb2Z4HosdD
BZd5IigYIM68lm+g9qjnjg5ZlnFv0+V01IEwy3YzHBm/WgbjQsVXTZa8dGYwrxwSxIl9ZwNXowkN
hdwoOYx30GkLlu/7kr8qaPqobIQt1+HnWufE1WTh4kwL9y0xzgBHuhlWNLnc2MvQXmV58QtULBBo
wyMdsiuBZXATG1q5aYIF2fYrlcqzfHUxEQM7/jy84a5DLCi6igAzWxYCwy1xXo+ykP8IIOzMXkI+
lHiWFda9soWXoeSyOu6IrIGCWgW0Upi3meQCUrOQVnwFudDBO3S0Ad5LfZcr8WzoE61PiPkueMSm
phCfnCVhn36GueVzq7N3d9wflmL79TZWmTMK4NTmoXWpVGB1GcwJf/8MLSU7BeqlsAYHnXHVDe8a
qxG7h4qF7svEbsrhs40FiT32I51YXDRzr5bTnno0BU3qkoV+5PuqqDOMiF+Id4rCiUAtMPakq81D
jWja+eBkkp8HLo1Em5iego+XjRaXidkWWo4JgGJA2PgWw/Pm+FGJbTMs/6muNr344fwTd2pxBcTX
45EDsdRBIlDa7cbw264uZozvHFVluHAWXif9ugV6y6OVg889ZivEz8gPNb9jPjvcFyb+CPC8jPT/
bAjV++eC5NAMKIp22rLWsnNcHIhfaVlhR1P3y9o1lZO4VZQ+qMm8TPvLimpFdw3iptM9zsWZ+0Sj
BDrdu4zRWVxIW6ImxoM4FK9Pa0/xKOSL83kI9IgdNykrBLSMo5NVg0DMrOSSxtDd4cNzrWD95+8a
Eo/j6y1EykT1rp7ZxsteLXFQgjWBUJ+fv2AwuhORU7kFcEfIZUedlCfxCOfG4TTslOu4uPjHYUz5
IEUDJ09PP8wRDvnRtMfpPXUNN8xnMNqrmJSqiYjhhhAtyhG6XAKfurgOzxcBzWQDso1fyeeTUNwW
gm3Blry24pX3oVJVObiNH73/bbwo81lV2JXvMujJdgqPhAIG/I9Jyf0kgIH03frFfitUZ8GCTPPg
Kse1KTi1wTtsiTBt45huIDBbBxFxgtaoWpP7Ah3lV9gkURxPtW55U+16f+AldLDIFxbnZL2/jBTB
AvLD8asdvr37phHMQDqYTi64XKsl/MP2REVgmyNxyLk2UqjdCBMsmhRmzNh+IDI1ok4QsXGcRFOf
32giV9dw1+rnRn3AfWWe4lehojMM6+zhYUP4B8LGzUwgsAw729yUbJOR+/FZRAxC0RwgdF7kDGzI
H5xMU20CilDnY2HRTH2FR5P8EPZORfqVKnt/gvwDH1xa/gAZzLrIJiiIufqGdIT1TCqJsBqr6Iv4
sNzT4iSRuwNTx2psHCgADoODETdNfqDAjnN+uc3qyrkmrIodt8iiGEpqAx+Q9lDF5voMaA2O7g5h
5Te528HHrJgEQKQh5RiLVovGKJ2uqF0ux4+B32ch9tQEv4MBP/X+j013f5XQE+sy0OzdVMcdx8IR
e1m0AYa4WJt1ezhTG+n6x3rRjV6MnZuXBjkxXlQQJUBWUpy85j1YPiXz38PoeEP0BbI1R/S5mgR+
Oq+teiQD95YJrvUwZGWKGGoFIpRB/J2zAzCz2douHKFtGBM1/EPv4Cj9Gd5y95xyCpbpc6k81FLa
nYvN2gnrKvQfCRzdimBMPurF5kxEd/lqlnl2kjBOht7x7Tqe+3xNia+IPSjMntkSzH5WQasmJHpb
XyijbHuMvVonSa5ScG2xzQScO3oNCrCTr/bAnaZkr+wftutTOiZXG3eqTtvpVP+eIJ2aSorRuNX7
Zv+En5H/a1jW5ChYGJrNiYK9TV3GB8Zk3p99Wlvunk2erdgTs2nAenHoNc0PbnQv456789uPSm+h
MFF8wsK2c69UwQ7qSINU5+IoL7HEiLzJ/e2ohRvS9zGtFSxgfr8zC2xf3Es3N37/PspAbOhzOGAW
Dv45pcYsbLAQMHET88QTdUG5p9bV/XdGXdevEpw+cyifC5H1A8vo6iiw8kw7vEjoyxilRSb6eacA
GPeQ6q379Zy4+8lkt8qu2O9mIMQsTa8+rKpi1iOiPZ5fx4ZqRPJTbsgJ2kdp9Sr30Zp6QrMP5rMO
EAK1zpRTX8F9ld9OXBkvFnDw8P4kvQGfCdOLeJ27DDhAyjwjCwNAlS4hcuVOEapcG/MoDRWXx6Bi
U5qB24gL/YkZ2wvOi414R5bjj5xO2Pt86cQsm2m6OsmwfptQUV7OqH2LGaR2Sz7NvmSENZfIY1yq
XzlzFYwouSKnYtD57BPZ3+Ofxex3awN1h2zkAAfhzrUSKLZUbLUqxdw/JlDvVPn+F6tskZO6G4qr
59pqq6HbOuMaez7PATxuI63zR53d734bQ9Hq+ojbdVTEORyDFCBUzWozFkhzTlPecutWYVs1aapo
9GjJM/NZ5Jy/EgzIZDYqHBtTEwxkfHXJZrxH2Vlh1C5GRCefdFt6E8Z1L31Khp0++94LeiIKRcgF
1ZMxP+ukC0eODxAAYaiUFt2QH5da31RJi7Wt5k0zehJi7oWk8Ri/rb3+0iiGaeqiKe3Rd9g+OhrI
drzgKzAZyQf2hHPPUDq3Bs9xU/q1uLqzv2XodyEIHCF4/2+YVrD0fu+5svIqBGmwtCXaz7fqrtd4
T0KrA+1vD4cSr6JeitMWfSxFYyCZqj6w4PH+vyhqFplUtMq2J4i5bQ8xdfvgVOX8RJbSfQGuwHrA
jr0w9HuOySbpmnMEb/3Yn6mbnwv3gzZtjyVV7PbpyG0ddtFFq8Z+gJbY2BCC0INUaCzaur4Q2Amx
/ZOhNrJ1f2b3dGxacuKRu2qq02vYDzXsZ3VYIqqaL7nZITWYZP/4Qc2B4HDT2wMFoAg4vIARDSvw
hkdl+nQr4lfuOH8g3oDxiu8S48DiHP67EjmDOTZfo1SliCXJ8B8B2v+j/GmjpvqUnFdP6SAQdI0T
3jy/9UeHtywPn+LQ1TpTol0uMisKj/PAeXp3w+q2yyIt1EqvILjbnI1C/rOhlLTWzqKPJQLFZHKW
4vazIv1Z28G6sYMinazyt8uG811mftlgV/T+edd+rfQb6Uqdevj+krl9JHLzC81Wcnq4OguzYQcX
fu/lVHGxtkSqHBaJ9haD3nFJj2L2O7Cxh/34AYr7FclnicAC2xaqOMfy2jQvsVUsvxRjzWKVCPt8
RopSvu88ONdZPQO7kqMpVngPjxRuuwoTVAwyi6LkNZ/LztC3l0sio8i+CQ9M2L8siNmeoLJCejdb
DFKX3OjAnduZxlMdgIQyCVVm48oyJPimbxy2ZV392boZ2pw4k5cMsfvrb+5hQBXGIy4OSj0as/cB
udJw/1xhXni6PcnR99uy6DbTclVSG6nIHcKqo6xXrG4VBms/amAhiLOHFqAHbCuIKSUFHA08+stW
V+Bi99aYygfEIjLSdDZ4BKgVAz1K57nNgD6ffDuayGuIJeYqiBuiXgPBpdPDxAvVfwj0KEyxP4WA
PqRXBqwwii2EmWuhZOovyr1UM/IKyqbYIO/eG4xG4YO0MvAtg6T6u/J3mJQ010GzQHwd/648GmI6
OeGtspVkqZIIMV5GRRLeydVA2Kdj6oKNQmWEAz4nDb5ZwW6pcHlPrwrJsMs1cvPlSmv+9ae/nyYq
FyxS716kqz5+eZ9/V9PTRlFD8N4UfMB2uiPcJxnoiDD7vXOJ1XDNRMYIxBngVt2sTnlELINC2dvf
FDvpQM/9DCnZg3rGldtk7lXJWakLfY/CW+zUUEqLU0OOssxlAGKpgK2gUU3mIZ5CeSAPzmbuK5c2
gJpmD770oy4fgPkpE516nGXzdQyK3P2aQkgOTp70UgyvWohbGnc8mWNdMxJHiLYiOKwuqR/3GaPc
Dir+T42nwmmHLytG67XcZklcx2+oYE8sbRku4TQpx/58Eeq9aTMkm5ngPkK/T4FtV8nGFbRkWbf9
lknANZdXWhT7343OtmvUaUB7ybP2UJNXoXLdBc3VeQR0jguI2KB2nFljhkjafZkqFIi/O/icNicQ
Tf9Egc1SUh/aiTPAq+qeF3ZCjwnrvRfm91D1JHhEO8ZUi+1L1NFwlmCxjB6J7Z5V2AuYl/VLMir4
0LpaxXjmUuch9TMjjW3zxXlsDHWLUKtEGRCpi3/OELHQWeK6PoD3Pr+c/GViZL+0tyRAP4Yk+TQ5
tGghd2QLRy12Jd13zNAcLtygZE9BYFpNHJLY1EkpISJ4nrLh0rBEId1iwgaTDA8ILaqT5kbqIzYT
WvRiOTfl7vPuzvSNymzHwQMgNZ3uYGLcKeo5x2qSJL22Bbfa8gwrjYWcypA7/FT8vRpCQ8Xk27Pl
NyZMn9TDpahIExnb2tkq58idiSc9IUlVVb38kAsyjbTcL8cVkQoNU6Qq+jFclLSEpJesGGiZAX9Y
6P6SYLBdTFDwYHhCvMnYB5wchHT/aO76/LSaf/7skE51DcxN3GoQzjk+yZuLg0wqqky/V3KaD/Lr
gJgylFMl+x+8Y6WCfuOHLsMYMU4tbh6YGqpGDbvacFhj1efNWoTbPhZN08er0VEX3hZCwgtMczYy
JIXC4KEBy/QTjdfPoPKmFWu45IjDh+7vy1qTLT8Id0aco4W60ZunxKg0o8YKVY51egMdPkHQUnj0
ZSvJJZQ7nkHi2z/EbnJjkRCz+cMD0NU308kdpCVlrfdjllf55c/qFK32TGbQHbb5uZuDEkfGJh+E
xMsvFzyWYTAdpX3+YlUbsJu2XGhefZDmsD85q06VS6W1bzGB1fbCtahhsXAK6XyuVQIcd3cWklK6
PJnkkx+YVjucHj+fgVX/zQ2PWzpkK+rIEorS3UJOM+ajVYF/pmH71BsQxdQ7t0lQSjSP6pPTuAdm
aKUhlpmAR9GBKueLfGQb2gBoTBYM5G+PXYoR5HW8G9FiBeSspRq3G+0UPgeTV6JgB3Tx1ISHrfrp
ux/7usa1vm/muANVsXypXWC9N3mdTA3+4veQb0x2S8bXf1wdsYPBcHKqqcQZBybxIupnmyLslcEN
EMdYR0OSLeIioERtsTdxDfkf/VlQW+CuKUd+/IXG+Z/0ikM5PA3kB3X302QduqQM8kkLOY3LQyqQ
FanPqrSTl6S/2nBxlRwkp2JxlfJ78rb6R8TogKdyWUgUfLYQgPGz0REBH1awgO9Bd/kEGijK4fk7
a25WBXhPlwU7vRMI+A8MYB7VXB08IkARtaTtQUvo3zv9G4/bkhuscOUZ+82rZZgtPTLZYMNiwclc
A+HTkhB1Y9z2iykFn83zu3yHSdwHGVDpiyBW8y4jaz8+UHrWMUkH+bl87SBiC0gwgARV372RK+GO
wAgs7yorXDXZmer79NnOYN2dvvW04qf9d3kCkJE7SIC0zXGS8RW2qMlU1loFhnuhHYCB9Ez/j9Pm
HAXYYGkfwDigaF1K7U2A+KWNhhRZhqZH2Qc0nV6U51vyOHWh0NZMk6IShRJUj3UqBaphM41Y2Enn
LjWrdQ27Ekv4zxAuOsv535i5SK9VyASug9+wSWVY8IuOeeYgi2upZLHhtk4FyEVBuZIbOZKnav67
a80NIfsVxomA1Lx1xbF1ZN3g5lLzHfccjWosMSgW0lUPrP8iR4SrXWVFgor+aBxp2h5WdMwtH599
QuHgTcpn5uc3fNqFKi1v+tCOFho7gCu2uX85jeWJa5HlacUmIPFC0B8W8NDr4k4fBdgXY8j/+Z1a
Rr892XCMHBGLka4LfU88OK0HwijDTL9rn6MZWAsQNb67kbkPYOwC8Yn/yOwLusji6exVxg8cAmox
CGIIWGL4YVNq0rZ37UafkB9WygM6qKgYzvCbeQa14phSdwbcf9BP0Zs30LsIskge2uUJFSzJ2+XU
o7tM4jhakzeF3g6qMu3CM7PuWmoIQzGp1CT2BQ78D1rmsv/ObnAQETWva2E4PJ46PFvDRj7ZyA6x
dyHmBUPgZNAUWLezH684DevHJ0bU/2EjEuGQNFXcA/U+mV4KOVL4h+gYvY285M6ygGoatWa3R26b
Xt4p0Vh5CbF5i5KT8wCuGSZrhSe+iX9BQHdeJkaJ7Tm0FYlNNX/d52s1EoVubwHgJed5hq0Yl7Fy
n46h+Brnt1y9B54jI9gBTc2Xz57nl24TQr+lBawBou8rHkphoyOF5AhkIek8dELBrIa5Dy91SZTy
/JRG7meH+Piivwx/Qy4E8TDyD3L2DYRPsCUskrtWLzST390TPcNDUKxjtpqaO2AK8YvtEXS0ORJI
soAjzZRsHlO4GjrDVD0SZ55CvhbPlcqmpD1wfDllfPgj9BNnYymZANH2OOU2nWCtOfdBN6CpScoH
bwX/k7zRGNvzTemxKUic4RduIabsRUU4mYL/cKwa+Xk0gZaiJjSRvtcq2Jdq5ELEwS1F1vV+zney
Q215vlyuOQ6LIGf2nvqZ48u1QYYIKq9Cd6lF8hALV1PFeiyCICPf0LZ1PLjcLO9HlX74rvOA0LNx
bJEyI8/E7FrujhaUz969bVOimiTiP7D0NFibpN3zgiUsd2HnZUuhzVwk4vOFGJ0FtpN6La85vubq
iT35ImjTGw0U2hdJUjGlgfzWPFMOwfy9Rc5FDqTmYtVqdbFAPaJM3UxJF+QGe+cI2GROP7OrC+PC
b2WlREjdAXFF+3jWiP4+jODhnIlfQ2IO1lQ3GQaAb+ovRE+YaR5xwQL250hcv8Mzvx5S7i6EYFed
/Eg9AfiB8I0Ri2aTMwUUrNNr2zCiJnVEtQlRr0V9tUhUlNxE3fNkdTri8HrDtHmvRjKxOwhS9Nqm
jBo1q+WKLResnZxia6mEvjK6OecqyC6xjdRrhw6LonHuHaWDEgrMNucb3omgUadtXXIGbNt3xVBJ
n22K/QJgMD7fDTdwLfLTbtYYpNUKQWK4QA1g3B03NU1iSRKX1TySEVBHAwBNlIIB1u0CTE8o+Rja
UzqSZonrsYZ5yykTpg55NNKRivckBddsfpDZMkzifZo0zXoewYq8bdtfmYHErk/p0yL0eY0pDuEU
0W8/dQwmwcrWC4EwgDiS88GlEQoCxpwH97xt9RaPf400jYtS6HdeXAim0WmnSHfaeRpBFw2iLHNr
edkJ+jslQZOp6OqONtYJqphzNM3Q5WrO0wgFZeEqnvnSgIjTCT9ZmfYSgP743AsiAqegREAGrxBQ
Ulme3xjc8K2uYG3MybOt9bvztAT+m3IZCLWB6w1w6FTLNnjGWv0qmuwSG9q3JVXXl0oA6rjIhsYM
1AwAJmC9KbozmjzUCK4U3iMmk+uvUGppPfjoQT0DFtaeEcAl0AkOidaasBN3pbgc7SKJrfU2+ToM
XRYkpL0f9w1RvEIxD3q/d4GB93kfTlr/Cdy4tqXoNN3rZB1jH3woMAG0RXi0ZlOuhZLAmZ+fjzfm
fHo7r4KHNiBqrlC42C6UFifAmCvyuoI1WcS8uo6XBapVDNTfsF6IkSzL7BB/AaeVlyari5SeX+Pg
RAnO5JDOrjbOEckDFkqY4qVSqpTouOUNTCXKPTf4t4KJdUqTM6CXIYMesU4S4PR+VPGJ2YSS1obo
p/pwdVpnGicksu9tgxGqItljE9+DzlXAPC2OkoBMMy9jzylnFkPgJAxuxr/BqNrJHB8eqVad3UEw
B6H17KAaylhxhnPqGVh3LHQD5RruHv4eM5gxk1bhse3cngFMhKFqLG+kShXTob1DmqEBp0vM0A3j
A7CM89LoY2RBhUsJhCPBkHb5U/91nmkpNxSbmYpsM7YeU98sU5Pd1mMxH+jn0PHEKKTZPOZga9qN
VReqsK2t6ckUA3t/fdSrX5b8Vp4uFftkMIlXx66mXE2ZWW4f5BGVJCSaR5QEis80YQuH+r4tzR4s
kBuUD+MfSn/eVpSUAXOwbdhc/z2NjiwU81Gl0KQNuVreEeHnqdLtwGIn0eGUSY/rslEW4uPYffNq
v/sTh+vhVoS4TZ1g3kF/FmwfMTguwXx0y6DkoPznCGCO8ZC3RWxLcuHSNm0lXp03IQHnLRhDkJFY
vUAGgTw/jZqFXC8NB1SH8ogM88l+VfctYLwe7xjf4UlU7VgoG63ZnYVCPVk8e3lbRcDjhUCJ8NRq
pMkWdEKCYA2rBHYkpKc1UInbVRynJ4bQUET1pwVndxxc+4Ge4cnLs/w/lc8LoE5ssvjsZWM/9bqw
fBhurkOiJAFTUmSJUtX/+YMd5McbOB47ceKXQBKOdKYkWIFe3wPo4YUcni9trhl9wBUW0kDW/AcH
gm1VaVQR/YQInORswNg/UV82tMnCrBC+AZUFYmuUZoBI6NuwbEYDqtNNydljRMTMtGwl3GWziFIJ
vInHLL/UYwRebqI1AMEaj4k8F5pqyevME9uGkrMGzlSJcLawV41KimFEzWBNgV/2PASg5WQah7qr
emgd70qQnBum0tTRFnjbh7IxzoWCg3/MDih3Fb3gfYqEhPUq3YpxNr6RgwDVePz2DqlRYm/vfQni
bnF2f+AuztUfO0Eh6cSSXM7FfFF58ASszZABCWzCBkimxxVKUVPJW3yJqJzOPw8/Uin+N4yg3ZPD
JcB3+1GDjwf1ANRrdqPoORyPxNFt/8nDp6BCr1mxt9G/Kq8kIqKTCYBciVOdeGveu/PysyWSfLtY
s8uVa2gRBg+hwwVxlKLHP8rCOLqsrRXI8A2J9tF1ybsPAuudUWtj461SqKiyc241mAz8z8qfMMl1
C8zHRf44bL3c/KZKkF+pfuzJn18Qylhiz8gN+w+c6+gQQT6n/BIwpu5dha95ydJDGXecU8tfb4yt
ANuLp75lexT1yqM+88bx0Fv+9IPYb6z0VY6CJMtiA9BOUdP5p8byAchnEM8aNkt+dSNikxJlaKin
qkfdoIHRQxPagWXUYfx+ZQBOYSyYqhypgpy4lQyH6pl3dhNytDaZZDt0oGUeH8qUse/62uTVezEq
6izBiiM8h/rtEc3T2/JvQ8bVn0/kjy7uod2CFwbjTc+Ear3aNuRqd6BRp+UMvfEZgrifVUZemJ+r
vDKGsZnetlPA98q5cHj/JMSBRHsIbYOSXbsgR3oc0QRqFQ+rMhQNcP8QsVGTBrwTFLEFK/lzVF6c
BzzJEGi/lv/iPxzSu6FQmmAdl6DamfHPJCK3EVyISnCuIMCdTkhieEaabqL5cHVHeKDqIkNfZbrz
SdBiefRtIkdbi0MvBeHKOEw8Ina77ofiXwZf+z90CC61YJz4kqbtGCGS/C3rCB+hViA7Q545vQCD
JkW15EhGK8pHKWhBAXJkW2hzWoDvW4ZF0DmvuycsznzbY1yhz7owa/nv/6pW8mQlE91C0F164ecn
/jTcHXa8Kfxi0DnFNvE53XzeguiIGMoxbVndPFKb1W5xo7BkloGc6eQcMfhoYuULXGPLTUzJ2xHr
lTgYjYodCO8HxSlJp3b6COV4WfVgC2pdo5RGKGMqYuEtHpy6gCCUKOmEABBwWxwAg3SfVyLWK+UA
7FaSJgfmG6UlVvFMTq5zuOoK8EAB0FAaqWCHjkHjOHKE/+21D5lySliRgCfZ+CGiyMKznimDWV8z
HS1Mf2gZ1GlcDsSsOpfNUX1XtlxHmpwHIzvrrewy02RGMg8GLUwbOnrkpu36yNe4qETyLK+lupl2
r7BdERyuzplDiwbrbuciy7cTshBJ9G7gzKMlXfCr5WPToJRWaWCZVfru+dzl27VoW1HI5yg1g+Vd
OG5TE8ayoBLHt9s+kO/2NKi/4HgXfiPAoBYQpvIYuY1GIenVgMN6VA2I6qfHPci0wwSU4TmuVUoZ
kcK90UzUkxD97+AEBqqQl/+t+FVViaPBQL3K42fFgfKeobgrtGGUNpUdt/oJ7NgUuRglHvfH+Znl
68eLEUaswCUA8vYyls9TruAqIt5jU+bcVuHaL047EaxXkiS9McgzBOiItecjMpWjQ6myH0Kh0wTY
2X+WP+hM6d9+96CZWdblmf1I5ETM4Qoov7sutNM3e4Knk3eW43rwybOg+5P57LO8hVbd33QHeZJs
IqjmhKARN99ECMt+6yvtRa1rgHpnaI9eQTApsv4FbMJo7/TQ99JlSsc1NdmUhC3SQSYP1Wi0RL83
Uk/jWiZsp1MPZvOQC6oeh7mbEwtynOiNRPX1lPXS2/yGp1xJ67J1RQQwnYwDmnAR7z/RSTiUgaHh
bFMW+C2kk9cfDlv2obSDySkK59PrYzBXXxzQlBpscJRqFgT63ajAZFVszjCoII6EkVjlsOMPfmro
HYbpyZCbcbcO+Y+uWTnN7oGy5l18Rs0sboncK9ak2mGDo5aRZHSKhs0vroeTWdZ3eby0tyUdsLgq
c402Tv7wi20n6sV9f1EYHACU2BrHF62NdgV5VnOpTgyqgLHsq2vVXzW61WwKLFwOE/9FlTlsyGIH
aS6jeapntCfqt3KoRL2rRi0oBkrBRd4AyqUvGBDQW7ANqDcPJpPmCQdqHSfDDvV/sNMvdcB9/BI/
3jRza6ez+F1f33mqu2fEihL9ojk9ZSpalFF6u4bNztBnZGJYHOYS6yCSXoqi/RTmXr25bvUC1tmB
ImvC4239vwvoJWyU5dzfXfMkxlfT12FFbsjk7/igRgonXqM1MMnpzCjiCvlw057LZ584fCO/RTSH
drA7DBODr5Pf409M/jkzumEMpGhjfn3xFegxhOm2JG1Isspww3gRjTknkMuoH20kxAacEjniM8Pu
7qvr75UU3rpx92YHjfBu7WbGO4m/odUMtWqTvtzUrluE8wwSpB1ojsCK9CrEN4/TTP09LVsb0FWC
yXIjij0VrHIlCoZ/a4HKfGcmX0TT4NWi2Ui02CSRwvuM76DAQKVbFgx7pOUSA4VUk0ric01yZKY1
Bk0isQ6tCS0xRs9gYOXppJfKS0FOPRnUWt1NMZJdLz8ZdHBaGB7xBTfQpYWD1xa7+9F13luCSdwr
KsKHJoffDlIODkAjv8YI3+45KgqazTLEkV+av2TRI0oL4O4960uIKcJVtMC7Cvv5Yy2ycPbzJWir
CtqdjqdWPZzXbCL1D6Z8/DhQIziuNPBlzHEZZghaM9Hw9TzqVsJA/YpMZoZh3i02LQmF1zBQ87nO
1/2o4Eht6YtikkTfFvhRa3VZy70HC/6kflQOIlM1S1pmhwu9l/DTuLdJCppOMkUqBcTslu8ww4zA
yXe0v6Q55zfk4xSAv/cJYMSZ+3FVlxX3RkMCGEG6KDZoymwnC8MTqmzx53GtRdh6v2YZdPFJI/B3
RVGFRsbHTvXQdyzZnj1RxqOKeSi8S5ZlVd3d9vWy1e4mx6DKsrvebbcF4E4nJVU+zQZZrSRgwjem
YAO2kSMRvl3Hl34+YMJj1fUeH1DYj86P4WKl8VHdTJsbGkjvQmfVBnRUY/7HPqM0AVea1zA/PHbR
ZMlZN5UvUGxpp3fuebyHHhy/BqncHd8fYOeIBMzLCuloCob4/7ESp/Sb+PiplOCxh1Kq+HAJdZwG
osJJBxs9/OgRcOGzqK3n1KFwL8sW7YqS2uejeVKOmev9KRJu+mkqMucpATtkXuwuZ1s/EBLmuxiX
/ffcQv8RESdCHP7jWVJ67Uz5BfASSq8n5d54wIVEtVONCWt3HV1NQ4CMz93EFNxRnsmWj0rbnezC
yWqll46fgtExFKooFR2XgkEoxLCuSY2gM2WliH7AFyLOMWv4rjI9trRxoi6Ti2IaNDn6RKyiZP2k
jTNFAEkQDWu7wkMV53nyrK/7PvpXx+GgVvP8hUBMyJKC1uIcjjkclHsz7emZAEZniyw5Vol8pVkl
dhBemU6+0/wSaIANFdf11JAO6hJFtF/ZkAgxWuJ0s93c3k2Hc/1EIXgue2PC7Y07mj8aMBIm5dnm
SwZG8A4gQSoAhLSw79MedUndMWqvsNlNqmW6+MGslgYqRuXy3ovCOoU7GyNBbtBSuj2YCV/cRRlK
7PWS3a5CIQY6P0OxZ6xgBYN0jJOzknM0Arm7XS91+wNp3XWvcEY2eLcqwDsKLaoqS7+FdmZEQNPm
orMm2uKrVXNO3oDYAqCDRpbrDrnOCnS4BJ2VhbfBKLjTt5fytMP7BmwyxbRmYtiOb4rn80HpzXiS
t9InPJcpeSFcVr//1SsuLXh52gQSLB58dYlbTEecVF3gbfPGpuXbAGPUSeqXhdaF7lnVvz8lHSst
TaScwvKd9ARtwdhjZFloOeJgw9CaKli/NCpQe04KJXeM+LFPtYedlBTFeXLPPnIoU0kan1nP8WO9
sGL4jpRWOFtaQ4Vl1L10zJpnj8sMZE+pwIa3Xe2bwGQQ3m5bVud3beStbeCISOaz7oogj5epuQBS
ltjNa0CpT13/IFVx168w2GfY73Q5qVesTlyMsKZtQ2x22iwm8j5mUDY2FfY7SXntBgC+1b95NYpX
YcicO6xGjS9FEgJPXYsf+5AzRop4IMnMEAwL0mZ1/QeIgqix7rmP2WdsOP3w+A4BFqb0g9qkk0Ck
r6VK8VR5Vn/U9W8XawYz1rmn58iliQR01BaG21AU2Y59yMrwRjhzYDTdJNtVM6g6nX/wxXnJpHTn
OX2XeDGOpDTsjm0MB+pxJLqzaELcEyoktA4or+6IINT3Tfl9LoTryraqoqtf06Se9/IfIF9o4C6/
TIuwIXHHUqTHZ86ylpu9/lob/FFSKB/Ci4S8EGAXq7j5zZWt0A1JO5qw7xUBo76zSBBJaufJ1c54
cBD89J0huEUxNfuxtLXWxgjEugaLRtnlfWm+kNuY+849jpVaiZw6dw94pYaoA3wqogbFT5hcxbIU
0sOx2ad4q2QEosDtrcRydShwYRhtFTt7/fXaAwTMlKStXxzy9YobU+tAoQ/K4HF3WW5y5HdMB2//
wqTOFxR2oD2WUA5I+nDIaRBZf/d0VXc9Au3GyTdTHVYLoRZA0BMX2SqiX9QgyxHz7E4AJYDB7c2C
YV5vWLrtLIjEhXMv6vYL0vUn/+gWpSpMuF9CdQma5EaCMo9JNzFsJ7OJ4mpUFOH+tDmzz3cCG6UM
Bv4mBWSuYl+8KgNaD7Pzkkj5kPJV2hvJXbbjmCd3Yw2d4po4idZt0S4CCpGhI0l+ABkMlcrbd44o
5p6Mq0aQjaoJaZFHAzQ/cVdcHRzLjxZFBYH9Dy5c+p12HYSFIGFpUOLPHEdv3rCBdDz8anCME+Sc
tc9FQ1q1cFDcJqID9plRwsO2peUp54tyR9vdwFO+qGwv8CmuZHeJacJ7S4lTARrY09lxu/7Stfdd
QtKQBFY/HiWjmYUQBpfA7fu+gIkBRO+JO5JA0VaCZfskNSYGB1bkXVHemusbvBoRtvxzLiR+pw71
xCpuWYMeup9k9PpH6G2/t1NRrKcrs8nEmRMuOYI8bVpUaCs47jprJPmVM2ug93nPYEecF2ljTlLR
YNeuNYAfUljYEDBbOZUY1T/vTY9rTt08uH3bxvI76ZZOMToim+qctyj818IgdX+GG7GtbLtxqaUg
i0nDvPf5Zmqz2H/0UuJlCTX+V7kfJWQ0xTQz9TlOgWj+/gquFo1Naz2qJ/VlYV4WnCCSb5rShiu2
x3t0hqzFiFlq8en3WAnQ9I7OH43b92ZjrpOiGgmSqlcajZfa6cOmq+NgDCeq76smLS/wqs2IhGns
t6/NE7MLk6TxCqRkFvSpY2xJ0WTzZZItl3u/YsfacRSoUBYGlRtTDh64aeGiRUFFFXWa9c6dGQiD
8Tezd48oXPyQfGkFKYOnuYonGSfDSW6MMIdgIAbkh/9IwoM6gEvebbSGFwA7HVWhWpQJEG0VjJd7
cs4NwiqPQEfw4UvGL0C6kf3kNTj4IP24YUxGtArJNexrh3po0EojfpCXtrN/LhB/IwOoE4YsBvTs
Dcviao0WUEA1aJju9P1WQ9WEh8lYTK4jcIzn4AIoYDn43nEwWrKQZ6xGb7tT++aU/b1VAfOr3m4S
Kf8ZNvfDUumLRED1rbB6Axi0+eXaQASDRgzJ1AiL4O5FKz1MsklEjwvXRzOZiMw4nW+4A5JeiNY1
k81DSHLZshH2VB/FobIrBfRbHl/Rv6svMuC5Y34PlBkE0CbzHyRl4DDFlDkZByg3YyKDWBIvj4TZ
LrV1SABl7joLuAmsC3/Dop0D7eMkePKN+Sod1fmNBXbiW1mSNlMlINnLjoMHTN1SyVVGbS1Y6zDX
oaJwreJVzPs/AeOcEvxEUPiz6X3HNpNlS/1CHGKKz5oTLP8aObgVSoTmkdRlnoyy7+4ZFQMIzDEU
obVgv2Vi9GUJ/4gTbkk3PHRR0dtoyWgYf/rAknIkpV4jJWsmGD5GetlUYT95skmWScuoKxjmwN4J
rbuTTxMfulnrBofZ+vK3ka5Xm5MOuRXvvP81PMPzZ11CiuV6MX3Lxsd4duVic1Qpe0gbNmKGp4mR
r52V30f7hr9GMHsWyyKL4ABtJ0x9rYCpbHjwo6/IZnReW+KDUNg4OzmlYzqXdJxSwnhs8zfe67dI
FIfEdIbJlWuGwpcV7UD1oA7SoyiyqjYdfakHW+f8bOqW9COc/Z4a4K7S7Y5TafloTGFnC81xzPcR
b2pit6YkYZ6MJqOmqv5AUDh6HLoGN6Q/Hj0kM2BooTAc0sVP/un/00QLhFELj1riZbvdg2GvjoRG
ueUya3OF8xAgzcBvbz1B+CNsf2VpOGX64U0O09kkVXSOBNurkd+3l3Ktym2nOzZ1jX9YPKlOBNx3
y27huNae7WQ5WwEfQvIynzHWq2mmlTFR586Ln19qJKhtuATRJ8sv+SLgbnIjGAR/6utM/UBz6zKF
XTt3xhGNTPqze58cC6zo+JHD4sG5GGIT3Q4K61g6480gSCjV3MCoxfZ4rdzee8PnEsTI0qOUH3+Z
YAflMrtbColTwcN3uxIvo18zYiwygraZTaxjY0tPvVrR8Shl2t8l4MK0wz8njkNCtQe9Pug5hD4W
HoTIHfAYstsWjjEZt/u2wFEclE5WOwsU0eVIMT/PJJ7dO5+9vSueNhVCMRkR0ZhTN8vwADEkX1fr
OkCMgwn3fcfQ5IMRYTFMsH21na+A5BEO1mPusDf3tNLBaU96Y1zNgCXm95w3wSwOHn06gP61OdqR
n3oDFiYm8VExf4TuIx3p9me+D3X2EACk0LnvUQkGA1MaRptMw469f5ViIuITPbJ3WSDkIrbSeZLI
GPNr5jd8WP7UoY9lzAZK8t69PXpTIAwhTDQ0lJjr1ZMN2ZyWGvs//+k0jVSyfgHIQj3A3X/xSz38
1OUC/UTg5NvBldmiHjvE597qEA9m+fu4XNVzqGdR4GJSgleEfpWO5kjxILNKivWIqVDo2FAJPAK9
uaqtuPv5YdYfj9AkE45bhhPt/f6n7879cmFJxx7VwWWb50ptXk9spzKJbpm3gSbB0CG0/45yRzgG
3UF6thhUhGebloixcEPXVFcBka21BUtEE3S2i4cDqsjZo3OZWQ9kFGZdXPHnTvDlZbIzzLgNgpOH
8zxRT7m0LRfUaSoD5rCe5zG1kZgoRzH7RsqJmSiPTdT6DCYRVeiZTmQDzxqXsgg5GcQg+9sWxEGW
gD50w3s/m8tuH5iMQGCFm1Mahx7FsnCuCvjz51vPUctcJ7sPljD9N6ke9Pl9UahZCtc2A0LcBeIm
abrBR6jdWpjmh55tlFEW+qqeG/nT3KCLlWL8u+knC+nChnb21rq9cKrEDrGp2cIphfttkIrIkUMS
fJxf7Bq30i5mK2M/F/PyA+VIAomEPE8Tst0r3Lh5Nqhi9tiwJUTA+EdpJWSoX7ZDCt3pr7lKdEVq
h3/uhNU9AL41R9yq/K4Hj9akrnbS+42aiOVIwEsUiskJp0f0xv9xdAdw1u2FXHKvCS0d1O77k/f5
9ZoUJuVmH4+hAgR5ffwGZ/jb6hUQoAq0WkdurMY77v9j8OwcUBpvo/omKj232O3XbcTjLjKG/d94
2hqtvbrou5tEbP2YG3A/5LUFOpfACIb3mpqCv1XrPnoOTKgHUcGMoH5CNVQiWEjNIF00E3MPwwQQ
O/C65URLGPROsV2OMhdQeTx9qT4hce/Y4569jo9ENcq7adIi/5CaddAXJSHyU7anHcw8pinHw98z
O6/86vevBgpkd/GqcIz9Kxb4eF8GVcrcru1FmYi3QBJxlYsaPx3OB4iPTeOf4/xbU5wPYn2ERv1I
UPJWkXo05fRiLp5PAvEB3iM6AWOGU5yyMuNRZcE292JbpcvMCdAyCGX02LMS+vMV5VMJB+Q7kf2j
D6j1iFuyUX7MgdxK3yCOoQo10/zSuSyJGSvhXVnsOwELQpu4yBrJIVKBW7dmwVZzH5fQfgMdyMOO
/+pzPpAAcmoJEwsdrmLT5yl45ERVUFCZjufRJnoczB9lfSjoDHwEM6wWUsL5+VPqGH/LMeQqprSK
9NfZ2Nk5r7kfrN8UNgPav2Mz3Zf90/1gI40LcIbqkWAFYJn2Ax9tkJlPfA0eqgpTQffM+VsZIzZ2
cEljKXerN+sLLZG09yEmyBYF1WFECJnfTuPxqBhBBX/4mXYIItbScbYkz1JTKxUtJdTViQ6DLswO
6zmAV/0iHl6eK5Zf2/9MC9J4ABu51GFFYXysfDgVGvqpsjBJQ07F2QL65t5/MtY3GDMupRthLAaC
/gf2FyxtbtSw9iYSb6mLuxIS8YSg+vkYN7Q4LmAewpokDqfW7xMz1z0acMT817i/sLDrIUkTcpkE
/Z5blSCf9+TEzUniA86yR76Y4zsgReWR2ZCX1A253ayV/FUahX1FaQ34hyq+QR1m2zflvHPJZD+q
UagFHYXklyM8Su/Q9H6G3t08dHmZbDHyyP5ZLN3OgtcsDChW3xEMEq0K3QzjfzheK9Y8Q1BS43dk
z1419G/p2aJ1TsQ/xejZVpOugIAwf0fk3QFnloA8EQpPXrJJtWNkDk40cDOEZlkGHc82wHLB/QC1
7kNuYfRIuulDjNu0d3LyJTamhVyd0bfCUJxH0v+Yahqahv6rREBoEus9dY7SrOHV4AXlXXSu24C8
hsT92oYurjXgZ77D5zXontlmL38M3zy9UUy/B9mxf/7KA5imhWfSlc2wVbjXB05txx8EWHyTsKHI
O5acE6DPyep3Xxb0AYuc4SoUH9bU9Zu4U5T92XARYg0y5Y4vKETs/DH3WuxGg5qnjLXuHmQLUOBU
A+ADXTGd6VVIu0ZIyKtRrSjFY2l33W+woz1rBtc9jNk8BpGO8VY32Crh5u3S3dUOvnPaHR7e2ox8
JihVYhTSu4waSIWgEGY99vB96rBtxZecso0gEEsJhf7F/NlvuTW0dUmaJ+gKy8Z91l8RFwJD4fRV
dTavIsN8H/EvCqSjurG2Oqs2sgt5ZlvFKO1IX2uOnZDArx6GIyF0NM6W2XMzHF5+2VegYJQU/BhE
8jf3eoSSswPu8cNAkOcfTFHixD7JfKcVPG2KV59pUgM9PJqbd9C63GELJjRIfvjGEtmi96me2tU/
mFQc5BIp9kiChRzsRU/g5lHna/iSFmhdM+cz+QTwDagQWURJLRu56cLsUzMesHMm/jy+CZSB8wtN
0PWhtEFYO/3jw8tMK9Noj0HcHLBE7Y5E39h2fyEoTi+JrUP3hpnC7wSpB38feZR7sWpR0yxPZJO0
BaZRbQvBaBwjDTHgpcrJw0NxaOgMjvEMp0N+1OzDvE5eDaRjdZSwCM8BEAvm0KGaDoEhAwJsU9Ox
cHLtSOl+yULbp8P1MkKPM/WWnEiZq3B2QU1Lb9uAALPqe3ht84568QXYFX/pjkfUC+xWOtUSjgxs
PG/uM3yTzwGQF9iOTfLN82nASiUCUrs/Z9xDkpEJWSDycogKuCgqpx3j/qGQpf2fNTrELC8iFzeD
iAeAIeMzclkxFCIspgoqeHjYBL1zTiIRJOe6f7HKiCLO1qaIZDEd8MF4woMTVNSO3K8m/AK9bNT+
NuV2g6kJlk5oV80WwKP4uTip7LFMY3rFlnRsHOAz0PADa1z9EaEw9GZPSg18Anzyr85P2kJrqJVH
ST+N/jRUTS7AsyzQu2iA7TANq5wb7Xibgik12urzBQHQXE+UnuYplWXtpRmxLdQ4a2XlZ8QngPLM
Ik6tHfEAsx0v0i4LHHf2YxP63JSA7tp7Q5K7KT6Yl5XKBK0tK60GYPqYYBmxnIgIwwXIoz3l/D0O
FXydQ2fIQ9LZgZ6WOO2ntWdpdJxJqqK3Q/6KzE50iDnhIpVmmAsI3M/wCpABfLYkd2m72ksfQpLv
/nNUivhZoh0fLEvTQ7TNZHZcNEmedrUvtCUAKeirtAOYlygVp5nMbNe63Q1kpDOC8u8r7yYFjSSG
ePD0Bz0W7uTKJKSRHo5cwKdCnSC66CBIaGas6gAYGX21L4XuFuxqyInuISkJlnTOudpiHRDBYt3+
hPWEbNjPiOB5TPGwwJ9EeS7DS/Eln6c+1jJR7m8R6bJsHd4KS8xKxk352pOrc1jjp9DT/OjmwzEK
brJp9KG19rN6WWZKp2TkxCCq83GfbslzkEWoJK6oKLDjLt13xnAlzNWwOJt1kResq/n91Su9Bez4
Rc+RppZn07tdQhMJ0CxPECPq4FI/0p7wOec83+7d/iLhCss0wip85SbPGSc0yRNyKf858dpy3YUx
6iJX1xcNOwgXmvshOJGUZ/jUA8D5xgpxrwi0QrMTNucCOMf5wO1CKn+xlSPDeby6l+1wMPWXWKUY
KrlBZ+7e8k/nk9ByO//aGexzVnOE6poVYNRYoFV64OEHys+1p8HhYCI0WEGAoY/dSTBcpXppRetU
iKYnEVl0pEslhtCExiyXptHiS9IH4w2QnWJq3kehebtMKFucRLgFsnal3NgGjh6fAGSd/PeszXZu
65gj54OmalGaj3/PtpiCRPxk505OjLZ5AyRPCPYTjrpEgltA9AURsyKFjSix21WnzHoQxG0KkHN8
3IdDqNA4riulWQfB0yYqXkK8o+A2hgoorwFALqlmO2UAs6EZTJcxjmo8DrG6DvbC1yLd4b3PEPKC
pMIx1mFJY2sTIx3PjYL9ufr45xLOPhN50wU5V5ABhF0g1pOMivN5fVK51L4HaEmIfih4ZAVSWePc
Vem4ZF+uMg+MQLT7raQc463xwhZjK7xLfNzrDHeaRJ/NogqtLQRT6y2ogBpKnYOum71ukD6e2ILl
t875EHAH4v+UKO6rAPvNsoSo10eJat6wIfxa1rMPRZhT/Zoxam1GbHsd92azTT2IHdsKMIxx8CKE
CgPLvooxJ0CcgyPdAK0IKRBb/vSS82TinL/TI6w1i9StJdFH17S0oYjlXxT+FV15g8ljiKRK8qPT
8xBFdpTmJOOumDy57IOmASHznOpsOQj51nwed1MDpRzhdfPrvlSrw1NV4VwsHBcVAV1LhN6zQ+Xo
6gv+WJBkTrrauSvhSvjR2NP2ldDiiCrtR6CP8Hf5nSZn83pUkzZrybaoVDAmPgxlJ7skxo5pRA+f
ibC/dnVpfWqSKWB20dEeT1CgGWm7t0pmoy/h3ENWdfootcHFPsQn3jBF7X+2TpmxPxVcj+RYDD3J
wPm+xRMoR4p2c64TR3ZbIFFAAvUoQTNB3BYrDcAwpdEm58ubHrglF9BnolrS6qpIvnlPWLBpblxK
p6uJ3eNgd5LNW9mczOHC6Lo3HZ+iEF3uNBksk99UbEbP6Wj+xEIc6krKu1lbGVeiJ6HPuQJVyCVh
mtKxYbDkcPy8c3JFWilfaLdEKjadVZKFo5aptgMzHEa95RbrT6Dmr6Q7syrjHvDx6qB5447JtdF5
VbFnFBXzrC4PReZzlyUIC0oV4ImerpaSkaQscEUA9BVGg5cqqvvYeuzYHyNiJ791bNZDa27+rZ0Z
w/T1UBCtAyDT0YrSz4EC/OuA7yAbgWOIYQGfvHzpK5yrqi/wQjkB8nzobXrgxa8sNbhgZMSU5/fm
QjOpociaQqyI1GDox4b6B6ydEY4egn9Rus3O83KITUE9hRx7f+5Us3W89PRTFRvHEBmnBbCCLgy2
TCXneQANRZ0CngEto/A9TRLD0KlyNRZngwIr5dcpsyWP+Cb99AKjoOBg1hewq3NI30Aw0j6qGRwQ
qpYIElskTSOUEyqmfpYOH66KFyki3eqfhRMVTxkH1xpG1//fS+gTf/aAejFZplxlc+mvp5NIoG+m
XT0cLliAtHoDuU8gV+x8k29XfhBMA9DMlIBSXFMLJydnqDPtVlUkPtHYfCJtcQXCMgbem3VgRrd/
Hxa0AYFV48iG34ASCvGAGwpGBuYrVa4OMGSmNs4iDBauDnL+qTLmFtcHxir4OumZ2FEZry28szOr
A47MOAGLD7VpYdYfM7tSGV3yQ5Xewi+SEaK+rMLhzbVVdqDl4MpcQDLr+wroYP86eOcxF3hQPfHz
+UEPHetRQ+DSLHWvq/Qog5iCaUUp1c7ydMi5WiYnFgg90iLOth5HqxJ9/TFOtODy1JS5pBaax+nx
YM06CL8YjP4FVOg372qCoVkfs2uxK4TC8jnTwby4d1wVf0x9ts5Wwv4AbY3gwzmwrDJ2X3zzxn1l
DZ06NzcfMA0CpZ44Iq/DrTKZHzPVkNY3/b37pxaZBcFN0KwOwtHAz04MuigPg4r84bsjCdnZmk90
MkaAOrbe5YcH2Uy87iQjX4qWrB6l6JUBop8XhO0oDFGAot9BubrJbFpWrdD/N48DPxz0Sy24hYNm
6mXuXVzZJG0WYItSp9w2avSXAHRnZ5oo5e3XrkBl5+P90PgUwHOvhm05TIYDhhVSBjO6gidmyrlv
M2sDtuS64spubqcuysH/eVYK2n96zcqFvKolNKk/NnHqisQIF47LTI68A2u7hvmR4dUd6lCk8sPY
aqyPinXTPulCWTfK9h47+Gwley7cvEKj3XWDnjANYBUvFFKLYoeVJtOxeg/+W+wOyzaNOxUEv17Y
sWbyiZ3h7EtJHHkY86NP4WLN02UnLrzn99oOF7EODrQI/2foIyD+X8s6PLAz3TWiW+ddDHqtpdqe
EwBKy925nk+dK/kLIYRHpE/bnRct+OadO5mJesp2SbbYqW26Swpmp3lVhNNwaxAzKdIGQse/T6NS
VPT7h51XH/+p1zRpVFB6Heo1NW5+LF0khU95MR8AJjUJoQeZgedDu5jN2DTEDbdXvv5mMjmf2+I+
YvqlvA6ckTlitzxTTFlfsU/CHo99235LeyrKKHQGCoJA3GeON8WktavGbaemZ38VfaMGNQncpJTl
9eVd+pm8RcBJU9s73I4eqzxAlvrwloXc+0il7uRNF3B8xr+lnl6SwbX7klhx/M8soieqdue8D8eR
pfCet89q6dW7t26PkWyjGOE+j4i7mEsbn0v0jIdyjRFAX3V/f9RXEUklkIX19wpdDhtuYxEVB6PQ
8AtmHR90QSv1+l4vgq23U3GZYPVscQW3imYfhFa/BIq2713YSERi3Mk7Erfc/ISuPro4HJo1Gk3V
XEbRN/aN+DbjPOMB2tXy/HHAQ6tL4s97kxbS3lygIkRh4uYX2Gknt+4QQYRynzGvuzOdP9K5+8TH
ERaPFqXl57CcP3xKC1Owdm7CIIkmGYSTMEi76URlAOI0EvpfMTbNYViaKH5M3ENaQ2XuvSk2flon
yWYKRmwLe2PMFeVQs8KRlJdvm1C1rH2NhOZskUeyq0N/ltsvVVRKXl6X0ttG6bj/u3Ch/wQhyzcC
Xv7y/m8lbHeJYfcb5wTiuBnkIzChWCPniqg2cR2dyU7EiOk7ejsi5UwkIfslXwCabYQuvLRfqjUc
dFTWR2xMEprk1nvVRWXhTe0oXh2vvGcgjOasnrU38FRq/vTKIRbEmqv0oADHFCqEeBGTKj76pdfD
HAaIxlCkkx6fKR0S3oFBJoYLKqwthd9FVZbkYdGwLRcFAOYMJqgPo2ck0XXxTqQoYLt9GN0R4ClF
8s6ihAo6p1f80NoNd8w1nIc5Im8PdUHfUD4yE2hbQAd3l6R+z+uANBVzKAw4faQgA86SQG5QJ8Zc
NTQU9/ojce8Q33HDCDm1CF4bXxk6CjU3NQ08E0yxDlL/JXpTqjk+TvCtMVLQT3MFJe3QxIPvFI/T
Ic2nbx5w8W4ikdtam12gLx1qRq4WpNMAK7ws/maK/3J6+93Uwg4asZvDcZlsNGcskm7FfUshX83G
E5sRACQTAEJrpYaeV92R07DdlaBslNhY2tF/XT8Irh6ll8RFZHGKYFgIlECcmYiQyKiS27c740cp
vG6BptusjaFK0bbaHGKlHOWLSgkoQwT5ZU3oyJF74n9cpFGf0PXisH8V2++q2huMdCEDc3Rd2BEw
Q9czYD+y37gU/fsJCoQph6lnaxaZ5BWawwGvnsWqioic5aUBCHWMEXMeUZWQM2Sb6bEzGXPbIG65
Kae4LSBPmxs0AKktSmxJ4aEPs4DvF0YH2d0iOOWdWF5LWdtJzGGO3e+oRPqpzaECrF0mChQ0vIx7
y+AkvxsUXdzJCUju0mi4oOKjD7LDH0zpFGg03piUUuU1qxgldKMhTxT9Lvt8lsEc2u7cTHyc7eza
bA0tTw8VF7f16eFdDd51dV99JA0r66YQcVYPkfGprQTIV9NFlbsqYN+b/fTMDkV0KfKOUOLF+yHh
XvLAS7v5sXoiexbWlNmiQzrlI4J3yUT6AaOqxUezDinP0+e7f2NV9ic77fFM3JEMYp1FooNh+DWD
cS9mLRuCNZ/kpmN9+cU7ENcE7T32Fb3kEWv7KSDIRgRruBTQAkyTobbrFrci3DQskzMSZICyP7nG
4+jklTUZqBKmRfuY0VL3jh7yJUzLV5/wbAJs8dvZ+rIVXG1yGQUOpJ/MRIk2bms+mVghrVPV20gL
tWdXM6BFu4Tn02Hr+NMmqU3oHYPQBtBbdODQf2PodS03Yo0h36y4BtLdlxCLG1L7xl9qem2FTvFu
uzkt3GloQXP7eRjj6OeDDlmR9qF0mSqQ97csiIWoKCePv9i41+R4PLFh7U7bIhCWeFsAy3lc8JMY
6REx50KP+HVLuoKKeN7T4np3ObhwBsZlWyb+TjtdzDM2HYnX9sWhyj6Z12I3fPdiMyii06Cd2jLW
Cb4f+lxeGU4ek1GPipxbVDfqnVhsPrnD1v0ShUjelQ1dqzmbgCoJqNfbcLIXW791YGkbNYmc5BWD
MY4KEDgy4yYcjGfessUrZ+mbkR6mO8JZxdOItpkouf3m2b+qf25AkTIM5G7I9BnZggWsbx90YI2l
mz3e8VbdHcMnTZLlE7rRYR673ZUMx+aYVeOi/H4OgWzitJ+53bLDS6BvYtQLTWdOtMcN7QW0XwpS
IPjYVY1dU/8pob/OhqiIO6E+I2y3Rtus+DcFBF4lYy2rp7lgkn9DxNE5Ydj+lWKBFVCJSFCFFQCG
sfyLnX7CUsDLLfG07wMdftnAuvGq/eWVfoPp8RvTpGEnQzRAggvkTH8Qa7MlNQ0qxeDjFDIiODar
CmwlKv1eHlz40nlA8t5woEkg/+yhDo3SG9pOnLRq4c8XPun7sMeunSdY0jyRxIGWfOpw2U6Lgzs9
tYZ8OV4e7w2QrQIf/iMYZiZqAYkUnEVdeoTlefMZkIN5en4fJzNisQf/HSx4EMnO1fUZeMGHxvdx
rdOGMjVdVeH7Sfbq51MCyHppV7me5kLpXlINJx9CxW/7PMvzOYHpX6eQQOgZCVkVOp5HIL6u0Ut9
EQzs10XlFm0aOFqapTieBGQWEP4F3SW29tvfyf1MgS4eKUR2C4aR5eSzdp9D06UG3FT13ZPWHbzd
XSVQYG4imyi79riphNGRQOZTzcANdzZhzoz+fzIS4nhl/s/qzTPhtm4hpCzSGf236pZk3P8g75f+
QNZnu3I+aQxl6JSjWJJThente6on9x3gFGG+Yw50qwwOmwxgRkDtMtDPrciOAD1iEJIcDOxWjM3A
xUg2+JbzttbDcjt5ALD/jRz0G5MVCqAYf/Sj9vdxr8+/8OMkqtMAQMLa9wQ7Pxn4jDaylTMdytpt
UlAfdPyeFysh3UpX85sETXnLAdmFIa1uGSQxnCf2+21RJUGU43U+XBCoXMd1FHTE7+EOx0dStZ2u
RzbNyV6POpNCr8Xwhtt0uWMUK8159qORgcK454fjOPu15YPT8JGcOktZPlLJoAdkQq5tZHoUEATJ
39HgYzbLRs3DRx8w0GeUkyLTlxr1kzbUD0vbMl4wghwb8KFIQ+TkfWa6Hz6blJ57uPIIHx9wOLkE
vZS2TjvbugU368hPdH3N3576UuVpC9S1bVkWOGaWzB7+OvWDNtFkpdlF+OddRpsLV5Y4uvnaTd4F
9fHltsVB7Og9nMWEU0b7XAHTJeUOarG5y58ZCoVa2rPNYLi2ieaaU2aiYJen6SolnpsLRQdU6ETt
8iJh/qGnsYihk2BU2+KML1hpmFYlbZvKyvgC4MkPweqRTvu1DNwOzy9P/zv7YGPDYvZY9sL4fffK
L5FuqHIcuSXuMK7oaRK/t3Qf9QrlMWob1ubnVsQzv9jWTQ+tZLgNW0SaFT7++KH9nM/NxKzPUN7t
G3PbBYWboW/4+NfHfpus9x36ce3z1FxL0oY/i9th3U7/8lgl4VKwSX8cvwGJCpUjHqkJyZYkmE7Z
gU6fXrQy7PZdykQ0l4BdJq9/FaZzD4LHpUdm574XpThWsrAHno3MOYi4+CY0P6+Cml/FvdyVwfUK
YPf6eunJWXp2B7YSSmq6N7/jVDfpCt8imaNyYIAORD1nL1MD3VzVaaKxYP7OcubofTC7++KYyWFP
S8WI4/daGyMxKfxaOeuYN/WIFAN4HpttEJVRs0kIhin+oOGzMCUyR2n1ywcSO7+B4I5wYMwwzhPK
kvuWSZH79GWHMRKY5POVMleCWg+BSz4hWPzJwtWRNEx/NR+vft3LDMKQbbzqhxR5NR+dQ3q8QUhU
Iz3JKlABSLnT/3wDcsBp7ZCpKcAuD/9W6zUr47EZwqaueC3q4nsa22TnJVRue6O2tL9T6vUt1cc9
uM2aVCS6YGU8maaxHjqsNJYTVElwQU2SsjMVXl3J9/SdsYHcuTW+faPi9zCC24SfnGyQCUpERZol
1TdulieuplID6EiF2Fh1W4ldBG2mRrsQPNIkYWKL5r/lvut8K0/KAq8u1Hr7wF5SYVW6ffF32NjX
eXCjtqpxl1MtslT/nvp6BUvujC2u1GcsZLqLa6+94TxbpUhiU8caG7y/6eag4x7fMCYCofubJKMM
2GlRUP885+vM4wzkKL2m4lLhCf7y9Z12LIZAvcjGn6o6Y6YEh7Pxdds89mygtG0qy6YYHIARVdL4
Gpg5M3R1m4MvF23ZtyGxWaXhfma4jbyVJKD6BcuSBZ1TGc12Wf8JztdE/ihsNKb3o0fCQXt2ynk4
KVkhsvG+ROGDIC7eEn/tRS1I3pQrzsbGMwHIAPDR22cO/ryptcRdsfQvC8c2YrqO9SaXiNil91fF
Ojl0/RHE0BAKxXOjsbBcoqmKELm9f+HMerc2t9u9h11g/Z0Ifgnav2Ov8rwS5Eg2tTF7QugoSVGq
erYQFTz/E7+zdCPwU8GoYDQe8/mXayYZJTZnwT+Sd7YS7HKq1cjBwXRMv+PZHweEJ6KClokJXUbW
iHx6a8eawQfVSq3lNHObbC8z3a/RKdSFy+qEebZK0BQ8uI6gpS+4fAZF8h4Zep9FvwvngFzja9oG
2klSdUuGC6wCre5cu2rc5VI5MxsMWnSWX48f8dJpvZTSLcrTm00AiWIpEg/NGIPufql0P1eCP4B1
aVjgwxpUbJc3uD0PxDhJwJ6yqDUPdJqrwBCt5Q1fLy07psYod5NO1qXs0jm4MebE63vrL5Ig8sRc
busw15UvOMsZRh47fyFr1Xk4FN04PtvoyVV0ofCnq1Yt7sKfCfu/zF02htIat3JTLqyhc+YQBPRq
smfpi8rs9tb92n3CtDwQfHPUGNh1dghVL3UhfGlbpACW3FJQtat+EwS8380+KSO65UsSB6Gv2te/
fi2eQZZPTYL3GDD6KRznJDZjleRvHcsfD/tyhZKZ1gGe12qqvPjCwqlhEAuZbNkktjxloGPBrPSL
qtdhqqv4Hx+Fga+2WFO32eG+9YuvSleNZh/mUVh3U7OCvDPRhoPS3AFPB720KyMNBQuTnCqBZItF
LdPmDKTHPlv/nkdzKKswvgzx6OW/84n8djiScTVu+VSgwMgOuzdscPN6XDKr7E0pUkuzid+fdKZa
dJRF/kaADrtLa4YNavcLI8NVXuwvq+3ucRXoHjjmeE+zdttxghf+DBvX99yNk3xTWCVeqhK+kKIu
12ka2FAbkZ8DgmX2UiV7HeXMKTxvZ/Acq+swASqvyTf61qFm703WurGKiouPxnmsC4L1fLE4lZgK
BCTRMHG5NaKzKjWT7QG+I4Wkrjg0/nDUgokzLPYt23y7wfHRUMGKk2scT5fIADZMUqQNppzaaCsp
nDCvAJcL1l3GjT2zXF1mHvVr26BGILXQ/ex/Hfov40tWe2ymGGPf1mPCxJ6khtn95FgR0PQLzu5+
XpVApL9tyvZzY41rHQKZ01QoL8pAlARzqs8LV91TjVKRxTSk+laEtCc3Xw4Y8hodQSxXqbo4nhG6
0UhCITrPRCwpIETPpCXvLS4emqpwWMiKKUsTPrerre44FLonsIoHZAaCrAZni7ui/Z3eXfKUdslw
y6RGulcXq6IETYEAmbcn4FL6X5BkM51e+TDZNo63jYYGLPDOr/6G8Iqt6ksVETFhZEmDsigqBigO
Ixk00EfTqgz9FHWFI9K7tddukoZoqBeyPzlllJwGXDjf/XlK+K4tMPFo3/qT5WRET5XywvELbp8d
fgdNQuJjTe11C3aX0C9Aog3jKjQFwOOVVTlZFirjJykq0VxhqW0S81s84T92BHtIXvPNRFm4CS8D
5NyzvNgPayDDVLTDeuwz0GSZxuVQ/+oANIlyg2NcX5xPkLwO/AbdyqFGsVijhx5rJ1pFJN2s1+VM
0izKBO6qvGjalYfAyWRRWGDGK9s2G0d5xC3lcUrgGaAKX9iOpFzdgfWTF0Lt/flmPZMleTc+wHlg
LFw71zKh7ALvCL39PxzvAgn3TaAs6Kz9fUH/I1x0G4bfZlY5d0ZdSFwYo6lmw0k2QXjUm4g8YXM+
5ny6LtMlYSfdP/0/TIHycWSzpkLL0NPTihcNiauVP87o718PxJVc4eRyNQegMNJNAjVi2Qwch/9M
f0DaLxuBCeZ1zLqjWloGNeuQrHqS82Qio/hyaA3idsAs6sup3PMzKjxRaj4R/O52X2+m54KqfDgU
qMalJ5h46U9wYE8ob8TWjGF+wOecjufUPIM9eld0Q6x0FtvxPgN5Ltl5pxOYL3py2ffyZxFg05h8
xs7yUKTiVL1BJ3szLoJoCg5GuWXHupRTQlcvLt/w9OioyrlMua2G9ojRINTT1smGHwfBqZ8lcAtY
CApE6RTlJhvSoNwjvtRUBbxTrD7E9dqX1z2v1dYj7dLkRNJFxUl/hC0x5WjkUdYYOQ6hVx19nm7i
+cM+ZIoznW09QMLLBwVkiOiew4TLZulkfdyyzSakjBJCso8a3i8pSjtuwn+fUEfS10CrrOtyByZK
6WSsS+IgZw+/tfoczTjPvZAxcGr7n6RDktskvfg7fAqcLIYz1jWPEDuuMJk6T6xBXz5G6AIVA27G
baFoRyrbMGZlgwCvsaqNDb8uNnPVMnbbjrQGud0TOF+vyxs8s4RHU3pyKlDjhc1b4WYh/EVJGgV9
hsBf30H7ofJvSRkZLYebeXQzRRDnlqKZzCM7zMg7ZD1X4/PtwJYLdiZiz/NCU11dlvYUlInP5i8p
cj2TSkZ6gkDVIA/KDjbCVmd1PVxLCF8Y0wUsHKXE8HaxkTwoPN/Y2azahW2quacNbVkmPS5NDc7k
Z5gCkE9J3s41cagRT0xMa78Zjn/Tj0U8yhh/jHZbkuYBmzu/7UOVjiLpyNj4gnBRHIYu00biqU6g
URmgbPphma+ilVIY77RTqRWytO5AXL2PkHXTC81aGLgWjXsHL4kslvNgMqm27qPras4muX4AjDGt
0kmL2yLYQSDXCOToDfDQ3YJ06uC9BJv0CzoT5eTB1T0prg+MOit8N5l+VHQrMHeEn/xTjVLEmjER
zqrWOhdxPGmAiQERtHBkIjHLpCM1jJUOvD4LcmVenjqbwaMIYXq0vpu6HbZzv4NCEItiYbUHKNAV
OTvKHmaRHEeFJX0qywdigh5TaQF7rSFyxUXj17H9gFQSNKG0QjJdgfwslQ608iSCxglEe3UFmxzT
Rp//vH7BN9pLo1wJAwaXq7lw8oL9n96NKZ+lf2uiSwAl4Q8p1LoFpGsB3G0m3t4WczJdpcK8Ff6w
9ziOzSGXqHH4MSu9kADRhhC0TUiPY9jA8CZ6kS9HMURwKLwoIxZfqu2slQUllC9DxNDNePnDgl/k
EarjDQMbR88KN3o27Dv/PKCZWQNi5+wU3xLQMCcSRzJJpn5YyxXeDULeYB6hqXM/vuVRH+J4nfBT
YMc4KLNEX+k/jDM23m3VZCY8jSc2AYQDnaYt5bJ0QzhP1GgeaMpiB4K+yUEhvHhggrR/1kdxAqAU
VNmM00OfPMlian8TVdtWQQthOxzQukKQ77X58LHOxDng7ZCRhDnACNoynry/Q2S8Wg205bTNOJkG
pY7dpcoOW85qOfcD8sXqvOxqABU4iGleVfSATHM+yTqmoSsOoI3q9oAAX1QgXh6e0FetBlZto1t/
dXZ5cIkHDW3+EWewQRVp8vZHqvU9s5+U1sUDhbnQbdMfLwSVBNsjJUQVZH4WxliFnlGG4cfhvqvW
QiVJ9Ijf+/pssdmHLnG4vjjcK7E4orMHa6c3kYKGjbAwkrGAxBznWxV+nUi5gUhQWzmo939AY35D
qPf8qmRQAgrWVBAUcqnTG9QgRXcs/TscbkdJBS6Izh+GNWibI9Y0uV7kmNvK6eXiog1pQ/NXR4yD
g4E1x8hX394UNJB6HFt/GebOlc8UUmbS1Om/K5lPMOafDXm0jSJqiyx9mVywQy4kEhZEFx4Qw9sk
sT1OWUi0hZuA54p6vvTbmuQ2LdNvSOQQwJGnp7Q1ILiEdouPtie/0JmYcD5rDtdvGqi+Gw2qnzCF
FPONnmRKYpIbCsu516bIektU/nQRDPEspi5rI1PTLMmPIcDbw27OBaLD+2LzdRyKm7nRFbsacJL4
Gkn3xauSnUNg7LKBWQBN+bwxpjqeV4Rn3wYFgNsXZSoSBGuOCkID43N7OW+rEA932w2OBrvnMQwr
TO8Jxu87+hEOU+thPnqVziAAYdfnRtK04gEv1mofbPa2y4Vq+9PsYRkEZ1nd8ulRx1mLBhiWyBiL
xqesThULZt79XF0FuCK6BSa1ZOD9s+I7quQTtnhLFkLm4ZX0vmm2gWecNo064sdWF8Uix4qCp0nx
eQo0mBsH1hRJ5v0GZaIvnhTjLWKJq21tC9etosnMyVA1KAQrfAqeYWQvUor6uMOFjz5IwTjM+4w6
ftvBGBdzfQgWeUUwzLaaSC5yLBWenWtwrbqhREJpn3Y7kPHRIL5pplQqXx5Gl03k0usrsTdZVFaV
DJ6eikyb2Bmtj4RPtlV4nX4Ph21MPWrNAPPB1OEkMfvwuhMU4bZYaGBmeYk+1IAE3PUi4TqBcyaV
+3C+DRL4upKM5gZOXTjRZ5ZWzvWCPIxd2AH5izye023M/6dSk2H+ds14fWwEk08If/BYzmrALfH8
u6PnDBA98Uu1GaUtVCLulNjmp5NTBsKOJhx90+qdhHduQ7eBT6DPSBpSdBQmobFv592bB9F6XYHs
kSrHHVYMlbur8AI7igkFb3gpdiUm/DBPDr4q79BxR6Yt0L9sad9aIwqO2dTjUiy0RzLMS51zzcXu
CbBeFcXXaPxES/Qa5mdkzdoUvfFQdNPolTwTr2KWcBg08/iEHCu3zznS0F4i8fASIER6L0pYCc1j
/oUfvs0JPTiRbm3VKogkfgqG2ZIlK4XDhz1dUvIMf6NwnMFF+lfyZGZtVM/+vjBsJplEhmwvXnjd
EVz+wDfvx83MW5VidJcNDw+ufjxoB1vqvsz51CbK1sPdvlKvxDbfXpvZj8i2WtdhroQknaN/3XqF
KQkcdzd26TZ9LFev/1cGIkmuxETGTAt7E8VisBZz9GHR6rCGNrQIwGy3u64Igr/6z4h2xBYW2omt
lEjiEvZBlNrmy9GruRJM731Bht9vU2L9lUo84MUeRLKiyBflnDiFGb1s+mOkiSxa+Pwbqq1wuHaN
vw7TxZwzt+E6TwiaktiZHRyxxlmj4najplmwLyDxxeJRd7Z3EnsEbWMV4meSwqyP0N3Z77LEis0q
+iToMTm4VB8iOBtEUnUU4FsBN+TkycN/9HwDp/62l7ysrTGM2/XlVMKfkPYVk45+y1ffzOkDv9PH
JW+0OEfPH0ATlWHtuYkDx6C+aEknWkRMJR6niuzsWxncJFoEhAjIbJIPLzLQiekMN1MbcmrxQpoa
kPPqYJ95ZZ3fIdm6Trdfhd1VsSpHOR8yyBTim5tNrxKDv2ZCOIhDdvWPPH55cOjZGoW6+vAyBll0
4vbAGCW5pXnuFd8bkoIQUgAledLT15j7wlTTZc+QKuWtmO4PyBmqQPSqXshma5ZtMV8mMULp03UP
jkVAxsYbdN8ijluWchGKFSNJ52OOvQrZQxElGbjJPB1IoAoLLWt6LPK8rKOdo4f2WXGl9zw9NOCt
90RjwioeuJ57wDr/qU+pzlLsIweNCsFNXaCBMjsxp0rtbQeMsQTrEItd+DIBHWLxrE6iLwLjfiUa
U8IJEfB2rEBFIv+D20NaViqO5CK/kBOYgxnxXOWGk3NEH3boR8nCJUcFQNqWJYOeSmXDCxuhh0xo
F2g+EibbfWv7y6SQE5Tm7d1QWwQv9Kfgrm+NJ32C5apd6wGBjKLmp75VZPTivRXTzeIxWul4pWx+
tZA/izE0GUbeYommfweLwJJAxx/npfftFZPHo3HndLYahUsP5VhA4Sif4YRStZLsxkPk8GhR0ZR8
Aq30E4Jx1xm5gLye7s19fQWBdyfGHtHRAdhInQL1CcCu8SXrwoV33ojTc1XykQ9mQhFsq911eXpZ
jW+NcWmdbxqCMFQOJEIQ8N1Y5vcH01vyBMnqnLi27prD++oeq2hNrMd+qbZUi8rFcMpvCLb2m55S
LQQGDXPgUESCMDTLwbS3RUmtzLYUr049XjvgfpfChRhZFB2D3CLwpbMFNy1QMfCYl9Y/gEnZXDYD
WQuLqkpJpg8VbyFEyD8htkgdBe/4VVgS+ccQ+mrpRPN2J2Odjukmy5Fv/l1AbDkaDzB/I7BAPYF1
t3R7QfPJlDtqSFQ4phmtptfFX6nkqsC7+KYNkZRjtJh0QT3rN6YU7k36kmYWAF4qLuUcFMUBjG8D
hVXBc88ArP5VdMvCE3/pvVq8l2tihctq9OJmx4zbaBBlFw8U1S02MPwzmAwGZ+NhiyfB5jzLJiY5
6N7qgxMhwFiHZnV2/0SDr8na9xoOLYxy+yMixzyuNzt8ZANrDUdcqMHTDqb2NmpygWIrli/xaPd7
OKD6KQp/75l3mUPQAj+U9vadKzOgz9jBY3ko2QyWzyB39Z1O+QpjZJW86KPcnz/FHf/dA3PMDjao
7HV0s4TFpP+jHc7y4+Y0A4zGJDdTdrP6sssCBxxUDmJxU14rHVZfCjDk0XyiUPyKt1UPpeC0e/bK
zUrmEm8+1A4yIMEh/9vjtw6Gxekb8fsIZqtNwgVWZRG2biKLSNT+c4AoNkWDB0d1Deh4qJWysU4Z
SqxlJi49cYs4j7gZQCBYo8cUeovhmnKFLXxmbmreYQ4GIPJVgm5Qa6E8sh221a3fihwLyxJnPZB9
liJezru453ybXKt18aHLq117eQ832y4UPG0QMuvsvIkLZKmKHET6f/d0COxGck+cSRkA8zFNmjtL
obh/r3tZDkU6JjgkHGAqdTOEvXKfQrvZx6RYZbH0GUo5BgLnIiWXGGgTLFIIiKFBmV7zdRQsOaHA
oKDGfzB2leuOUuy/LDC7xYCF42+6FlsK68H9SrLG7iU8hCakPcb7BAj29m4F5LE95Jk8XxCI1i1U
nEmq0i1KxgMkjI7eVlXXiqWoD43CIIH+NNRHvdoa/vGjIi7nyYgm1XkIFU0eFi/eGU3+btvJYLN8
RkpaXSFBtAXGpkBfJivMJsfHGqNt8kfp5CY/S4EntI/eXx5nrAzeD0wkg8gktfLi6R8HIkxf8Yyf
yaupLHVUmYx4MMOODmqDzxM1gGEKz0nfCk7NhUMcM0MpM3xBX7N6QhN2dFgTPZBPOU0XQ7BprxZH
H7PCUsSbxWPoq//5sjrldxFtOFy7EPictPBlvkAQJsSCBuaELTllvsXMcGzUiOvJtvt7mST69MLo
jVXbGOw4iT87XXWs12aLv9Osie2HcuJ50lStf5SzhR6levgee+mL4j/K1YN1PBU2tD791nPv0iWr
2XErP2Y64VyNjVVrPMJYIYoHkztOAUo17ukFbmCVVKl40MDQSw4bJSnuvxitz4bo8UxwVKGzp9Q3
ARxVjADZYtCO/Al7Bza7962OywY05UW6lwatLd0LPwMKrJJ9WbC59pgoeh+rIqwvpn74RyrhN/nY
4IAIBidI5vGfJyCzXOEG5V4l4hWrpxuyWTWu98pHtYTNyAJRmFGYjrtVFOcIdFkB4BDvKj8rQqpv
swys+50AnZiNaGALGDzK3xFOvB0sDMDR4X5mbcM+GgY3je4vJkpiaHNHcbZMLgh94Qhoye84u4/3
BSOjZx5EqFx+APEeGvcUYRWuI7/C+j+tSpWZfkNgx3zTk4oK6SAwN5QfQxcm1U+mi2TqTi2nf5c3
OxVducpbMQvi3MeMCnpJq0SY6IR1ngqZjrvtV3qj6V9+Yw1ehVa9+2hLEyCMOh1EKKCrC/kQkB3Z
I/Kqt+Yjw0lKMVBPK/fVR6SKDSppyGIT4lu9dfyCdOEUB1s95KmrvMFuRQfXEWmPaBPYCuuXtkC9
pUDbmLlq4hM24CRU4AXMRsTDln7j1C3kL4LQlhl5bZ3kjRHIK5fS7qnMSKSiiRBoMrMhP3/1ocfy
vSdXzbVyFSi2nPZlXA0ay7aZnV+8LCu/MjCcxR5w2bGekf5JiEnS77YuXilekodjOq3FYMGnmkok
RpuEFoI85KXXGuDWMymQbh60saSS4FX6mEtpZso9Fn14qfSD9KEj7IpQcItRnTTIkF+gwEDIU9WZ
IxVOadzFuzAukG1Rn1e2pzL3t/+4zXxqmQbpyHP3km+WARqFt3CS82BQUNthaW1P0ZlDL2Ez6AhV
QBAFkWUrLGk/F5QTDH3ysNZ58A7ZXP3RKYd67IZsuH0n0SihWTihHOf+tqUpjJQ6th6nzd0CWGkF
SL9SqAU5YGeYM0pE56ZwAGCMff8o6UNdAcmApRY6IQd3B2I9XrtvVf7NF9oXPeX5OUgktEc8zCV/
NR84yp6B+XSPwMo5RO03c6zmjZIc2kti2xkvTGvr4gJq9c19QDM2gMX++LQjRCtWxYUIWnGnyo+F
7CL+wygVPxH2QI6KLtGrJkIooZjqjDjo+k7laU4VIjqnaT83d2B7B+cirE6fJNaIumllH/gy9QSj
vdh1qS1gap6euM8Z+VOrQMK0boeyGtQSI10S8ekPZ75LsOZEwHE3EY+wp0eKDdYQP0E98hFerh6E
swTqjhCUy467pw6S/r4HiKRIeV+3smC/MeiPb3TNnni8Mhg3tdRyB3Assx3HnHK039PYSNHavuS9
BQefH+a9IhER/2PgoNkHMFj0xGLTWxmAUHuqly+lrDl7LrGeYNe2RIZaDbqAlWnLcIrPeZPqS9mJ
xwrtI+tLsvJdRGADKhcuVkcpKsSNy3XTZg2mTLeXjy1kSf8sC6Ozfp9h4I+v1gOwWcJ1xnzfCMbK
SNEaDoR0jSvRu2yhGzkZFkm5qM0V3JKaT4tS5suCbdUk/9fMr34Jcus4B1c22j2JTVKejZauFRyk
0zGvnXfmizufC9WaDY9Ch/G/Yb3opSBM1lxhPqiLRNVrY6ZPNPaIzaMR5Oll/CK6Zij1lTJkmJR6
hzvCWjV/y8JUMMFyVCShqpa7/68lSN/ZW+VfM3VF7E8/6RiGTY9r6dpn5dDr50SxzsCOobj9oENr
e1Cp34BFyfE/kID/cWl/QsfPQBcj2K+LO6UFIHke5QWkkiz48SJY3+C00HVrUx+qVQ2GyH8NCZ5w
QUdBPSzGvlx8yhfos0zUOzglpzQhJWr4QpEzE9T/i1mtU2X/cAZCyKTd8FcKlZNSTd8B14D1e4A9
AePylCq/RcSkHUxGx7x+v/5QYFDllDRSonoFU7iizXFjHJe/KDFFPi4dAPXYkCe4f7daMEH2JwXD
bf3S7qR9wK+uSLAOExGWFxxG7yVgc08CFzTcgCmZaV4Uk8GhfYMmU+fVMrNaO18CIoSgM2DbX2Jh
3zC5bX+9a4+CHhrqw2HW0u03geZXuy8SSnNKePt2vWRrq8XimOy/NpnwCEOegZRRu3PxIl1Bbd5y
A2cq2naAqekhNHfAHywFh+XqZsw3kVftfN4q+9VF8BDFDaS1UPWll/UzoINaq/4hrqy1w8Q5O8KV
kKTpVYlAhAtFs2Oel37KxWGeCEVpncEuO3tavuO71s8+GuHZ+DZswHa8hX2Vk3KHs1amPTOS1TdG
2PtGfcvPVbsAYl4hgYB+Hm3kM0txNvrqjhmghwu+dlgklIU29ty1AGfz3A/wWAWy1s3I+82MSE0z
LuPBvKPzJnJ/wkxQVfsNEAJwTjnmncHVT1RVB2Hzl2FnW/oUtKzVX7boFuNg1d5V+bBOppUQn25z
Rg7Hqn30C1f4c9sbS1kzlRO005jMmzPqtHv4N7RoL1sdl6/U1L0BAGfYGRcaLW40jmq/wo0TrmZk
d6Xm5el7hoQcsGhVus8MD6dXfYFGBrGrRS0+2H4JyjQqmHgFEk6MgI79vSpCsEpRiaaI4DMbi4Nh
aERup8ccp3S122/jp2RyyenCoo+tam2//SUJzYM83MWP7p/h647GOCBkCfVuXsO8Yj091dI3gxvt
/3sis6eo543k2d2GfFbE/dDK8GlCfiIWzfd0ZuXyUj6ekVzAXY/YajA33MWSvNISVrCba4P8nHXw
SgbtS2pEyoACqiY+sk940pWT4SPGhAB4r/scQbowLZtoYLDLrqB5reYk1Gn8zo41a5L49AY6T1H6
tvezHkimKZwVnOaE0PbFRXMbT8UtHqCkV40QkSWe8zYPbskXO8IDmIJ8kWweqVxJcwYfbjsTV+t6
k9FzcqbNVFv9zp1zwh8e4lOLktLov+htZAVdk94WvJArUSHgfsBviOUngsjnT51FSKfCAhH5vXXi
bxqbol7SpW05cTcLiG68GshkrmmZtF+zSdGuLE6Rf5hFAUeeXAEh9Ez2LnnXuEoBM5cCyt/cyU3y
Gs0PoNSwsZEKcEvTXKkCD+j+oiklfUC+nri6Zj/iTseM1JDSFPqFklslpWRQH7gSIdR9Y2qXGcPE
sMG60c51VFPEM41xxokkgY6wrDUv4AikbLJMfpzuBu1A250xB765g3phmtBwBFa4aYE+sU4m0GLG
Irh3G74JVZ43GvVfMBuBLFvvp7jkSPNl9wwrs0QTVnNxtwDKM4IpCGuEMH+JYBvmqXCVxgFs34+j
/ghy6ELBDjVxlPHBfSeot5kwuiFnkoTW6gYWaDt+d3AtNf7m8sSp1Br/JR0bAkGJg6R639fkVgKZ
DKzA1GfeZCdpM7XEZhf+HYF2j8i7Ypc5YWPAOWQD1dhZiQCNZ3PbjUDXfwD6OSNXPjoGKH41bXfR
MclsTc8uP5mBwoyFwg9n0hZnttsH7KGN1R8KG81jEK2sFi7frDmigeocG7YBSTvUhfL/lLW7mFZ+
A0CztcNnOJvnwii7A8+FFf/jxH8SRAB4tIfIb2oAVCNdmV08wqoiqw/12eaJNAxCVkwyZgXl6vZi
bQBnq5efubbNm7BAXQnAbIft/24tKsO2QZHOxBohFE6pwfkqgNCSndr3CL/Etespu7txyw0yKqNc
sgpuSNj/FShhXalcuesEzac+cfgSPl2Bgl/igmaLJS/RzpRlw9SQ4k1kD8kS8W7+SacBqXJZYNTn
MpAJaRYDnlO+MUi/3Y2/8SN4Z2mAxZureOwKmQxPdG/qu3NpzbNkOxddJPYfehY84C2drq6/MAvR
PH1jVWd84lbYlvhR8QbKA7SgXh/i0xT0TzMwjaLSrCcAmBSyrcUxP/sKTWe3Rjs87joR9qZ7v7de
Ybgck3qeaXsMh3lX9idZqFLZrz9b8Cymxi3xO07BgVYOLi27gG1X367O1TAvFLZbYZtLwTzU4Cyi
UKxCxYxvA8zr0kHDHIxXVxJ6w/eoA9k8bTCJGDeRwjpsqsWhWt1xk7RFTArX4Rg3ivk/OevjIpif
it+nzq2oKjITdC+hLW3QDsTiepWDrsBtYeA7lTBo0TD6Xty17bmlbHkDTc9RdTstMrjsWaRXO8Eq
zNFWSLOAKqYl6oMQ8OG7vo0if39F/clRPF8er+7xZkyCZLJR68BbK3UKTeTpa9lhhu3y19SRa5U4
439sV5yB1cZbq5RH9emWWnNVDNSJ7LLEjsXTrQ3BEy2I4nhdH66U/ij0Eif4VtzJOzzJZbFXUduC
al52PEU6x4ELR+FC4gLbhuD//exnv2Uu79lfnTL8c7T0ZH6e8VvgP2uEPNBo1FZkcbQycPPnmL+W
qLrEoFvL8ULNDo4sTchEqVw5ytczmNRFuRbyIYME2EbcVQOHfD7FtLla7elDFo8tMOBBgp7Bt603
TdFnKBXDI7ROzlWhYRJVw66dL+bKhrhLHaj6835EVYbFodNWChfbIe6RoC4gJ9D+/eZoSyIF/eio
cmyQ7K5MlKIkyX+fDvjSicO52ckaD94mfDF4o1lUIRNBkI/ow1ltFJ4jHd/K5YYgsi1hUtLkq7An
GBCrifJDX6A1tPHkjkW+dPkfZ9uUo1TuaEueFwndqrnMlWwVdoHYEKjXbl6basaGor3ShWZllz6V
UWxRKzO4MUAX4nkx6eravtsZg9MZeQNgt8eaM7QfRXzK1HP93HQFFPOKYGN2n+LzNRDCdrISDuJh
pYFozlNqoY6aIG64xU+Osf94pKsLUMbvgM1VlBZhssTabB/3+K2deKd/ssRTHw2a4eaYtE11OYgo
ANdLAMeW4IwfuS3hY4h4yteNIRCbo7nHc5EmrFms0EfnUClLk2+uBsCnkjpN4hEF1nTwWjWOMMD7
8lm98rV2wDw+n6dPeVo/h5QPHdML1PULoPKZFNeFeHixkpfOOuK4KQyhoeDGOTok+58HN7dbSrNQ
hzt/nsGEJiqN1rsGWU/zbMxL+xwIEIYK0sTHXCJRI7vRTr78eZPNYxsb0NmlsA670yf0JdBwjCCQ
1Cpvtp5PethrSX0ByjmnjnmIaZNeqcxAp9YdZqrJiS9G1aaay+oS/16QNzIR2LrIFSBGmZop2kCi
OS27xdWRMJJeRkcM6nhxO2oQW5JJaWEtnuXWX9oVyTDotKlI/0q+4MHtnycSHIbXYlRCr3IEoegd
Q5lDheNF3zykBf6sQU3RmbtDlGdYUKODb+9a1cS849OLd0Hd5e6P/y587OVppNHif2Bx7wZO8Ov9
q6jKT6n6HQfqqvXxb4syUaAIVSOWsBdmF4Q3uzlZ6F9stOkdh+8YEkwMmY7Zaw2tQvb+gWYv39Ch
2mD6DGnyfOdufFVRJUXkybibtCMi8dWNpg8y3UZJI1a0wzvf0AkHbyqUbLNrkf4nE1o0EHKyeKb7
p3XJIA0MHTSkerX1veCF3PjPeOlkKouD2cdIH6IxVLf7M0pD55WdIpl4TFSEpTHiQk6Q3ZlSssRP
MLXu5t48VO88rs7f0X+wwJqnnpB7s/q6/rBTKOgl0xHli9vclYDt5AvRcUzTA06w8rCTLUKh8NNJ
7jQuQd/g5ytdzfrZ+mfDK5ja6QOImPxHxRjEt9DvrgC5miWEN4TmYDHWkr2p6dwJuLclYNOsgw7P
NcT2du7L3r4eTVLfI3vrDfQYvDegwpIx9cTx3g0kCvZMQeswZv27bilEVLrTVK1EqWLSnX+XZVIZ
8XGoOZqhCKqXvkhkODRxZJyrQN87jMjqdcj3g6vDWV0FslC0GAAYBZ4sNWbaZJepRCqYkSMZ6tA5
P22VPhcc2RUow3zIrxHKMLSN77DVz7OjbB3JPXauEGHtuI3cwuQ52rOK34EQCpV3XxlU7yqEQvHR
8Qw0vyuJDziKeEx2gadJ+dZ/jzVcs+smOqYFZrB+mjrBgY5BEb09ZvOrVhx8fVKKN3m0oKZQ+XXf
Drp5bFy0cROabnE2ErQ40QlSm9AI9paqv6G522AhQ8aSWpG3gAV55OymMYe3XloPwV2rtGm2/lr9
TKEbD+FivF/SIbsWiS+VUAaXVSQIk7gRcQd9X2rNXjMdWzy1mFVQpT1roAQQ1dSRnCeIdCWLbXmg
yHSI++ZkTmLBEfz70OOYRYcNB27Q3f1BkR2xpLEYP8S9467tigYNcgymS7mq5j2i7OIijto7wbdr
fpJys+4gT6GPr4pvDsYldUUq6Q86c97JU6VZve4JDfk/9e8d02KoHoWrjxEoelIKv32FxBeMhbUo
8QxPrH2hF2EEd/3+99iQj2pJkdr67MCv5FF6FQm7exLBRShAZxNGYH7KWQRIG7aGzYq7z3xFfTk6
24aaXssOfo6FoOrW8L6GFZCfVo1U76bSWaMKIss5xJ2LrnTFbHbXQOX/N0KPkG/ri6lUr7EZ7UFq
OAozjTVD7shrdYyOP2x2obtiMKMgUtwMx/XdbNFr83ZaLonH3mdcysELeghJgD2HNIGMF9bVxBbc
xzyPJStt4r7sfWVby1obJ/g1DMxNJtsJI/OhJ+dWfaPlBh57Tad083x2wnv25dxz2s7zqWFAamYV
q69paHqwyTYOwPAycJ54zb9d06X6DyiRUlleKL6BtJ83QPHY+KmdbPFCk6L5DPuxvxwvCeLjVnUI
bgUWUpHQoP09QSzWZz7R85gxtSSebHa1E24AU/GynaJU41hzQP74cTSWSE0noApEo8xyJhGlaDX+
BKkjPMZQ3GSFt+E4hnNxxF2JS3EF44GomYTNRqzTALtm6n6sHaA1p6zEmgM+liaVysLvq1Zyio3M
qqAmAcW3C8tTnO8toCWAm2H1aAYhKyi2u4PxLgUpZm122EFxyYPyYC3Bv/ZYCovekIdKw9/LGuOr
DopTtE3d6iweCfziqmMr7gy5eyTdKZg+ThHP1eO01mZ0s2MeBXNXTqXpOWfewPXHJAiTf0f+S6va
dc7OgzMD180U/yj5jrws2ym249FYD1l0T8KVDOCJDz43UjQkI/3K4usQCsv7PxvmitvDOqLwDLUw
PZW9P4jVy23OeZJtKt3mndEOrvwOPHtuzr1gwmiQB10BI3fAAf/U1NrQpRdUhIxZRZ4v4efe2s80
BPyC7no1VkG/SPucKytXOj2hrkbt2hHMSCUYdh4kScNRH7Qdu4CMZ6IsmZYLgGtZfBmugdXztFTE
CYMCSoaJDZkeDmYX4LKS5dzIzPcqP12Xd2ix7nGn1MooST/pPmcl/ObizGfUaK/vtZCcp1TqybJn
rbSKEIGZ77C5JpuY5w50z9rhgSisYhsH4kBo4AAPIQjsT5f7wjejZjXVbZcZ2L7iet1M3vd0tW/v
SD5Vql26iZqY3kvuU02fN54uS4Vp6Fh22Emke+3beTFwIPFmx9E50jcPZ+KhurA+puqng7rl0equ
bJvumelvCYKfEqpN66b9/XLNrE6oaOgmAJL9lwJH639izI/dgBFxwzaq7i2CbPvwUYnwepqwdnMZ
kVAwPxv7IP40gE55FB3it2VWW83czxQelHwSvdvG3z2tSUbuFCtb1Cbao690Mj0L7hG79x01puVA
npL9Fz9TEMsawZSye4gIC3qW5QOhOEx+i75f08yv8s8p5euuLyblExwJjFrq3qgdFX9u2BJ63+CA
TZTwKqynEs3eVFi2TY+/MmB0DsB/c/kVXtekyf7V1I0QI+dkn2yWT6EescqCzDuMq48Ag2KsuhHZ
RYIg80inxG2B/2ZBeOXjiNVr0Het0dNxgIOmqfsusf2VZl8OuxJNs1GkEPDBlO4Qm6LrjuRpNfpQ
iwVERlv7sYW8qshYi4/KgjKc/V/BJ/8vdTJJPseM6bgVrAiuI1V7hw+F3rBryUw/H4mpGT7A8Yh7
ji0JTwkb/OhbuLCGKz06eeOShoRQdEx6yo0jwTcyv4MShL8SvOqD7GkxSHtc4GTup/0UsRD7Dgwk
5+4WmDwHdRJOI5DynNxwwC3nBCZTw2XJsEzYrAJyMcqaNu70zugejx7VfOHPwttl1/vA89FcTgOm
nonyw9GtR9cRo75nyps08fIwQmDNmJg92xDY/wKSTr7Heg4PYv+RhcFqZMjEfvoJJIxVai2e7+6M
XgdDbdC2k2dPKgQIAloGqeWxG9tQIM71P+xmIbUZDHqc8tWX1SmH+jPShqGEW0mF1wOSvYWqcuey
hTXgN6pVLzyPACD6wHmuiyFxUgVqSrIymQuX6+OUsqDxEPD1yVVLSK3CfmKUMLXrwi8g8YXUGU4e
PIOXRqclmHnbVf5ghMugETV9A5PEnrZ/GJNeCEhSDcksdvorv+zDdetMoaPCtOFmI2OdwGfqMnCB
kGy+Clgn6w9VQaBZb/RF6gS1mL1ua0E+qCtJats7AelfX7scEa+qFqyiu2KKHQX1HkhPJOrKJtiL
GplrVM8AINZx14s76Qrzg86iB9k4F6LE8oIaFHG0F64j8ynwVBvBA3oWUp6lozWhOkWx/P6sctFX
m4AdBp6KdZbBpdKeCWlGlA98mg0jtY5c42HP6CwH4O3frwwwyB5YgcYogldXs9drEDBgP73aoyym
Txaa3fFxsolBMGLcmexWO3Kbe1n7M+tupJ/wgYh+PEpEPWA1D3NE4Oq/85+6c4GESfkCHO0m9Wkw
WXRbCG12x31ES9vaW9jhno7i5d2s4/6eHR/8l1q+DTg5SXSaEiqOQs+GGXQS32wm49K1U23x0Wmt
3RLNwewdOWFDi85TtYrmWqWtRaBnq4501gt72/v6PjG/aa1PqgOhDzYGAO/NT55Hhf3Wz1ce0Zqh
+D4HW14mQocwk4OvAuUMjk0k/ymNFZ5e+nmUigeFp6UFdEn3adXhGh4dZc6nPXK7Swqu7mcCkxlu
tPsN9IPbHDqx8XRP0yfdMMZbUdEVO6Ih1T9OW4KgSiWagRx62fz4I46oczti3wSpx/AgK5/fl5Uc
4tk2+P+YVW1Z3xwg+XZQwU/Hx00QoeUtc+43c31RZIf7EesArfuNecNLSwnW2HAAR7z7B3M8fRfb
R7eEFyjeMD0R1RegNkn2KLprcyq4ssah3BARoCoCvbRYZoY34/upulK8riTtYqRTa1Ah7LbBUfyo
DcVBFfcfdPd28HHKKu1ecF0v3Ny8JVMMPFhuohHT/Y25XWrtLSkCaZjJ1d4cd6PeNEmvvl2MauFV
TkDGC+X3uG1rY290/sgAKcVA2OTf/PMDKJiknt37pJUNHydMF291UFpCgtoWXAQhwO8np3OnJcDV
Iot4ey/OYB0gz5nCxK8o0xzO+cff3FXaJShUOqmmX31kyJx8pjJyWKqnN+USZ28yNYy2qgrAiG1n
m/Zz4++waGNSb8UODgd/nL7NIf+oUvxJ9/F+lrliRyKI5W6OE63f0t9s/EIbKpn4y2hKVLfFbmIg
RoyjiCptwU+FID/rGcJENrtzEdWtdEWNVHuL6bEj1usDrXPHr7wmE6E2m9P85f0gz+g+sXS6rDni
5EN/I4CeFt3JhpxwbwBfdEJm26u4JoD4MRDH+UnfQazEL81pO9SIvNyti50PlKyLKQ8SSI6FTO8r
9Jbd3V5MhN4lAbC0+nDgq5FmuIy+sp7hHmbuHbF2aPoA7eFlqIVIHQOYrTAVTSuEIvxL4gSs9QEe
puiPK/TnYN7SKc7fI265WZUvgwARisN/12hgzNloI+EJQCSGE/stIudgdsnvQ0Z2nRbbyPBSSSyE
wNScKOHNDVr4qKcB75GN093WWkKtNjqlbj3xXj+Ujy4kKSRljLlKksBGzQS7U9Up+jkF0CkAJwDg
G6ddqeESM46clM61+R+giu0LCSOt5Ow9drGOkVb7yAeXO6dDUmiXVCrJVJV7w71FI4dRHF5eoWaT
oXOBi1czTzNKjcUIcIdNmnKTysYeRFd4CX5wiiZ2d2xcqRO28PRyVbBUWJRDj/sUhigacRnCgDdZ
Oato6LgS/Q6Ayg2BZQPj80cFD8Ja8bYAlO7NGxyIWBTvRkoiIQOZxxyKYXUt9GwwRMewxcopqxvy
JRVkBl+ipkSoVZ426chwlAXR4dmKh56hoB0Zx5RiLMzNsOy/Oql+z/o03abUmSLZ4qPyK4jzemc2
+pbshB72xa2B0hzE/L1GrWt5KsYae46STr0WV5I6fFjIPBPg5Od12uXoGO6172LAKLCwqIMnqiGU
GtT/t9ER5NCJTlaJqo0LTEyVzyv2ff5ZVU6K0CV/X4M2M9qurwgwgx3Csa21AJInHmOyGjE78zVC
wXZj8g2EUtLZxnq2VPe8r8Zbti88RcyVbenLkP+zB6EcQRk0go30qyIdvMk9Zq2tvtyut3EXn8Dc
4kIC427fwroREr/hDWPgjlCexzdYTpqXdshVvC/M8ilNdeet3Y3Yqlzn2liQaJV+vPmYNJk+wz6A
rwX7AbO7LmIdPBSDS79i+V4gnMVhznGgJtUBT1b8YhZzLlYgq1nuO9w1StgLpeIFOZDoyEaJK4nN
sW/Omj9vmDpUqZBczvImtYs8mukrVMCpDOFTb/XcT2bZnx/MrtXmML6Qo8hEKCwc2sgtBscllgK6
Ymf/RoAuUjTsiLSZOH1E+VoiRYlgLLeni4bX+1oK4fQ8m6dKgJtQ5fkkuAU3xfiDSYXVBGB2cyGT
TdKo3x73VjAruSGeVL7/RgW0vJsjK7Sfq1j3jalukGykQi+dijsY+97+NMaxtLZ940zslVh4yssb
KAJqhfkd3ZaTL96rnWq7k/fc4+sUOC41Qo9P/UsnAPkxSTF1Ja7b73eyEj8uJFy7D4oIGVT84S+j
YVFGYEG+kCNQ7uRH1e4NtmCAsCccP4kehpQWsgt8x47Y7cERZ9s7Sa2w1EoDuYvSmOes0ibl4b5t
lLdgdnt52m6BB4iHgmkxHrcG1dkJ67TWUUe/S0AsJmm83TmW2IIxWoSn35OagmmSzgZks2t+BM8p
mN651fInYhMCM58KTkHy+1+V8t5apXV+v1LhHGsyKvaqtHCZp3dtE91wQOBlcAXprQAxz7P27wM6
xgGy+hPII+F4KhyBYun1P7GPFt0CRQUblzA8mlhK/QEbw2k7+dSP1/QrcuNO7fv3c1I6EhvYDQgL
Nb2tSIJpgWr7TzY3c+zxkbo2S1RhnmAvhWjhP+8DlppbfQ+u+X9KSPtjLy2btOqiFOvH34VElzHt
TM9Ah2Q0QBwbemRfV9ERmL5UmOBwSPgiCMFoLPzcNMLvZTxFqaEYipBzQWylrLbNsx+9KUFdZmlp
KRvtBTU0OOz9LfHMVVf1TQRc1cnX9xqQNfLqfXAmZiSPvkbgV+XwxTktyvVljpY3A3Rjh1cWpjnn
yl/Xsi16hO2c7FmAXrihdcZBYPQdmCWyImVd+zG/nDrAJDkakORTblj4te9KDs7OuUxxcSwwwMwG
olS3hJeh742XHhvPklY89VE9fKrEf6CIIg81mrJdb3REdHpjXk1VqF+187fqac0kvc6KVowchLcd
UgrzS+3bcr2Ec0zL3bZpMiGcult/G79Dr/d0KRfTNWqJrob8hw2AR0fKjJcaZtEgJ4zFsCOgwXVb
ArIgD+5uacPYszdd8HYMyGKuZZC12ePwq6ejLPeNmED4GzypalMiSd+8ek7ozIqVn0IRiG1aODza
ODcTNBxhLwIwkqj27slPVrF+e2YZS/V/KHrTVtIDy86GhvrLvQToungALAW3wpkeBzztYhO+IOxx
fDzJBKOrc3n1uON3hzaEWtfp2DDi3LxS2rg+iHlmIPMT/USp8nJ91bo75fnsD4Mm98Nnw3RQ/T5u
fk9uaH+auiqpidg2+wOWywaOhqFw4X/cSFpqLzdPZZ7EvcpuyOTJty+Dg7Ejo1Zg/00pDmi+DZ+I
IAmrBNa0TUX4n+HeTOu43hwIx7Hezy0kjoY3MbZXI6wqjCFsHbuCLol0/VhDtNasvohkiNGIKug8
JhwYigkguDwVgznyktPtjL3H8DWlcz8Ql9TfTDPrgbNUCfyXldIYC37wDpfd8m401swtqHyEBWrx
FItv7LXUQ59hypHqvPjDWJjCaNPur6OPWhc8+B4GSEa1RZwQLfxVoAhAKjk7LJzdRWK5ACgOxTmx
asonv+/sPjWYYyo9qF0tJblz3uHvMaNjQlCE8SpPADyPuKdYsI3ba2Q8DMeqN/YF/Djm/ZBUQWm4
L8pFgfhvHbN3R7++afDOj1rylxONNa6E0Pdlg72GRxAeiXx3+m0fDm7ZFpsvWtr9eEpLklAncOp4
XbthgE69TG9iEJUCjspYYc9TBc5wvV7WRE8yW/ANmVwRni28Rq4fSSzhYG6M0ZaskfjmTqOzq8/N
/KgZQhAyhaNDE/oOeJD1DrNL8qElgnOlv/XyKS0WUrDKSlAId+k6+RelcGDjG321gJ1k1zLTk9Mu
B+P4KThi6NHwx4mUx7U93rhiF9Ldqmo+dQnlVIEEk59sUWTCfO+FQhSxPSK9N/g5c2AjHkA75ivN
7ni3W7DEaTEzPw9GWLecy0NUYnfYkE+PMB9Yy0O+Mo7kr1W4Xt/XVhktsCc0weYIAANXO384yGzB
omr5vyiacDCFpfz86U2KzfXhdjBFSns2jDxSmQ165PEYlXxF/YhWQoHKKRzkH33NKGFvl1jgq4KD
CeumBvStQFY7pZJI0M7oNmywP5GUtGf9nwXY38RcsoWg7s7JO/kIRXDlxIzWeVUSr7EN9sdn6/rc
wZuytWeb+NzCSqtzgnewI8P/BNqJdxXfzxrMVn7BZsR5U8pXlf0y9/xogZOo3dkvHv+lHPRS+bgM
NSFyoGGRmJSJZJDaebHiocheHkymDRGf0qmVksgQiVoVUWhX4KOzwyjm4zsifg3cgWFaPcXbRiP7
0Ey5NGD3THoQbRToRfCAtqUEc89+o1Ibj/CzuqLOvPcNcXdkQ1SOynWooTlcKcIeKGD/+QLm1eCy
cy5Zk5FkAtftsFLPUstAz/0K7GXr0cZ3IxVmrZenhw2kNuWCf6fzW276qTvVCd0XaYCNNbuCr1Ek
f5APCZQFCsaChGp7ZIIhZAbkw8MhOiJ/JhsBoHRPldXuYKnGTowpf5jG7F+SuNjdD6Ae8fRLxhin
1jA2vsMTo4ON3UBxwySm5kWzE8Czx5si4yfTF36xFkaIoE3xg+TvAr8J1wdbW8c/24G6Cn2+wNTJ
hXTxg+Rx5BsnrVR20IOjrYQJWO+UYvInw/i2bZg1kx/vqCl1RuMpRufhwE+LifL2Z8BnMv6ZWSHQ
1zHyYywMfcEYY0GWo2x1n0uz4eGJoDMnv72hHQ+Kms3mLtBrmJazWBCsghF3bBHjfGfSVd9+2GxN
jfEwtcfcVisTLGgZw3fv3b4wAC/cUfLAsd5nwcrBAu4XWWhPbNOpNGZZPptkl2V2OexGXUHgk1kq
HxqCG3n+RnWsWi7JGliicaiH6PyNvXHxrcR+jhIGNwG+vHdTdUctn4qVO86rxd6Z7n8bXSh1ByFx
P5/wriIOKGRaIpUWlMOHn8SA+LoqHdEUSREgTXStvj3zH1nMoo56y0cFHlXrBgOftWFgHDzaelvY
ikW/O32pTfOR1takk8+2cLKQub9zkdiEazzt5jq+UL/WmZyBZ/ugwWs8sz1RSCkG+2FDnHx8SD8+
9jC66e1mfI4sTJdwUH95Je8g4MaqlgtVW8TOFM5dbuEGKNqO/XdIJhx7NFCwsAwUNYcFGIdUE0tA
F55WEuJIspEX0sRAgnMZgXjwGL1c0y8eALCBFwkuNrPkIBs/+t/Oo5ikkhJWv3MPNCx5jT4E94pw
gIlZqVZfiXGQBSBveVd0CLLbNe1XVR7dZk8zEkmtS0Y5x4FP7aCIV79EBhSvWAhkEaQdzGMqmuGA
U5z+p2//CF0GV8as/2u5tq4JFIdAZdMcelNR9PZGTfOHeJ95VL48VrWIqaczZBMLPMDtG7tifcyd
LEC1TrozgdKERFxAPOhvRVwohIOVXhqGSXlnfCPo+o1IlB0Ymj7aD73Yx69mzuX84CsDodqm6v7+
faMnD5pUYCVV5xEdrSaBLmWWD0Gcz9EctT0ktfl9k+nuJQKjX5bHGZ23U4KLNUr2PcvHLCqopr0q
Rd1R1RiscbqwGcdKrswPWYrKG74nCm+nZkEKwd52eoPfC73mQ4zOEbI23mjOXpYUDM7L/54cflWc
+eh8eITTk+1b+YEL6l0K1KFQPVoQ0KBrMkiYGWZrnnTKlsVLr416Ayv+FoC+hyiLiTht0aK3Gg2W
InYlj/B1UHOgo1oLjTCWVqh2QFv9oPKh+o2lurK4my8B+SQ54vC5cNQRmsX/bAiT01Wxh4pq56wM
uoijZJMe2O7UWUazk0nRocP3yhOFpVIloFJVAImLzNySSvOQ0TFx42wNChvSGYWPAdcHKEqfPhWc
bCzofr75jLE/wh5yvn7W8gE1UF9wGc/wNxNH5INof8KEQXU3Qx93J92LkeFEUMaPc09L+Pt8AOcK
Pej5iyn8/jMApUdTPeDl4ESzCqWrWsprfYCy9yOnEXtQA3m5YMgk4aTj4kJpZK7GUln/9/MEYZrO
VLHzCJEK3l3tgxPTNKPelvkkFRcHd4q/2VUw1cAi5GdR2aT2Xp33tH2RvzHgUB03QhtN9Q3tMVLA
cTeeo3wV6v6/Mn/3NUkanBvoe/GGtrqp2jGCjilWCMsbNRxsVX+fImnXXL5y+sgEO5iFYnG4VHHu
KjvPUJ/YK7U6Ps/1MPXMufvhCRFVNLdReuCDB4AL3DPiZZqZWMG728J67PhkSzkwqd5RipFZ/A2C
PZagMBphAKQEa8FfZ/iPik/gHQrQj7jRAVAOlGScdNDhRhcssWkyZ6y+7xEkHumy+IUVgbwa5nHt
ncEXDEOsAP7n8xxf+8GdrLx2KQwek1q8IaBkW8zDvGgpwyMoBGlfiuA7TbXikw/ZhuHd4cFMVKfg
A99E5SCsNlEJvdCtXHxJCInPqw2vGRGnZ9YQ7sVQu+RnYppjAl5HfljW2IuX2M/7tzS/TgaZsXwT
X34UYjwVVRaYEDaK/TqraFpExyoF2mUTJZPdrkedLpeXqBEklgjXMoqPMYu51tes91lxu9SjGMub
TRCbgmbLHWaN7CAmUx/5j0aJNfLJASWoLXPH9JyzuglfmpMusg1OhmaiWNefzTNEuNoOOuTEOV0I
uQtuTQiKMfeEiVnstsrNMScSISUu5JhqMFbUiScXrkVNzTJk/aeBEu7b7mzSNkd03FrkrOxaq/W/
pbKnMJlnR5W4yvvI18niKBnXcjepoNXisrHwby/gOTH47Fcv6wYvZC4gJgJ1lxP4NS/Yk/6y0PTS
N6AlQCgLqotBsMbQqKtJilD+nBMzyvDXgl0cIPyLu/2D212nNsSvFc5L8lQjmbMQ7ymzDhM+a5Yz
U7HEa+k7fF98ZrBeCJjQGNjdp/K8GoAJb4A/sIKbMeFqRykag/zHG5xupg6QxhDzr7sJ7B9mOk65
OE9e3Fd6PmWz/tJD1U+TbWgr5iLaUZgLlwNOoXf+j4i/edN7PmQvzsKvcR+duEqVY5fHr4k7f1DF
sYJMYO/6cPtgwZxi2etaRmkpleHzYHxpERiMkqNNhyPYomsOCdvSpm1QeCzfIe8ocxhLjDEwkZJq
WChJTQWaB9It7j8QwnFlhrWsOTKnQzLi+s6gFvr8FrGF0bohH6hRvvbzVZL01YVnO6GJ9ZlrzP0r
tptQrOeGNlFXOQbKCzKv9YIoR2cT4SVIDNI+Msdkt7dyDGxA23Xi7512itf8Zq4YlurTziZb+rly
L6eTCMZASIY0YTc7trymF8nxOoMKb7tjSbdvR/rEYT7yYMbwWD26kOY11Dl2bJQxL3Y4/rfigHzC
R3tV42iZKOea2pmH22b5hEzxt76aAJBsSVFRXD07gSXtZ/6PeT4cHq/FWWnZrcnq4Auuwo3ra5Rt
e+OTnPbMWL8igxdqbheygUD6lP5FGBkYQx4Cv5DuQeQumngPbY8HzxsbxlIrgxmXt3gWWrjiR/d4
+nqnFaV/CG3pIx7bQfPuJsiHG8mKbTovJVvT5VMBlZCExY/Wi3/WuVrgGyJlgW8Ozrxqw9A9eGlP
B51C0WBg6WcevjJ+wCYd0+VIR8JTAqROo75uoIbQagq9LISuFP8hiN3tYaUVHUPOJztVHPx/WdIP
l6Mk6MYY6z7GGn+b54luFyzEjlxI/QXCVRYnogAZxVChbSQPoHBKQh/5jdrvOeYnMrjORNKxvKTo
ina1WIf7b0MLs6wUDSwUF1rbOMGR2xQuu1gXpHU8Not6Ij9fjaTVu1awSddEwGSn95QD2/iD+4Ad
xGFMeN/emJHdu7T9QxFqKbE1YAK9Xi3N31LWD8ZeRD948OdqIL2CNhuS+Kri5gdxj6t49JY4GfxN
RlctwY8NF7ryTaHmOmuYZ1o4yxXyPejrOsDxK3oQ0a2ezw2dUUblrc+4xUVVFM4AA2FVM57GZILG
WrYyk09JJ5Ykcb8mVTzvO0zjzZ/+W2LCqNp0dD8FE/ABbdqJhYoc3Y4qeGEkq52aR+6yAezt2h1W
OzbB+1X8OIrey1XLB6YC/pF68aEforA8BEk5Yj6gOGmnhnFeBLN5Rwl2TqAikDStTdU06HWnz8QY
9W9w8U6tg2QlPt4Rfmkts+g+mDF5w4FccKNM7JMcLs7uNdMTU4PmbiwVH8SXh57lHbADIN4rfjfQ
QWd0x3qAndokuEwp8JAAQEwWDY3elbZI0dKOaRYHzgHyExBbI8YE17btdPJ/1G2ny0ETWxajd0k5
L43yoftHHQFbWBpLSqYLu2/+N4tjrqlGw3BahMKscQg39wxKjoPKg59f1lHYp4gbp4WeyW7imPV+
U3RIwOvrmifB3J4mEFgTMZLqUEvgQX4uz/XhtbDd+gQKHDwvLw1MZT+wW9dVydA0cyu3Mv91ZdWo
jQ4YYbCFs1b/J2EyEA/uSnGN5vnuWMjGSpH1Wt36lvCFegsLpM844RaS8psh4cjq2dWI4OqtfpMU
z7IzunBO5rvUo4Imyx+sK8XIczvMsRHzZOKjO6PMeF5dK1Q40Qiz9MGWfOAV5qTSiqlhWpmPjnK+
50UnqTn/isZa/QBUZ9hAhwjd36y/B6WqDgS6sPFcexN5JQrXwlgLHopIuiojz42wzgjmm5H61WHb
n0ZDw5w0cuLF4OLIOxpL9G9P/pW18aCVxe+zvnEZb5uHZ/i5ZoGtmUcrauAYZTSI2NcWIe5Z5t3e
KWsQqA9GFBlhqM/44d6dRzDaZ8fVgjTGu6B72NrnKyItU8NfgHTUl6JgKSHVoF94gglUXN+OldeZ
kn9r43Z4O2GkxfR5aJXtslvZnkzbIuO7Bzii0NIRYvrd51SjwZSZvLT3EbPv3j4Dp2mz9uZx95wo
yH92weeB2vs/k5hx7cNWJjqAOYwLVsRJQjrV99xyLfCKdib4zZSnNEYls8KCoIRiKXAcnLZyTFs/
xuDmLI6MZ+ZUxkcP5tDBZntd5JGph5NJNvjlhKyfz5MglwIpFRUhOr1yrIF2ZCZtPV/7MZdumHW0
UsGUJLvRUECIfiNfeZLbcqSHmOviHHPsf67+RBcCXKRsuc6LUweDEnOe1rkEgivzxpu7xIVUgCnX
Xz6EW0nGkbPBfreElEN08RLo/6kQwV78TOmG0YpcTM/IYlq0yIWq1E6foYDCQu0LsYJj/fb2Phyf
QZIrAXmisWggtB42t/FRVdrZ0jzWatr6UrUuGWXZiq9ddBAYq/jQ+TOD+4CcHAotzDi55FITxdQn
iptMHm9mwQ2LSil3LP7HjgXV2eLl/BfpfNWhSakEJcqeMPi73O5B7oIqzqi33sMZW+zmupDsInc6
MbCfoMkjJgEzadyf+6c6Tfl23B8TfUuDtZcFauLhuavTcIF2lGiTGzpQOIeUo+bBmb4c5L+Phyn5
Pt6lAEULyIJ8qQfK+1t1PDqWFVVq5Gb9U0b7yfS2Tbfp/vkL3DMntDPolqAKCnO9rp6OaWxnQceK
EMAbGxitbDZSEP67DZ9txlWVUenAd5ttXOllWAhReF+GJTrjzp4AnlEI0ZeycudxyMp9j/NgIgVh
WoGjaPDhSvJNA1bQkayhhz3K/kiYEoX06tklAO58Qwdsu11WyXPaDNVEr3ZVsy0/iNzFew0+uaMh
4TgbJNQtWgo2EmY9QWKrlC3dgYl38ymgyFCoaGTs4Wng8dVFQ7Na7M5B+tBLkDmPT5wIX4XV4y+U
Vjio8TyABarjW/97qRCJByTPum6cCWvWrzjtF99NFPZ2SFlLTO3WfhnjbnL/tY6Y4JQA8tBjsoWY
PELYVFt7AuhMGZVEyy6c0kT9KiN7Fh/o2a5V5WELRYRa2RXbyZPVYUFdSWZSzzs9VPfwVLaRGZ8Z
TgWgdDsVhULODitbmTOgWS8G5f5zbVhP7x67+0vrk1pni0pTuiZ1BnTbbfIOgzoAYTnCYoQyYwgp
HV6ckFg6E4hGlFa8lOCI4sk08neBBCWuT7kcp882ROFiz1XEIxrds3+MXoedS/5uzSdBIaNT2Fcc
y2IkzIce70peNAqzH23YrhXGpF1AbzBO879xVjma6ejTz3hRru27V/wSYEvC88i2dnNeta7gdecO
gvWx71dfW7eKNk6LJT8HSKxL105c4W57AJyVVxphkxF5mZhKfkwe3l6tPKw333bbN0tcNmcDFRPr
GSLGvlg5NXWAHlzjDPvDVL72q+uoA19vpPIXxNS1q/NnTGIhNN4nYtIjN3Z29B9p6t5JgeDR8dqV
oINWl/pVdZczZ7Mrgi4EV6oB+Lm/M0/GFt4K6Ew7cCf7itBVFjhIPhfLYff/jYXBFXlgOSUXYkK0
8XnkG3COsfN20dLD1gDhifyKmJgXQSJe5Eez2tiIEzWvEReV9HyWr5lMINs2qJ+5BAgqh4/4FIsi
wMnUDIynLTTKaYqKMw2QzcEyFMBEhuhZXf0FwiRYcLKqmomLXD389vM5UZLvNzU8hjOY7dur3GGT
WnkmMg9UtwhwaVRwq3zxx5AFHUPwz1+MYOFZUmXJGY0UgIyjD1RX4QwUbpkYJ2FHMww2FDp9+oNi
npWVd3iiPzERyCaGpkkeURAAYdkQyUqo2owpe2C+LrBveqPJtR/iYQ91GBSYfvAjABDLdW20HaGY
IeRY9p/LZi6ZFRx4BBVHSLChHCXgLWAm1CdXsvml0EY49wz3i0l9E5q/D41rIV18RSOaEOxQcdKL
DItDVLbrBT5wJP7KeJjEqA/i0tnKKo21Rdc5XZKnWqY4ueVrtB6ZcCfp6NlBDKbtUHA+6GYDeAUW
qYCNDVgv6exrP97U/fkBbO5U+kMPiAa8bJ0DNS/nRWNe7k01F+Xg7z58ibqLzvm7AzPND3/WqKWA
mm1EhoxdICGSq2bn60NaOquSOtdT5jtPrsOGmcgnWwC+iOfq+nyu/V4WlvqbTAAIuQje36oZhxJ3
QRkb890cF2TRCdIYs6T1/t3yV5wEHDZfSTpdBt0GbytIHbPxyMsduMkHBBJTGuCGuk1pL9WdHmCC
Te/7bIPUVOaPuwbfjlqJYUzMuJLqyIbD3d4zHq2yPPppKlDnHfIzI52Oh5D5lbgdORm9qD7rYMeg
OoF28j44eh7Y/Zi+ijfPgFKKYW2HdAv9IoPrRdl5X6VSMr3X57G+jKnggbxlhSg0CVp1n08kz2bI
NGkHLT3UvE0+M+1jeMW6Q6JvMZ8xdZcswjL/mk/Y4qvx/3RQqpGbB2Y52bWtQ00ZqX2+R9jzAXDu
sLKgxT19gapHjWfFvO2lNt8DCx8isyVs9bgUtNXYGTV0eMel3oCvKv1WnoEbttuT7sEW4tnJEcA8
a04XM/tRsU+lDslFod2wtFMkfEp+k3v3sgKdF00q7WFKXVb3l65o6Loaa7umje24bZg6xQvgiIog
OriDek7UFTe3ZB9LExNsVo+57iKVVWYfd/GndYF12JQNLMQVkP9yVsp2LQ5khCdjexNL7XA7EU6o
lG3jKKgxZT1Y6x2NFVnl9SNA1T2svvqN3t0htL1pA4Q67JvIAOcF1FwskXpQhFLpecE0atW0C1Fs
jWW9/isHKFY6di9FPBl9MNyipffwCCQhVVCqDErbm8j7rzhyK9Gjky7SAVn3RvE4zlrRdPsb0Ew/
DUn9Oywkdof/Dr4jLn5X0W97bj3yJj/Co4vcHByRpcKXLIFoZ3MHyP0VVDWB3YOrazNzpOolSVbm
Xpqz8UP0NbftJN/3jhwW68zWkwRguxztcGwAlhPCEcJ+OxFMD9ANBnyvNP+CFOLcMi628TunuaTz
qcH8Wy7fIiD3XcYjc7630T0vlLN1VUbIxi6TJAMeOXz2qvKdQfl4vtcaoe6INN6piC2pgE58Z/gy
etyU15QVpUMDOlGZzpUoQOId0qNrktnQ58/iUCsv3O9U9e12BiFu6gBqwLl6EUDnYZbn40xzrMtN
zJnpcKMv1h2/Hj+1RdxGbxD8VrfJ81Zi23f501dv/1JyVHxeFbX57M4B6Z1x/6RfR8Xc/ZCoA2SJ
QsZOIDUCuiMd5xn9N1Bqcl9iOV4mXz89MJz0SN/HriHrycZGIuyWw+TH70OA3hzpqZ/YffFCe341
kpGMTlVrl7pboB/1pkoii0AxxxighsS+WyAXklbjlUxGackMFwPtlMnywlOTyH7e2YXml3b0g/b2
dyOfcJJoRWV4bRL8wgpX1Ef/NeJKm2kWXbP26bPqPyxKR4BLLUH9i4Sh0J1T5U4zZZQlA/VkjI8Y
DnL1nHdvEOxzmd9WDDmR+f0DklCcLw2fwu9tZtaJVIV/Nb87x1jB5z/dBVGCQ8eWywNtiVvtDHQ3
RKnRaYG1oi3m5AXDlwSsxL+45h8LMkRkCPQvSSiBFAnN9W5Rd7Ipjadec7mKjHT7Hl7ShX3d6cFi
rv+yV2NCA3eP0y+weJYjpCwOpptQDAUx1JrY8EkwSVWKAaCH85HQthTU1qRE/e1GFQ47ld0hwG4p
hPJtp8iHC2ycc+ifkigMg561Z7AuDlSrqoWCWAoKKCnPrEs+HwytzayeTjFv2SV3OlCLlPYCOzj3
EBJSj1SDmRYwjKp2RnUGKtqiqAG/vtDYS6RPe+PfZDUxvcC+t++M8+kpy0fNe6kFF1+yp3mRSW+O
XznhAQl7/a+KsHdpXU3XIfTgUH/uBPpIJ7uXacvyJZxJx1B1RLYVLyj49ANU42hGXlq1WUHCeeE/
Vz2TVbBra/A9WmdGfWKp0OLM8Pr8XznQRixVa3hcQQem4gLVLg0EQkdoDIZ790lsV32xEkr3Y8BM
xxX42OD6bJUsaYF06Bbvfzidue3PBOwHQkiXKxfw1tkbl61iE1T7CwdRQ7u5kqnr7XgTHf6GMG+x
fwoHAQy861MXHgbZQPEWrzOVFgMql0jp0ailZasSxudJ4oNTqybQTaq+/3dkofVlfrb2cle/c4Tr
TeiS5MTPf5rUqyqk5GwmzqKUktjBPgpuSIS5Lf/RbKRfH4LdunPHl3fepDwAhwL8iQFRsc3txt69
NT8GQMZXkNHdTVakUOfn9gt9I9xQsjp++YJtO/6dZgJn2DGM+6e3AdtDaV8LGlZ/CQx7TedmXWgm
XaK0NMiYi2xjyxu9SeGc7D2GPKrc7XLfSM6GmTeqRN/IrUaFD4dXtd9yeMel42yo1x5QZhdvpgmX
I34Q4CzOUL+WzjoNRBGmLd4qc5yMZH/J26fBnM5ikOrGhaHQpF6n4Ja/sA1GCaDHWksmF4i6Z++g
drQF2XQSIiW+ymXdYf3UNDTql7pVJz0qS5UERmsPawB0YH9rAWEg6oRqP8zkfTO6Sbs7hE/c7fFc
w9r9IJSoewWGGGGGckhb+C7bkgj9XOkWeCxhGRGNveApGcfVU1h11xmavUCy+EFu9GV4XpA+ajyw
3VhkIuw0LsX/H6SCS2Ld+E7XU6+3dlZAHBvD4q5CZzAiNcX86pm552ID81r5Ia7LtLE7i/iFT0ig
VazSFVhBqb0DB8bWDsZE3AgfH0wvxZwOzdGHSuId4+qHlhVJCcPL9XLRhNrtgG0rze06zRXxscTc
VSfR3YHw25Bfc9Ki4pOR9z1Ccq4tCz8JwgDJd7ZljzgM2Rbu+6AlSkhCL8H9EkJ6Bkxt/SW7Drvo
/D97KP598EVSeld9OL6dT+zHgTB1xF9JBnc6KnO9mNx3OyDt+pio3BLTT2kXLa0LjFbxJgeR+1vj
FbNEOW30LzLFjl+TEPRWj0AeFAuv4QyY0X+XjXo/A2L57DTC+bsaLoo3EF5BHJgRMMrVj8MUYnnJ
g2A28MHUmBs59NYHWVcRzAcoAAPRXs37eHSFtSg4rkClg8BIh96YV45q+EjhZGEj0oB717euwfmr
3S2r0k7MLivqusTrvzN4UcyLQcOKP6Q+jPsBy4MpGuICYNkpqw7gaz+UE7lbtm1Fcx5A8YAfUeLg
LS3CoS6BIyhUlPx2rUW8nOryGwa3qW1jVlXaF9AlGq9vKgsN+9YlWO8cd2T2vcz2RU+N5ysTtey5
ztnhgfF2jdi+V9MTEyEHQlowMvyLsaS1GIhtUB1cqufrUwpemUbCEAKAYpAc1ohwUKWYsncrsD7T
VKWqmSzfPryWHSlBCyqhrGpheQzWbDNrIaYMbnzQ8v8e2c5Bh66jyslvGywkPoFQ3tzSe41P+Jgw
7szLEJbzYIHiuMDPZTwxZeoCcKAH9NVz0lSpaYmudO/nGwR6ASjTXgSQo3Ou82Jvg25i0mVm8c4J
L3dvQfAKSNh/nr60XElOIAm4NNzk0mZFG4X4xKfkQ3fKbH/ftVuGHjGAjBixT99f4PC5cCXrW/FX
jdvYkerbcLYR5zYUe+S9iFZBFZ0bBygZLRr3v4NzH5aoiKgc5DVJtHlAmZsf1jBiDCZFVFwmUumz
MZp97A8J4s5noopzPpkoIMN3lUsFIOhubdDsqht1ufIp6rTR7JdkNrXFE8P/C45s/dcnVW4qVf3o
fgXL2NaSixBsBx2FbpIpXkURUey82n+j+Bnh97WWrT84XiFfaUycfWlDKA+EdoiP0ZRWQ0UIwte6
osELt52vmhMarZsospUexuCnJNy5Dag1u02irceJYOVffqgU4MqX/rrVWeqNTd3lX2uT1A1hp1YP
y2ewXh0/RtL0BAFSwQoloXxOa9mFNwFqi6IK8zVMnctODMZab6gpp6aRDPP6uIdY8dZ87OZA+MeF
0vyu8R/+e9Qm8qid7xDuxGDpW/jUDCGv202JGGk8/qF5Xy1UDyHUazVg0aHNtbjxZMKJLtIwm67Z
VG10uesd/KrxTWvFZnty3iUo6ptVztM1sDJp3k+qHo8obo+aTjyNICllaOCJJCDV5sBcdWyBhYav
Jw7C9FIteNgyxnlBY0NAYZi2V3b7uH5P70jvXVCVXNAFFoH0JUyuahuhPXDkLnbDYGd14dr+FAGp
xTKVRTi0PZFd+LvtP/62Cu3qZMCCv787oejYyZA7bqMmJt9YHCsz8MFQq4D/qzHUqkzV4n35xlU0
li5I+wJfVEclOW55vjOgo+nMSOM/YnT10xhZUoBjhvyUcyObVW/V+H2MoQE+KnHyuR3Cc0vMf82y
SDzW3RR9jN8nzxc1xRfx5C8BoEnIQsNK3dTlu+VUX6ogEyNQSj0lYHJyAqrQLt4Ht0I5WZeddkhP
5AX1HolWYDrwciX8A5cT7U0/o2Omb+ic2Msor12t4Whj1R41CZ66zcrHmvxq6HS32OmBkQc3UaT7
alTgWV6fVcomXzedKQoDr+1oslnOQGMgkHx44twkBJXHOTmD3W3PZbpvDmFPa0veZZlDIsRFlCgc
7pjOhJ9m58gDfkVGaDZ8OGq/E2zFWuEBSbBRc9tQir1WN4/0GOyA3soLKJ2PL6Q/IPp9xz39thXO
2J2EonPAZ2pFLiohj/VDRDWBN0lGc1Z2Y8thhEgFIaejHRmLMCgGSmTrXGTxeBSaq+K4GCNsLAEw
95muQUafk/Ur9IOVcRiTnTkhopxDXR5v/TnyPTW4FDEDr7r4RKcXMnamNBkAA8RvDAC4b+ICavWB
Dh6Q/8FjuBfdIYdjufvAxuQWaAXvfamrsXS1YdUOgZXs6oyR1A1/qcjtdmNRYADve+carH9dQvp7
lrzfGXUFt/5t/tT8hg5ZmpUEV0mml/8L21o8pgY6vPog4idmDCi/J0a3fn5dphZwTlmJ1KlJbWHm
qyKcctGLeqTuLWY3LUJCVRxM2uhjADRT9gD1i08hpSmVSgvUWCbxr/iecqle54v942Tb8hDbYb8r
2sPp0eOzn1r6oOYTrhN1BSrgGaEP3C/KodZl45PcL+bBnlVIU2qceyUBztSPV/1LRLYBzaAma4yT
P85IcXNhuCwLZF7eOEQ3b5kz8ZEOYavmm3WwRn6uNqbdYUCXJ8oTtlBrBZrwyOeR3V0z2bnkt7EI
0aJ8mHrUgPLZe251zZ6xNa0FIkSunqH3Pss2djd12koEJScbQpdp92GMHnhPrrfg/Jl93YlPIgw3
CO7YpIb9JpCHfYMfscEZEysdXeQJy4xIG0edA5q0BEuVYgdniDojsVleVdBrUQEUY9OjTF+razCi
hBEFDlLCpaIX7mCpXTZ9AC8BgoOvP2D3f2Bs3FtlVgNAHXhI2P96FN4/pbEyQfy8ZTWkaCMAbT8t
F68e6zZS54L/us2qBEggvsOAw/TyhxRJ1EF9XeHLeDc+pw48KKG608581mPUrSLdYphyTHo8/lC5
1K2aAr3TJqfysVY3tWVWr444ThObZi/FvzH5YD7HIwwE6C1/eGX/yj9Ns5+PTIFIqpCnl+AV57Tw
ZOWhg80PAdPnPdWDLDDJvQizM8w5BUKromIB//zQgo63Ztg/T+N8MRhNG0+d2HzCllbltB+1bljL
j44EYkwWzWAuMURDYkQw6VMGJF/HXK8w5NYmKj6dw7GsCe44ACR6ilVklRB/ekjYgJntHKQFolSC
nGhcIVYhDVgX0+gnR0JG0hHgE4PFSCoYpLJt4/srLqFr9p3ATc2EVbr5B7klmYiIHkdhz1wQcJMR
N5V7RbQeV48avVP1KPAX/TUGO2tvrtNK6aGZy4bqWDGDcmQ+r7sGuJdEZEBrMPNRDaB6M758WVzQ
8sxmxVxk2zB/FT+/Cx3XaUbmxtZtydLnOokks7aOnHKnokoN/5jBeWTm7o4Eq5GXWgn4CFGKe8HF
rKtGHz7ygrOWdBqGG3+AKFJBauwUUlB92eupOWalwdRG8sOuaAYz5RKVJTdhTiUcchw9ia84quDT
TyGKGg3A+CmT4YAHcliGMtxwd0kISrTI4KKqVtsIeDcTXrs/j93bzj1JYz41itlDZhjIihr/I4S+
ABqsRdCHk52fAwbYd0TOYUUeGbFjXr0Hh5dykU8uc727e3CN52SpY2bENuW2KOsEX+fMj/sTtVuG
6l7U8jLnX1WS2wlIEiqdO/bWcCT1c2vU/QtBWDldTnmsK13vxThP8jMAEAcNosawrm6a5dreaxHh
Fsjo4+IzXWxuC/GhOUi91xVO8x5icEl5wwQ/nbwnklRxxX5Pd6gEUvHtQbvhqhKcpry8xGsfAkdY
r7VoHMcwchXS/J0KahMGZxam+oybjpiAHl22pMr7Z4o8JkXlyHm4qbs5HXTHxu+1FRPtMrTcVxYc
4SgGXKpcennrwAj3+Wcdr7hTV4AQiiiWUUxQ2MGMs2xNiNyXts1olK7z1xY0VKa1cQcgf7DY1lYW
KK2Bw/QDHXOaLb0AY1hW0hOFYpZNheOeklTohy5SbwLOpL4A/MQrNPOPyLDQy43fJAf9Cl5i9HYY
Ce4kcPuWwhy6oOB61mUWtB3BBk3Yr8yPrtrNf4zcJjxXWl0uoPi6bb3/f0QbTpoC/r5xWEg7hW5Q
EcmMa/40fKYMlPFnnSDTG8/roNaG4zRlSEMntDxELUZfVeiFmEQxPUH/3rTkO098H55x7Rs+E/oh
5rRvMsuDydVOewZgU0GKJAXrJN60dgoAApTjTcOpjRuiypqoSuO9oR/Fe91A9Hy5eTnn7b32hMO+
BU3PsErDehV9Y//brsUTdKfrB8agibGpoKzzVrRvFCMYUuEDgCdFvB/Ry8J4RoA49coEqmecoV+z
kh9iuqiz6iKFwF3Qf87nfMMoyj0SsQFWJCUdUUYMenQfGH/Lv65S+E+aQi1Wexop/qJjLLl9Wusa
3251Q+n90wF6TBflc+dAKSDsSXmiZ3cawvR4ePf1Qw9+es1HM+GQtoxFgJZHh1X7dxyfN35zTOEZ
EfUPhl6zVl/rbYYkBoKJhxALs1XNJE6O6QjE8ST5P4jUgn+hXN2Eo1zz2QLD2AX8DtTUuUdiXywY
FLeroLrnIRp8YlhRqkxda6S41HZGaLzC9F4O9mEh7RR3+vxJFK66zZFpwxG8iqUalzGI5UuKpddd
KH2eM7wfRZkuixd9KnXQISvgFPAymQoPGKs+S5DhSRKNUGoZXjN9/ISC6DFwdMFGEiT6B49nrnbj
Z0hMd/odJviMe0nl5xl97LG4dp4GONi8SUxBqWK5iYsgvygAdw7cMqkTRyIIbJRHPEpoTPdSRKPz
sIJen8HnhEYfYZDznISPIWaqyDfuhq/jDZvk7Yh+vlr6JnwkqmUOqn0I8waMFwWQG+oPGBcnlS3H
hH2b06FZ4l6b9z5c6RDrc9mH44WkHXITB5lyZKjW+io4dQ1EddTwGyY5FqqzOLAsHOBOjaRB4bnO
5WNhqGs8tMsksfWQtwf+ZE1z4/dw/O4yd79cw7HlFbwsR6BgPO5TzqqV8N0oA5OVA+Cichqju8Nv
WO7hTdr+mGowp+1XGU9ZZuWvFsYBQpJ53fVSu9KeBJqJ5CoVMD7HfjFphkhGY5THK+h7EK/KxoOh
RRkzYgFxDXNqKNvtF1StGuxnFkVeUF3Fc6ZNUlZT1yj3QsTAR3ZIxgKK6N2JTsKB8q9bQr+gVM3B
L9u9dRUIBRWP3DI2hYqeSjnUnru/sB1UMoFS47ILAkbf8SK7w9vOqktvgzoH+SlqcFiIifrjDmdg
U7K75wdgB+bWbzRm+QcQMJNFpsa6nwtLB66ESiHsYeNBBU6L+LvYbg9ypiF/ERDjdlcIIZ0iHx0s
pobF0ijDtTITBpJtSWkAQIeRfZ3lrnFM/WFYXyZT6ZD3TZi7/0D7f0jozjWeJ5BHQTT4fjfkWOB2
3EhcBhdoWUIDJCu6Pt0+ZkH50w5WenUT6hOnbsqN19M/2awzaQOotG5zcBuz61//rAYui4WRmlbr
HAcKX+gYvH0cHob5XjUO+TGPnSXJfFD3mB8UZFcX7zVjkPZOn1k/m3B1pwXlEfstpCsbwY/SHoY9
QaOFxbeStMvbnBMZon/qGiHCazWKDlXD1WvxD/aVprKTnDCwrxlQmCbes05OlfrtlZqNC8wlPDcy
0jm6VWE2CgrwEyCCL0zbPCo4yPCygA+gMkVa8aCiEYlJo/AWoCSbpAN2v2VMyOH3OYnxzjiZ7M5q
c2XE58xKyyqBwnUoAqNL3e+8rFZw9GScAZpsmKrrB64mULoE6N6evanjeXOKNEPyZT3I4ixy1Oyd
FDtsq3m5Vq8J4ze8YE3IXRe/mCb+K2eMer4v2lda1V1uvCBkwVn/kET4XEyTK5dBvX+L1VJet44I
iURC8U8EPEMwzjZXIUdWxJRyb4R8ggrga7IM4q+t1hAnFlOFqWpGFdomC/dH3hWWuQGM9gMDVjEt
XHit3424Y3LTZGzRcz/bI3dany9+4ijxwhS5NdonQNHN4J6Oe+gqQyA05ZEKIK/wwCUvDq6cy49L
7OeXyRAU8MYTcB70P4G8poeVD6/jgI2usheX2u9vHbYAQgUbsh/6Ui+2h03ECgipco9kA7j8UTkz
G095P0V7McSmxWddwynnoH53RfdkvM/3qvIYiEeVodZu+GrbbVPz3NtmMNg0jMdMdXi+dzVCJ1+/
4Nwx60fL69O+zAAP1m1YDrq8H5/DanJbz1uQXYix5DbZxQ/RWEu4rwUQnpzMVvED7jzsBCS4a/PY
b5o+U/itqCDELQ5vENYkmDddZ9A2cFE1/grYnvS0dFM+Gi6DuQeHMtG1tH7v9Gpd8a2a9n0+CoxX
eadikCeyuDFmTe4/5W6XV844CnOGWTYPLAho5aXFNmgjAeZu1HrUfehX2pLhLCim90TdAczz0ZMv
IxkLLg8L4vxKphVl5laMs2Cdw7qm46c11RT3K4dIYelhocylRjfQ4wrmIsw7eSwIL3FcQAP5bJpF
OXfJ/eRtH2ilvVTEy8pyb7kHLMPoY1ZgkRASbH9dvEGON7UD9g3YM/OYJxwHV+LlU/ubJ0+FBkcg
toaq0ldk+x8bBBP0Z/93euPXnXaclTwL5RZf8gKNCqt7SqpYaS1gDrt2nuKOogIpwCsZGsPBkSKT
fj4Kfzcmlr/hzVhP9A2ulN+ltS+XKqvBF59hSSzsQngrEQTC0aF/wrzVj7B3XEBOvFqRwqzuwzCW
rNqOnqATNkq+LgAbfMXMDQtFN0tmO71PSIHm4CSJvSOhgMzmzoEvoH1taUFFEiu7BBnx27prwvS0
Ug04QQoggumEzELBOrvUGCCyHTLJBCc3jTfWvvV4TkGNK0eVtRt/QGfTpwb35w629vKHXupJ7Ccn
5uYlhM2+hjq4Uc1xKP1888pS69x0/JNBZ/7W12WxxpzmQESeNjKg8xXEI737AnN77V/AMPHX6QG1
mA0Jt8G2fhNfqLlgCafSujl7y6XVfODm3cSdVCWdQIYNRT+oC4esiP8LRKUXyGtmj1KEKW80Oxo1
S0HFN2oKJx7hSI2r6vVCvOxTdMd+ZdoF+0ljbDV+6FsNC5p+Dmcvlp3tEVbH+aM+5clPGTndIcNZ
vGMK6f0qikP/5VVaUyfMC9wlhWxT8sV6QR5y9doTmr/SO9e+/FNS42HlMGYwG8UB4g6wBHleoH6k
aBJk9wdeP9nSekKvuMtYllBHhw/h6j78kbgfDxbrlnm5S4Acuq0suUg+UMF+835HyNWIsWB+EnZi
AHS1563aJ64SOo5tj24g+lxC3Fgb/A+UPFytmztmO1oVrjf3e0QeTtf2MtEioNgEUONsJ9M3ADiJ
ZF9zC847bQMtOupDmagRcBWtJ7sUG/mMq59z6DC6Gj9c9dd2DDRa2cu5vwvQiw+E0bRl42S8ke0W
TCjkovZaS7z6cCrQKD9YlSJEmOV/eNOQbU7JLaWLwsTNDYwMvkgwTeeXw0GBCBtHn5sDhUOyUhIt
XVdVPYHRGNAYrZxb/1pS7sRKk2UnfTsRIKn7WOKMIGisVYtTDSQ/xPBLsNW1Ew/r6n4hzZ2On8zz
HXQttUPnYmoGKsso2w9VoGf+8pYNQCl+wwwD7jRz50Zt57Z7sMSDGR132b1Fh9JVi4XsbEULPqN2
7EJAJCYXQEBD8f6s1HWUr7YeReSfPcJjptmLBf5th3Nw3Tgc/bqHRE52O1jBjOtcMMu6S61GyWwJ
MuyrQMz7QnO9eJvi8GdmXcUWAX8KZzd0E1vYQIzTh+MG0qI9QLkMrAnPCLvhxXq/JgplOe+GZSWJ
RSIQPXzHYhdCY/uzeoGjvXZahOHfVQ+Srarr8JcOw2+s0loB91rNtSvtHTWVYp5KS4gHWh7jrFA2
GdKykI7AANGP2RwdmG5qfs9zoXJPLVpc52EF+ehgwEH+MLPESLY4i19nj8FeYBWVI218XFK5gcBq
xr/9/eOWttf2aoGcdv59D3Fq1NrGxlWwaLgSLziLaz8xrJr87GT8LCR718Cmfv6Ye14mGnFjx+vh
IWSDN+uJ+QX5drI/kwfyrVIoTGFYI/D2xT0ftGUhvtO6gOw7XtZugRghEKafMM+AN3iSwAhWQMoJ
PfRYxCI9aOmdtndO/1nP2b5ykwO3HMu/pbeqcJ/OfqoBI0mfLI0Zz6kvsIIRs0v0Uq/VQWDv/Oyo
+SChmvrN3un51WKhj0+1zNM9GM/NTtXMBjPvBE/ulA8nSawKKkd6hWsT345rBQC37vrpvRrVODPQ
GtIiJTWiL4Wq1Xs1GGTZ339xe9j2d5LvdZf+HSAY10IGQBTPzTzGUaAPD0QpfFZT8inEXH9UsGtI
upBx8Uj3+nWDP+5zxWku56aqUokHUirtZf4sQ0JeOAtwXVpipwocTwoze7gz8OTqIzVSb7rwyKS0
JMez5NjUCSMUpd5/1cnkt1TprQFFOYh/MEJLDYPIdlAiRq5G2+D3UKUZDnlLpaRMPgUZuVzjR38l
AEeUqHitoZFaul/dfjF387ZiEFHDy63Q0n6F+6uAUw0gWpvH3f5WvGzx/cAimBuavIT/Ue24jZiO
dezgQr75CO6U41wjuU0CjEOz2u0I6rNXqgXYdheUQvc5zOYatp0GavbRwowMbBjgJIpDdDiqxsu8
SfvYioZ+vmWflus70zLWiYpmr8zONXMKxpjDXCWqXbUNT+3fMALJE/twrqJkcTdQgFU8r8QHY+va
PqbwJIv3Pwf72Czwvap0a4HatcZhFV7Sjb3L2S9FkaOeB3dSLrad4GTcNULp6nHk7NSCO2Eawj1S
XAdozZfTU782NENcKhY1uIBLNlZxB4jbhQo8/UxHXpJAlhr1oQSkx8ctv26UhF7uUJ4cxIDRqZKm
DDwYmnTYEHymurA31MD+hRWmtNXeSiOj5tUgLWDl+/XOleLPKEcKYiyymQjohR6sGoSlczDW8Uct
03QJ9U+inWJhwJExoCwHErSV96z15DgEdkLbACEMHzZKVA8HkDlLbsK74OvQcpwQ4TcX7BJSNd0i
dXvmzl1kct2QfIG0hU+t3IRgPRFz7NZCHBsu0jW2HFJL7qzS5Sq0kBSXg4fOJSH7QrZhpvV/D5+M
gwaAiuZoF2UUFobpnOFVkakjzQclyap4tYmWKK68QMou5ntgNOC9zdOoc+wiZR8xivbtZxCiy1Hh
Wi5VDVhO5Xh36lUNV9760WKsMG2KzltRf7flOD+wamkKHkiux6pH6l343LkbQJ18C6Ns2qrQdDKD
gc7ON1rjZweMfm0WWlPVsT6Msrf933sYp4rvL/75s5mcAXAL3gTljlIxt0jKscPmgelWmfs7CHcM
el5v0wWQwyKY7376/LGs6VhBsmTSklWb3sQnLOddNVZXcxcBt7FOcs+CBx1wFOuAoDE71Aw47tEz
wGCyCYcAidYfly9wZnQfi7+OuKbFHT3wP9+gJivKEp+4v7jxZsfWP6MEQe0bCMeVIHjkFZHVOdvc
K2mGxe8cS4RzutgYKFoYPB0CAc3vsSY1GLWNALqUxPxRJVAQjFAxU6sDJYEvi5MEssYQHOFv0GVN
R/D6OUqEP2uMcM3DQpDZe0veWtVlu4LTl1hxe0FOiPv1Y7+hJ+UiB+CnhjElZ5xtAOP0YmuFxwxa
wthKMcaQMNgOdVnbrC3F+t6oaCOgAKxBtk+tLF6iVwoKwP8GJY6Hms77YHq8bSKW3cj5xn/tIrfL
iPSFhJfh6EWG+Gt/Mc3Ga2scYB9P3w1c/MHwLYOKFQ+3cL4kcCJWyNS4yAtrLxfwvqUZmdseQNk7
5TrychH/JcmjY/Ryu+Gv68hVCiunhBrYG0O+/kgQv4L1rd7RMEkra82P4Mv47FmOjiJ25jD9wvIG
31h6m6zKAVH9WvXh+rXttaMAGBoQ8U/ct36ox9wMHpW8FEfMSClaxMxLsKwpnJd6XnSwgl6vx1ch
aiTkTpRmQqcySTptixBzrR9lEcHz+tY06pu3che5k/RnLOrr0Fon4Pt2QYH0SRoK8JStCX/WVZyE
hHQ7dmGhv0+dR72VUoNY8lBHTHvrKOY7FRyPQSuwNp/W4HsmKkrHVMLhKb/epP0ugSTwdjtDhzmu
0IZdwMnlXi/tBQmMacu8W4qVbkgctrG6fMaNnyo9Wx8CRKv/jQ5m5AMgzNzEn0pKPnzImLFOgGm5
zrUXB8+tEjA6vHVg6we8TqGzkHbGtXK2Iu9IawM8rH6K2c40GqcJCXFdvl1MIB0tJV8h1tPJzryZ
jfd1FglHySn42mv+QuDzh/m97Kr75ZnbO7R/NMo+FnRlu0CmUdiiX7oWjcbJZLKWc8FhxNBNx28z
O0c41kRu+cCBOou6T0LLMfF0FWaY1JbkWvMQb9+vihHJULPSOVoew4jH0gbX8M6J2j7Pj2tJLZpv
MFY0mOfvawpBfZI3K+qtD1nC9C0HbezhYlM9JLaIZyBXUYrM3m4UJnCtr+wj6XcYzJM7Lwxq0gog
9AqAPvy5DqisqUJCuRVu6turhYsK4A8/kD6fABF5BKZlEtAEmQjReugTlOwQqHq0ZQby/XHH61/+
6jlbVVzJwcflqTIQZkfGyYdBjrOVXHB1YCKsI9poSC6OFDIhID9l6w6pIDUMnh3Ura3i3b5PMd2L
mDnldf0UxdunDz5qzfEFDsetlhAj51YdtFQy5o4N2Jv/rbrw99GsBEmpORGn6BKtCzMdyt57/y2t
gIxr6yvd8icacYEUrI2wBjd5k5vzyEjW5///1YmV45FdUlR8hC6TbkY6O0ZJWJjhpTjvJvAxDJ6V
ifY5BYzs5fKp04AUagob7MMTyIs7Xfn9H9uJ3IEwMvJqU7zQCC7O4q32AhworJHFCmHQzjYmvyF9
F3ZxDZgr2OyLaih0c7RmqoC63Fk6UHEzQ8UUnbPI7S9ieoHrjEmG0CP7/F2+bVirg3giJhqF2nv4
Uwpg+PmuUtzTBxs4laYlH+bCNHmdMiviFSRJY5a36TYP0DJcNPEP/XCUkGIjH4Fd7HYSDxtNOlou
rF0YlQwfkcF7qoB/3wnYH0ZfErZjC9OQrYpUW3ApJReofWYU829Q5/shlr4281ImE/rxCf0T2T10
UdNoeivM0tzqFcBnpzVa8/gGztYbzekHQzVW4VrEPSWXKmDbTPgTASmsklv5Z867IphRSdWXEl+v
S8kyCHDPxfbuUuIRMUAg0QGLXoGq98MZsXuEfe50836eo5ULu063lCVt3PHUa9COepqv0XyMRLMu
SVzuK7fbiELWW5rS+mjUgOvUs2Fzy4CnSzzoOBoFlOJFgHGsiSNNHPJXmGAzb914BLPyeOivWylg
KE2arijtgmckOBSO0TlWZCDAGnPAR08Y5Vwmk516x0JsYvOo0hpeA0VSCr+GgTm8EhRgmvpdKBfa
DhAIDfQP4/D+n+O00egQfKUybKc1iUeUXyg+f1/VJe0gxLjAUKx1RWgT0OcJiZjAyobyS484P1bR
fT5vUKRN/+e2fTuUfhDSdPyeR7FdCairjzp2yEre6d9xZq9OO8duw0uThjkwHRzOk69LiLli4n2J
dBxS80WaSbkfC4MCnwRNJZFDJuSwt+Afnlcv7URbUwyu+IH93ZhHmGtW7kw1NHnknVeCmeJzWXGf
YquQv2RHuuW/2VzG46lvMjc490EGZxyBitsDu5+UJdeRJnHuYk9rDVyHYD0EqZTyAD/dARAZsaxb
jt92nvTpnykWZ+RRXjCrnO1H4R93rftRrON1o1SvFwD2XIc5LMGOIamxwkOT27q17yH9H6PO6Za4
Ovl56dflY0sDp3Zhc2NJX3mvTlRFJFiB63zTJwx1JM/z3MBafDX8lLJ98rPbodNpnJMd69eyaV17
R5XfKM75Ndl6pN9H2/CUCCwhKIWuAtb2Ml4BIF/T8sYvqckWHqoPyKoN3B31yM6kQQVvHKFaF3xG
4+QMd5Kn7ptdQiLt06G16coRZEwZ5I8yoQRBUaWD2kJ+JfwKkRKoCXK3mTNNt5EwXtWVSZxkKHLq
+R6jf+sPbLfbZAltfqhnGNtngbN/0cgvhfiAMLBM9eKSMmi1MuEajDOFBA6I4O+L+tjnwzIxWtNa
XznrDhv8+YQGTgmSG0PbZHonzrwPw58NF32fz+hPZ2JVWVTeqMupjKvyhAptUjE96Z/pYlGro727
BJPccRwqSAC+Y0ngXwjJN75gr8OoC30KR4WiTgry4WkKZYnNFsdkBWSE6FbOtA3dkGir83y9PMVg
C76luA4PfE65kJaImkPEB9RHSJyU/N7/wA9uvIPYjp6q0AhssVm7KwQyii0b0VuqFFGe/XtNDCNu
l27X1J0JwLktVg+2lyC/pENISgDAncEpssc18+2YLPseSk7gNIUtUzwVhTLgsyfo/LaNoK/Ubrw/
dEky4lw39kW4dZnQ2x2+ffPsxJ7iMtbRkdKkxULARpPz5eYL8kSVBNlNYbh7+EEqvgzJoso4W3ew
GhUaOgJG/tpCEt0QClaey4rUzgVN90HbjHG1ur7gDhJebUpzs74Rl09Egxksp84c7BsvAb2fldqQ
egTRSx6PPmT/BqxQwgM4WbP9v0kbeEjvzrbsW2sSgRhXXaL3491gEqunAeoxXBxKUQcIsn6qjRyH
uY9gOU7mnKq9rNgFqkgxgvZ512HGfVqWtCOQ06TZHm6rAueDIfq5b97Znto6RW+mwpFPZQ7gEXpC
hBngeLYJYbChbkZkxQcVjlSGlMgSUCO+U2MfccC7nGKP9e97TbjIM4Ij8eQ3g1iZwWxq/eHwYcik
QqPtEyu9qPyo/rksC9oG1ceQD+2c4OBuou1Dn0P3AW98HDzP+fGZsoGciKy5zVIMtrZm3pSf5GPl
2tvUWsPvHVD/sg1o9XW9JYMXfn9bJ6+tDVhkNs37u4/C7UbCDRYF42iT+1L1Xk/IwlyJ4ICEsTrK
Ojf9e2T990QFMFojiv5DBsbOk2Tx0jUbFRikAMsbkTVMvKxbIeAJHSqsQiDORF2qFqEjmBbiNj4Q
hTgTCYF8B9nSaXvEsjEidm5Z5/URIBS2P/sNVgEnKadRV3nSdccvLFB9rsfHYO5b6YlYXxh0L6FE
L/vAmoMrVSvFEBQAq3cnFasnJpEUFQU2DM381On+H6upYL7HRk10HnGDTzqQfpaEiVWgrMVNqI9o
eXsQiodwfdhS4RMZ+sUPsBVbD5laxq5Hs1HbXKXTw6gVEBCVSRswYmhT91tH9OhgCcjDZtbITSEm
X3NrWj1E3cGc2EoSxXn8YvrGshgz7Hp82KrnfxC/KSsJtM5QnWESjmhvbDtsl+HN41T0huijwK5N
ST9YMpk1Xm4Hac1BBqSsAAVhAsN122sR1vr9EnakK4E+fEPsmV5PK8/R69ChewzvRBeVQgZXmXnh
JZ469wstVGH1LgxKjxBukJhqENEvN+5vA+1VBh/XCgODlcf7lWAJE4XcUVyg5PJQlfegvUNAs91I
IRkqvvjcBqraABcTnr+ZeUyjJd+o3zf5KQXnLr5Cbf/ehYIRCd/9qpl859rASJhf0eehzJpxz2XP
w113oWiAX1vrgPD0AJKjhm6K31w/5Wt4IiQ4Czz7Se31F6YXYVanSJB8eMxmUivR7lzCT9diO884
EQ5kSOY9xnxQgklD7fqy4+AFW9e+CX8Qbp3V0ylWtMxFi1XtRNPQX2P6OHzaMSBELDH7p2+3jHby
kRKmJmtuzEG6K4GmvGzdVwyioMBtKbWfmbQ1U6d/2iQi6A1EYaaXkjcV7B8XZtKmaN3YmHlDXcYo
1W445Q90RrjsU+GWjCK0gF2keIuxdLOIsLkvyCNkFijbWVYWnpmkt3SwT7EHQ+ZtZv/Fi0yk0Oq+
NFbWBPtRdSBzqWUrkRRYOtShrerZVac+csQuvQ15cHgF3YJVUMVQtBvTWbKskfBvQPrihSGJNqq5
RE5X0pzH3Zc+K/7Eslr3Kh1nvhxNTwNF/L7LSda1Oe/MHVH1N+ja2M4M23sIM2S/nh6LetepNYSt
uvCxvtdwMUjzaDX1oz2Qa9IcgdOK7dWtD0Xivye5LbHxWhX1vph2AmhBh/CYckm4ZWq0Hqm+Awm2
+b/fi8sckKSoaKqjOMi/GLHlEIROCzy7M5eJxIbX4NpuuPDQ5PEaNQCJwvm/t1DbBIXwNBfTbdrP
u4dVSYsYPx51QRRePPKHZ5zpoq47cVJMl9KYeDqco7TSVx+DeptTfFpP0HgiQNJ+JAWwOiifQjmf
/30cFRi/MTErMpCD4Xf2gGjj0EPKVw8YCZ9gPqxtL9X+rzUi2DIPHJ6ZwuGNH2VlmvBFDXlMyzRu
wSIAouvzBZavmiga1xJDhthPhl4jaoa62WxZ5Wr6VxC3hK+JnHDvOnrTSg2qxG6UuzuLpl9F5fwX
p+bJwGUdK8i0WUY9SdrVfp+jiMvOdelbEejeGbmdqP4SzwWur6TE7ZVfl06Fxyq6AUAzVTkvkwDl
QIKk/CcLotPRE0dauZufHgJGWiucsjknUVKRTeU79nPPz9EQgiC1SwsvB6G5B+ozsQLx0BMqr9x6
WLTqgwZ434URgIdfdvWGiCnftDNb8ibwigaqavg1r2mZ7mqaT5Eb7VOb/bV2kbRiRdHxQjswOTAg
sWDUZtC4Wmosg33JAoUGAwTTSuYWzXCfLquWuF3SCvTngmMTnG35rbSwr8T4blm9dSW0XJUvhKZf
aLfmWoMRirBSpRr9lMZc1IKhgiOBtNK7ic8iZY6OCO3HHcRxGl54z+jYrcepBqcFc9XRQUlwguoZ
D8vmZY2KuHfbuxJR31d4ATqKJU+ubbSkbBDMrOfjqI+KPEmqOnCZdfmr7k2bxWBuEjFPaqqRshCB
9ttrPtJrQ5nX//tCGG7eGMg7L19D+gXaA5YYsuGW68XJbRt+jkddGGQYd3GZWH2YissTnHXXuIQ2
ZeKrGNDIjnZ8v5A+o4c8kxRsh7ktbL2M6clpUQcOaa7aeMN1IpZZ5LwfjIDuIvC+HJs5iGHq5nnb
wu+jsAQavPFVMNYf5CUA0uE1IM4bE47OX++QrCHfxFGf2zBdvIcIxan+AMWjzW22u5ObHCr7Wyz0
oKgDJNi6GZ3fiwKqVy/O7g4vTFBAGDCClkB3oGjtcCuPFcM2HzjzKL4IBOYoKHlporsahCLQUogd
BVJXeKkTghMpitXVDxijOHoEdK1N32s0igDhHmogKikmOXQq7TOwCxGFdDmWzrP5UeRcOyg71L49
q13yoi7DAKR9GXBRIrOtRTs/rjPDua2qIPJHSzhdO8ncoifF5lbQXmqzIpl7IUboADq8iguShfm9
ivV3ShPgUClHwfGiRnaw+4nzKhlOdxtyQ/oF+mnQszWpAPmutjcwyY8Z151kPf5ae9PXfENNEJS0
ByVXm2CxDJmyPnD4RS5j/JD3AP50exruKlg1Sq/ozDhzhsjMUquIECV+hExPQqmSh9UvKzdbg0cr
dLCq+Nt4NFBXreRFjrKobnbDBp9hi9r7K7gOcUMu2FLpJj3y7ZoAYL3J3/TwERMgTseuKvrV0Kpb
qAFcpY5wQkeCDMt16jBCQmh/6wA3Z2RnslCKB46MmPkjNlPVbHD0xrf0fFnPUyTCXjAYuYePhMrP
gcpHzhbP8h3H43Z5L2A4+IBLJHxytG2+z9naPGNW/XIuJZVRIOqQtK8/DMDHXyD8DMn3xDrvcifr
1JXXAo6Bsasvkb+jQjBmUHLCC/EQlseXHLwtCyFSbL+cDnt/I2GIGEThr1danEsWNfunLfh7CkAf
Eo6+4qZDIDtI0pLpAu5R5MdEU2+LSJc55tE12cJkYtxaIsc0TQ0Od8Cy4+S9y/JGUo9IzlFKQh/8
G2antA+axcSWSKmeuBpCLUMyp2WoRPxZRaBFUyZZS3eiGO2SMp6p4BP8cGSsglwSEqWEXHhaD8bo
EDI8tT+Q4CfqlbOliqvw2vsjMKbgBwy0NDZLX5ZcOs1ADgZBNb1DF3jZmDX9+yF6clkVffTUmw/t
Jh4ztSfK1eDv2USA6+RZAinOzfB+GOVggGjWoKdCdX09exjFvO9KksN0o+7J/iJOkRmy2MNVwWaT
r4jKpYAZVuAaASYCrZeYP2HqywTmn4kvVbNcD7nWxdlYLh5H1TcF87cFwXDIiEyEDatLHqXG+57w
bSdUwFebUUpfIj3ZiToo3sHX0M+rC5fPHrkw3dm3GV3UNF1F9s5glTpOg+WjQtI9lc/oNplfL7Cd
kkALVwsdjohWah3fkLktMUWZSrMsl7m6Oo/J/5tPhWajYlxJF16S3ZfnMLnf139Y65UuYaUGQWeY
hYsp9D/hGNK5dkJkFZqWhgPPc4qiLydeT5GbhNR5ZXcpniX3WFf5Gv0IJNRKS7/c7p6c/lyANISr
2wRp0weAtiFmO80JYI7kU0mHuOjtf3ZY34LIJ5k4oAeJg2lF9QPIUgjKQIuJUNcCdedEWxwV4UUx
gR4TufBh2g/ub7R6wLHkPqS18dbFuYg3m8G5I4B90urvg5gSGEfF9f+pxqn9Hs/IxYCGVL7JiC0F
ssIjbplUvVUdMq7GRM79j2e70yZkNW2BZvgQUUNC8FQ99Zlx4aYQ6994+0Uwgtz7KNTvUJ1dZt8b
J+5baMNxjciUJ9WMz478hrRiq7v56jJ6HtniYdJ4cJHLzuHd4ZWhaWMy/7BUK7pd3Y/RnAddjj7N
o4NXz7f1u347CQR8pcy2TAdonxqqragmVNjZ3hmBcMfMEoSAySkbpn1ncKK3nQm91PlQI8u3MiVi
imgzx3sYPRNJLh1iRGW3LwxptKDx90ZlaZcaqxK1JSW5hkGAWtStqpLzGOrcNih53bRz8K7wB9S1
6Dn3NWt/rJHmb5g4s58y4SXPep9czTYFPWUqiPHlEFL25n7plZZDv6KqplWZz6vIcBVAvz0+8/VO
kk7pOckfsa0Aa4jIsE2o4qP6l9Ro6U01LzPqaDIc27uk9527W2Ugs9g5ZEOjKgLllgW1d2sSJCHM
DVPkDAxuylQWoJL5oiTbZf0eevyHIhStUtctAbY/bBB3a+EgkkhbjdUmquQ9UDqns2qJ6kxP39ya
uh93D3TObxankBOGpf4CoXbhCJgQLtx9v/BnF5PUtfCZiTi4eDCgjwjMiPvl7nmADeJuTnj+fFt4
G8Gc4Af3uzTPFx5YdQ8a4EsUbUCUN6/tLDktCA6QIFm4ifnkI6AECJ6sfDDLufbZTiz8dL99xfTO
KAifdfLPDx/pxVT6WBZUgHVofWitdwJA4Bk6S/at64tsDOdq57cE+iigUhoCf2mUMVg+y6cOMA/s
UqutO6JgGDJL65zSyhUqNzUC0glqVPJZOcb/SU7sCzLUXB3q0QrARV3xELQjfu24g8/SyQqahuc9
bX0GHIOJ6+ut3EV8/8JvhwJDmEZY9Cg77UK2ueo5bf2l6SOJv9YkzHQOjp/2HSbAYdjUul4HxGzD
UiTY8VNGgTCxuuiykaIW3d+6pSLAeoiXVrwJY99H7WnSjbfXAuQbDm3k0NfOViqLi/JwkRdlb8c2
tu1ZDYzVTDqpBB+JWCh2fqQTymhr6+RDqIWUfGOJ+Talks4d5dNObvhJ0EYaklKc6rVuk7ZGJZb9
XBuNWLnkxftcJoiWh5sXLa8aOtze/JrIinH0+dOw3XQ1wKIdGZjHDHRDUGcC9X3CKWeIDobEMaYf
bGotlemdUHbLfdQGefDMoh3d8OR05Yz/yB5rQBylK8kdtmZ38/+y/w4WqKxgOe5JpSqSeJYqmOEW
fXNZAYP50DZAPt1lyaSWBxooOFJs/f51meUun7qWO4iE3SWgsA5w9tUe7+JtT7jnEIEf2YYdu5P4
IjmZ0BcKZ9flz5/+NG8eUuWdoOpVWUdA5SPaH6rO3Au3S6GKD0S7lBw6LLwf7t+JBwex7YuvVpxk
CPJCrVXubWQkmWyaD2rxWMtHw7047U48wGKaMxEANI6FXA8ivdBhp7xeFeTWJA9seK2kh5rSFKaF
arvl7sLbe4eb8M9aYGy57NtEY1BMec9qOlv6erfmgXgKsGlUi28uVKbJxjHbGgwDTJm4ob21urqp
TNDREsIgU0DgAezIh7+HJSDOciEh8cQG/3U/5Aky9xkR01CToP7QHjTEIN8g00fL+O54IKg8wxrX
MuMtiXUwXzZ8HJJhJXHzl2SneSBYwQ9cmm+xtDAtTbVc6XpJrKE3pHJbueUUDNIlLEocpqH95X1r
rUJmHYGPKb0M/ZOzPxCbNwxYanrXzJh2IvtUV24qRmTTnHJQuqwiMjxBQQKJCSvNzIr0PV9HtYBr
pQYO320bh0yBEA2aVMB52zZguy4ywi01AbbCxetMNp3L/eriKhJOudy98jr5ikzjUHI5ank8xa4Q
6HkJvVSFLdsDfGRt3oMQiL0dnZAbNTfGT1ON1kmQnLM6lRz9YUZzvdEq9vTFV00rh9OVJ7PMg/sr
8x/nNGEUo4YEuLt5NDfGaf2XaYqPX63zvKb+mknd5xwvNE6MH091g0AtewqIo0Lm5ZNV2inYqHkd
dPiHDsbBJSfZi6mhuZpoTEKuyMc9HRn1Ad9vnkhB0L0BKUT2EjpFwTJJAqVeTF+yt5TgVOi50FdG
fGca+OLyDiMVZk5VTFW3MtjgA9LpjHgzPBctTA2kHm+fzAEvshAYvDykMh4yVaN0keVy08sG7A+W
N2tG/EufjDhJ1yI2R1DQ2SWaa304YhNzj+rm7RERsPlR/8I8HWtZkbFJCZ8oYDzuMfMTnkh+q5i/
wa9GpKl6xT1c069RLFgPvqtJSgvEJEuRiDQf2+6NRH1S51U5SDJIM9lZMRVblXwXF8H8i+TJp++W
Llo0TqgJIoPPtJ9rvfqPoNSYfnmR7bLweqDtLGd9ZBVCNg7dRf8kjNbjZ/6tbiO13fBCPSOB1juF
k1BssZPw5KmH/M9qVFgW1l05SE06pcALKVNQTZssVZCh/LlxyFmoNIMAKil9yfbvCxipIdTpVmlN
749JBBpjvqPgbpAroOVyf49fqI72QRlSMnZ8iZ2Ks79Bz5P0roMmOhVRKHJ2modWM27hoB8C8KOs
kER2YA+bMQdE4Cp6ONY+ZbCMPuRYLkJiPqCKTniI/xnaVgbpI90iJLpreJuhjkaQ/yt7QqAE7skA
AS864FJfj5Hu5RYrP90ryZiRixHdXx0eHY7BzHsIS+4WC/myHijtHLEiZN8CRvJXa0GFiTZTAPaZ
auuuu8wR5r4rF1T98JV2i2bFXIAG3DECYkUnD/+yHDbOzRK1//WSmi3t+E5z4ef3Zjz5YnRWehD7
aCkedgENdyS4Q0KX2Ndik96Nkh/z5R/b+zvvBej+Zp5z7527GYwDTAO2T1OUpErjxGtSJHSk2J+U
8CcpwxMz1qhZuI2v5DgwQ3RMgf8g0kxD2T6BPWHthVqQmFODBFaL4NqlnebZbvaIr+SABLXTx1b5
tS1x29PL26ol8s1Dm3GDOqxwsIz9oeoCZpFqMl3WlJC8SWBJWm/SP6Ylgrn+YYu6euuUa0byCEyp
lXECyec5MSHnr+yz7Q9Udq78izOD8n1iqJjs4EB2J57fGCZ0BPhcZjjZkcf752d6AndB741pkxtb
QZRmnZQhoWNTIcfjESUxjyQQw/s86gC/ibd2QqRjiVZtAs6aQjPYV4lJpEtl05fdOkeu9ZeWWTCV
qxlH8zKLydL2F642F3StfEUkyBRdA1GSYn/BcdeKipOC/qCx/K1dv8xHaQna4f0P31wgjzGeDB4r
zesTlxyQBlW9Q1ckOKdvCzDqbRXS56b7HwERvtq99EQEtF0gxih4++mhtNJgWb/8Z1YuAItk03xW
u80RxdbcI94LqXioOwt2HLQ05wLh0NUSarGgkrSwj1RM526TjPjKFvGNfictoeJwhSEidZIWqLRM
FdD7+mbGPeBpkAc+iUvNVZC33T2P1hKUUkPbt11Y2RmFjqAzFOaF7R7y8tC8Tm7MtMOS+F71C/EA
LuEERjSUNGVQ7oxveFSJWojAH2nAKrWT+oaltOaKny/qChMsh3Lmoav6KBIyTlaJTMDaFnRBRqe2
iHgfmS3DkQU5FyK6Uk0GRNeJo9yXdb4LkDXizMBt0jniao8/XigYQUrM/xCHfIbGzWs7/AKDnIN5
+E/TD6hyzc2RccMU/+YK8waPdKq8+9oFe9yIqaFcuor/huXK61U3njDzwfY4+ty8PE/wt8R/1Dfj
O4PwkxRKtcFRTVpQpGhlnlq+u3kHxl8jHUstdFNXPKK5yXNAIXpx5nnfXUcUfzy2Y5gb+ULyGVlL
GxtfP7tHM6DABJZXAq7c7iu5pdvodX8Jo3cvhwUq/roV4WK/qV5DZaoo3VvRBIKt30sprXB27Qg9
tjE2VBinrAxrph4UEEc9UhkkJjCABDbAL5ZN08lB/LUH/yl+1y6XsL7R6eJiaemcFfe8AJke5Nrr
nAqkU5dwxAnkGd5sfM24HpAlMIa0PejlSSts8l3tToD/FQnmf9PBZQ5jQpXQRkz1wXb0RjRZfS9K
91lZKU50GzHjTX0KPJ2B8R1fpLB3ysHj224/eJU0bXRnbIKhI+rR6teJZ0h75Mh0zeHBAvqXYFBb
bDMKlogCwwt00k137SYvYA0ZhS3dGBvfjnfr95DcDcZaL3vXXAa9HEWsoQdH1l9PjmI6xstt/l1C
mK4K6Kd+4LqhVsJbYEDQj72fSPTQFpasHuG4YrAdCwMK+v9VgGtQC7VdxF2+rYPBGHZLK2ywEyAX
9FOEx9AodNNGUWe0VfxrEF7rg10pGskog7JG7qmHuNPd+c3+hOkLCGPQ0kgYSaesytnA947w2oPX
ZdBZ30JGkDhf7z2XO2pDdBJ3L963SRfpLIJ6sjR7AoUur2z0fwJ8MUraqyYRjEHEbif4ykX9hz/F
4d9ONA5N8jO9aczIJ1B52gtkKdC9qnCct0SGeHthoZByyHmp6lHm3lY19dwjhEs5ur1ESu7ENqyp
7uxP2LHVXO7ypefnT8QBgWQOyoCxFdUBqM60axhkGVRd1sR84zSGcHzTlXBL9wIxiJmbDTcQ10In
+cdfWZjo6dNWokRKzXZOj7YY6aqdkmwTDYD6y3GLngNRK4BuYpXxqmRbV/l3ywQA2AVR+vdPDBBI
aZh7XWJoxPGPIn/l8gNaNHAYQR3jxIo+tljZ5lJZ94QmJ0VW1OKozqAfOcnr01CUWoMbPOiHOkUV
G5V5ZZtz93x4qak0B4iKb1+61tuItmlL0m5o3EGrxws1rsaI6aQ89DZGKR453FXwK1dRR/MKCY3J
WS8wLv0s6DS8fbS1jEeehoCVPA4WbzlDI1cKJzC+jIVysyuQCqpE3yhwDdWiyj0AB8VRAJV6hjWA
gJVJE4wkTv3FMDfxSbAjWyML+vLK9dLLT+B8W6aVN42AmOBscq9z+bVkmeZQm9YN9p5tGQsOUFWp
+Na3WUMHCO9zaE0YdS0DY04vnY3IdypVMTfOSu6pFll6gn+yENDWPawIdaAn/onahSA/qTaJk8HI
kSXnEcGww+Omv1KeM5VvJvaH0gXy92SFkEO+lvmct4IgWtS4+gY8w9pyiynZjGFNyAkBpmL98fRw
3SqAsA8/AUTiSirKyHbHPvt2nzgdhD3g3XAf+0QwOmACQX1xu14CbP71UCiwabF6dUo2FtoA3lrz
ffSlijyATqU+AcnuU61X0sIuO9VxlmLc6d89rgSR6AJW138kNdYRWjRd7VrX8QA339Hx2szicq5G
namDg9h1fWHN0IkYGE2b9oAXcLTXH9oLTCx+ZBMq0iuAH2ZhpaK0IvQhmkTMx7Ql8IIpN5FAMrlE
qGBIsWFOIbaIUQUwCPPS2EzQP9FDb8o6yQXrw7uCt9ONz6GiTK8Sl/Zlkqdh0A43iv921hMTqqDL
zf1bBgq8P/rF2D8KHEwztdqcbYMBxiLcnBTEqWV865+C6ajo3XIMm8L1NQaYOtmwGT9e48h73W6N
S4VKY/oe4WW4zpqbLRgUK0hDyex4MIN+ZHDHbl1NqTyrVGagbYMeg4PkiQ8HYEZJHl0mYx/9rdfJ
xq81lV9z/dbD6CXRx4dcXD3tFjfrZFD2StkSuFfLGq3hRxLO+if1xJUXfCXLAb8XjS+1pE1qZB24
YROXgE73EBte0E/mB2DxeZNFAky9YYwxmi2cQ0wc8T+I5pgTs+7eOGhhqLlguDPANNlloM85V+Qz
e5pwEV8vEOlM57ge2A3aCohNv6xW+Ex9x9fsLuVF+7N4DqOR/d4j/qH1y00ezA7jT+0nJXini2jz
V2YcFRpzubN3JhO3zoJ+RfzAS0j5Zpk013p0T531zUo+Yhcn3KdQKbQpkV4MB3u7Ka3yV7tdCYzV
vU99MFgNwcwI2+5GrAI3DF9lTvzv05ZcJ7FSKjwM0rn8joMCBhYD8halYXL3jL2X4jSAxTiR3fxY
QUpm6099ZDnGpqNFqDZPkQ5XQgicK421elGIovzp8sFYELXRDNAPwh8FhZOy57GZUYxXDpzkEmvM
cBiei9LiSwbdKIfpjrL+K0gq7Muo+jhHVi6lEV6zP4jna8fgWO/N8qXHooAhYtvvLHszHChvfOuX
5lmy5uzRQEA7XvJdTaqOl7ipuZkNW7C56uQUDis7V3RbqHJ8gIobLoWlZe8QxwYHTgNSpijIuI6j
g97OnNSaV4JmwZyg0UgdkQVdgZommJ53UHLnriakahIEXGA+EXvFTVc+o6+pAsvqJiUYAOtAlVUg
wTsjR8vEXsKGJlL96O2YTURQeAuCenUeO9lwT3wWwEKLPjcG5XjaFgGkNidrfqWql3keJovOxDSP
k9ZK/PctvJHK5+SWpchv1jMJQA8ELILwsa2Stif6KtnBkwu8sTUZe0dJY7cMo58MXWg65YzLPXG0
Pg3dbFB1mOc+vYQTcrbKL27B6FbFc+sn8dg7VdD8HucrcqmEgMyk0o2hVNXcnSp3Bd9AKjqEgPW5
++FHtv+Q7QDg9mXMNl+kg5FvrUD8Npa5byE9SphhnTxxAsFYQe5WW5RiBTa9AbDmU6BygEeux9lZ
Vw00fo3EC6DZbFFoLkWhgpVE9MsPvOOgwZjZjSXL7oaDFb0eSwIUmwibxhPKjTOeG/yZJBjVeNoV
x5rqfOCbwbGMV55rsiOVpb0kkFpeJ/D6p0BovvIIUpj6KBCZ0Aj0UhK1eEXuRtxKb7Iw8bsgnfJX
bc4MeIa7i6Jy8/oPll8kyqRA6m9+BANp/0YzmIURKI/bNrpCs4wGd2e88vvQtmU3N0i4yIknHAIh
r22SXXIVXXzxLCjhntXDXCQn589egDTVUsue5FMZpga/NrztX0bpuVQTv14I4sK7zFsEgIKFmDYE
q9tCNMFadeCxrvCeiHYupZetkhYsvnSfRKlETkUXLSTmwTpnFFlFevToNOaPfzdixJG1wuZr9gG3
e8ws6DQcl3CK6rmH9Zt+OB7nRIaoUcwNFRieQsqudUism6E9Zg/hUMPLgCTJy5I+7i+41TXIKwRL
m+uESeqm+bC/70ETgz0DnpdcqXcvvl9UJIooVXmb3RvV/N4Q2Y7CHiYeszoVhsbjOmIzqhT0Rn8G
JCh4y66JUHoaJ91qUvFa8U23yQg4LoLnzHRJiPCyRsEdj5WfB5a6inRkjnYAYgL1N8bVZaQWaenj
g2ERg9AwZBU6XYpuhw+dRKRFnWPFdpir5K/KOpPyoWqQo+s7TUMlqOEvRlNX5CLRivibZGjp832B
6N8bxWL/53LLEUNk/nkup+D05sDCSE7pXPF06yz9nIzE0XXDXXNO+yvFnGuiFIapjb209iqcFY9z
IO4rpkY+NJesJpCaLStflc5MeXyfvwZhfATY2rrZiXZefzOL5zhQUrXOfzGaBm7Pp7xRFXDrgNyK
vYoyz+duxsKfxCxsLgS9063PpTZa7PqDKx1z0b8UxTgHJ4Kgm0Z3QTZdC/b3jhQs4PzJnBSDUhFr
zcOcKoElfLt7sEcXUPOO+NIBksfrvtXq8qelnULQ9Oln0QCnKpMop5ZxuWXLE5nN5rsCjrcQ8SP+
8FhaGkuVVvBtynceZiKNto8o2Uf85HcNaywBnQFpfb2vlkezuRVaagkoFM7ErzwneUAlY49f4Y+J
9lhVAjITaOr88bOTfryf9xaBxX4JMeZul10pwz4PGKxu8lyZiJQvE/lRIy5OTyiVZzTl0dw8RJJF
POuHf68SxHPMi55+us45fupH7V6nbZM6YSIc5W3pzAKfiN+/XxRzEYIDj6YPEDQtN4qEXYik/M6m
EtS8Obw0DqFb/UIXUlvCpuCy9sY44f68LDlOZZkOUg4a5dl2SbwoDGO6aRcHdkCxbCoBN1MZXRNh
uhxJZME9ibGF3BfL/k05Xk2rV223XadGqX0Ze0+0NYbGfWUIMkbyoJiwwW5+TNmskHfNgT5AoP1P
ZgGnI9bIzklF2Ors/AWUaHvaNZojqW/P4Jun5yvc4++ya69TwK4YsJGuFtxfoKlkL8o/GqkSG+qa
Jfc1iXF4bSu2iVFA9JcV1mw4TsYDHDQxDyOXydx+XV9sXRldOnmKCEHd10jGfgitEF21Vw2/2c6s
v7ppqQ09AtLUEtWIaOEGnybJKgLgZGFF4eTefw+iPdEYEq7rT6KnnLpiLylofzigRLyiRzrsCdrr
lT7HSL5ZuLg4SHbYYqs4V4eA7KCJ7M1gx1q0ZqhEkyK78oP5BLYLsH+R7esLnUeA/dqQBs+3wkvi
no6QUoSw57n/OKgpWj5Zj8Y5+vmgtMcD7wCn7pVrsfVbpkVVbgsuaNxQeebEs4NorgZvR5XxmF7I
Qfb8vKXd/Mq0XWXl8m1eKCh12xO/jfQ8iIbcWu6Qe4gDIzZ2ww6l6n9GizgIobp2qkD/lzLvlNsL
KQ3Y4O6w+IM0XD8Gp8LkktjLNvV69DTeHntlANNiMvH3IXuDVbrQmBioUxDbrbMRQ5df2pPNl81m
jFhRUBOQ+ovJnSvGdIx5xMQk5gnkNLLehqsus8kFTuh0n9wK4h+YlERMD2WbzhNHbPE5dsBUv2Dd
6VHtEaGv+iQMEdp6o6TD/0E6g0GnJCjS8ouYNwaTTqEjy0t5R7DbGrxofyAi1GLiKDvkqdERBxIx
3jz4Nfq8cylUmyqldlFdC7IN4IwdAxaWP4/3QevE2zqyvw+DAiMlE8bnCZAE8QBDSDH+ZZn3MjVY
RB9tF5fX9CmD/9WCoRQvP6+U8emOD/Csvrl7mY3VsMXdTs3Up/XdAtVleYo9CC9Tc4YJhQj6YbZv
qVVXB9Ijo0npIsYsQXkx9Nlbpf6SZP6SaXCLtVck235MKlodAchgJRzr1AFLpJVtFywaokreLji1
nj+14UE+IAR2PZgCRluRQoUZu8dI8Ln+eu2vToyAN4PWt9cClImq5aUbFuV27kLU0uuMNPBSF8a2
xBRIZytC1Dgig7LAAkHWcUl7wBxpXU+57zPETaTwnepVTvvZIbqeyvsRW8YWqwbYauFKa2X859eZ
eAR2kZDWieQEsOFDbQRq7AX154lxMQ3tc61ZMNqIFi5ldXIwl3l+uDcCRjQK+sKxM2p7k7sB2Icy
XO9KGMSod77e6prGCvdrswBY27jGvLmvktdAMCieQ+2rCCIGFX/CNonD1HBTKoVuYGbTBl9tDDQR
oWhxafdcdCnhfHfRf79dh8qLrCm3YkRsh1k5C6BWpwC7nKZDIN5gr8h7q7JyOokUJrLL6fHRJf+R
C2klEq7cwPhGTv4Vn7Pd5qX4o/UG/2B84UPwytcsW3xzw9exZgZA/eAsSmq8IbyOeXQySWYsxMJP
eqykaK02s0M7wG/jyP1WBJ/rTozaxd2M+FrL9Yf35D4VjYcReu0icKf6XTQI4QPYfQR+ZII+e5sj
WJV1v4LbL35Up3vmJlFMtIjSANDh41EahiSfgKS55LcHDs2v5c1nYdWnWWqyC08rdJRji3B5pn79
8KLe4HXUXK9rxhZ90uSVW6kblyPqFWa5kXTFx7JIi2O5MUyvedOuNIaabW72OIeYbtzAu21/125o
BtYNtrSIS5Rsp9MFQVzAn+8rFSvMe2SVrX3Su4jOPAyhkvqkekTXvRLd0phHXfb2TNJ8JOqiTnxG
cIMi6WB+bgC9bHvqJ4htxYTbEYgYvrvR+z4CLbe37L3nagOcBNQOnkxcLcNwjgTQ7TLprUtiyYQ+
1D7Tz80IqfrZrYG6baztAe3FNdcZ0OQnxwshyF9nxOAAwDAQXVSx48TiAIQS33zkCGzFYNXWKwe1
CUBwOsoa6+O76eNJ4tY5Q78PPe3dkGR21n1whZ74Ehld+VfHAWSFKenjgdqCpUVwptw21fhH6IJw
8Zn4/SYEHxqzzKz2y+/aHzCrOgDbkaKoJJRMZFGRJim869ZCrIhrzbBr+4f+CGLYLExa9lt4Ogjq
l1Y0OjaRLHt90NF3r3QS9cT/+WcRURVotCku2g1loYVrLjsB3RHTWH6GpZcd7DuBhruZwaQ4vkyw
oPHIj9WgrxOn+7EvRRFyZZjF/IXCK1zYN8pFc1GmWIhwYSGEbtFQGzRaVRMpPG4y4c2AXjI1JcB9
4VmbIJJLqUlBqvmNJJKHU0Uln4gTv/zBnt/KzK9ysGsbXVHj5oJPDQuVwcUnvKMGxnh9Yjsyqjpu
Fyv1vT3rILF8f/40J4v5eWcxjXlwd6hwl4UiUJLDA6rgO3QqAjGQue/OdSNccwdqTZqfOUyEhJhw
wu+t/M/LKUl+vXGC8vDukrfwk4iX9nyKI6k1dJJXGMiaCpKsiZLitw3zuNUvow6NH1DUEtV49bNR
FEAuixVVhxnS11FYdjgRzAnt+I4N3wCjngHdTZaqmwAkL4Nz9n7ZVd+IeAbw+AUw1Q77KHhsymhp
fynLYQ3oVEqkD4LndH1qCAH9hcfElUjRemoiN64fc9wqvUxDWPREB/eUbg6ax7Y4qfVhXsWrfDbM
YbDGOqWULI5k4WRlV12QZS3EOwrd+ATUI2ay5PJA8geqyj+aOvs8+DVZnb/vvkq3kAA/p9zQSMa9
5QQp+A6cROqJdO5QTzvjUq9+7tIi+UsbYME7CjcAL0pc5KL79B8joMOZdAyAPQZxBIMSrcowG7HD
rmyNbIba3bq9wWcqaDP/GVtRuCPddSdr6seMgGqZk93J3ILno6z+3G8BGDCoug+jX7TXVXKU/6u4
/X1mGbWp+JVQ3g0KmmBsw8zTwAzAzjZk9lfv3CY96869XTMv9usaNM51ZdSSCibuhHnkRiOn3QGM
l2Y80uaav2QR4XqKUjfYDLN0X8zTPc/4vq3l6BWLHy7175gpt2NtC9t0nzEl8E0FpiXzf9m9LVt2
c8Lf7xr72pT4egODCkcqzQcMGtBheo/3moqrntxEws2ejLFCcwxe0f25wXF2xvqFbFjYTAbQW69L
Bg+S1dTCxN2iQAg3Rr36ZV0yT2A7vj4I8HpER95VR2XX7b3QMGL1N2RxEWdZlcntyHSfTeEjj5T6
7vtCT1KxLBbPpSLEoAbak/0MhXB+y98h1lyejrDdDYOEzxjNXu2VN/MzPXxNiXSCIbeVkC47tqNd
dsFCtAbx8BVVmBDIsIIzk9tSF45jGSnCTUg6m2V5zM7VouqaOHN75wCakz/vbrt6mxD3nsgVQTCa
tBa97fchzDNPih7nmOZ2WhrYbvKpHcpi+PQwtlU3hE9oy6bjmCu8nFYbo7J925eHCBzNo+znu1px
lyE2dJTTRWR2WJDOpBQEYiudLl/Dbkg91vI+zwVBVq0t9G89aWdk6r4cqtAq3fTaoz1O1u0c3BA6
00HitSzHAF/XrJTU4mdIxU2O59me+qnmF6W9+Jmf89rXVVU4l8N5La8oNXYn+bIGcEgzDZtHBxcg
dYKc+gJGJ+i8OIS71WfFGAoLLz0kjc1falVzvHN2QTocmoLV996TUE7wBCj0YBWQgl3QzvhjmMZC
L9pagEH2xb7nFXKYaVhbmd0kwCc+fXI0WPirw5HrZpPzVgmlURjuBvkowm5U6+I9h3CFBisjZRL/
xyQeHaI4ewAOzqY9Kc0LOAJ4BnTB4PXwv2FPpsSdktUXhE0jt5lnOhewIqGLoFFf2hvyeo4dywPI
Z1Huao0k0pxk5voeYsd9gQKNCM092DY9FuEJdMR0JYNClRGH4aId5Cewhgg13Nys8KixYBuQ9b4f
kslgWLwD3fG9bC3hyeC00CUU0hiyIkuaN+04Ba33XAxAyRyvExjlItFYHXOTh6P2UqnueCtEse1B
oTfZyJf+TBxKJqjmM3HgqyShrKEAdVICR0Uet3MDnkMAxBvn//vbN2w/Pnbf0o+ELM28m6em7WVa
rZrZc1HgHpG4RgP8fh5Ngp2VHpa6K5A6iFiUCWNLk9OHV/KDLq1lI8iHqIy2mpbKx0dThzAn2W73
+KdGTFJmmYv9h1vSMx1JGqOmPpUJjOQPyTofAyfjrxV4gJzhbujxozvT+MSBqCDBqlkY9VHD+Ty/
NW8YPsuBIa8zcJr0S5dpesk95O0JpMVKvvl2bYffsjTtiFH6BHyl0iEGpZBFDpAy+I7e8F2wC5+E
nnVrNveo0b+tc/RWbL8Yf1f+enZxmf0gr92LQ3/gGXpleOH6WW3mgibPNrVzwpIuXxe0jJHgGnVp
XD9SxJWnhAujeJ9CSIMHIzJ0qeBrACmALgmYQgOe193os5RY8W0eGYq979APzRxhl7Q55sFBZvz7
YeD2PwRQRzJ4HbOFQDHAOU9Qnw+9DvAddTNht/k4gA69co25li4+pxN2FHoLSUWGiudHLQUER1lr
5hDYxU9WrcNnoPiM83fTduIgJlwtpDVCNl0pKeg7wxw+jD/47Rg8iQ+tc7ltGI3ec1UI94noVKxm
aJgqgwX/N+MvVkI+AE6VQoizdFEV6yyp6kwtZEBOSPBvqySu0jYylsWAjhOnjYKaMBBEnRblwEbZ
+8n+aig9/JAlZcj8dOZCdIT08KG5iyS6xkiMnSNnbJyv7QBqqFuLuiBXjjZfijWp6keEaAy/Rof8
WqU/ViyK3Lglxiy/SkSmJbsEQR0Coi4c4sfnWq4CHGObZnPRWWFqx+LuSY9KEFOr//B5aplmtcT2
f3h6F9B6+d2l55EUb3J+liwCuzCOfthBydkuxByDiwY+4hy1AE1JInaVTdxNapBelGAtgMgC0lq8
Ly4RZxfN4yhSBY7WBH+w8ZVpvUaBfXGlQFSlBiIN0lYSxd8neh8MfWOKNuU7+UvVz7mVmyGy0f/F
2szu62OsF45d+JpL9xWfqyrBCNb7SCFU6J8D8wnoKDq4wiAOzu4ddp0il/m+EV9obJC0RVhB/qpq
Fj7aRV6kJnEjbImyYhYEj5faWyLS8bBWqQWmLE8PQ07pxV8scafBjOqzqJ7EUhWxt481OKnNEV81
6GuiZw1yEmQlres0mLKTvpobg9xACp1/bWPO6+ayMJ5OOTur+BESId3qVtC0t4cIn1w6ma6jdZjg
WzeThDf18d8Byf8Fek5oIAal3O3q0wnVpSYvzTkWPcEbNZ/Q4yx519r1DxIbiHarRx5WW09IVMPk
G2mzQVzXkJwxBIHpn+pAhUgrwDh7UZ+e+lHRYV3FTI97Cq/sCzSQCzvGWMaRjq1kDjjp2/X5kpLy
87ztrm5Fqpk3kOU2RPXZZcii1JL5OWWysNAuoGb7FKoev8MmLIHHvw0qaUWTAw+uP0t0Lp2wqJW/
FBxHwLHa5lpha8RwxzFqRAaI5vwn5d/ctNNg4zuj5dTjn1jJN/FY0IkqY3Q0Dir2mqJ2aUyxhr7T
8QEDk9zvU84O1S484f+Ap2ZGojfIF11ZQfYr48fPwzZ0QyMdr21BmPlBr3iquzaNmjI8bQRJ0rrE
8bRnZx8VfB8ywG61nWE685cuZ3uL7CLErsNOR/v7BvPIlvEE4wqSFvo/LjeZHolEVVTYQZNnY+iQ
W6VjUXAQMu9pxTi4Tm+YVTWlEHMTIE4vDcghEZiKHMt7kh3FUyL/A8DJ1NoJfG8cKQbdz+YA5ydH
19cBkl3wXqBEfdTVOT/EdOqGbLwMtyx+QNzc9MFfhsxOjOfoZ48C73EKvaqh/ESSrn+qIJfmf1vL
T4O7rcHM0JoeV6lVfldC15bBCNtZ4CqH2tr04qE7tHiQaJFEqyKVixrwyUb9sciE70N/eFH94UIP
g6A4Ed2UjOsaC46OT7BizEQvoBCqkM6rNgKSCpna5ZMs2gt2AE+YkSQuIijtBBYkwJH1QnRjStWX
klKK+VO28Ei9/FGLXQcxqrazxpdC+2u0fHC0hoVMofLIFebHqAKH/Tgqj0IVJdLZwRzrwKBFPluT
iZtWGUHpldsaR/1ElabXKRK0jmpoJv3TB8kFbbkLwFEugPMPP/lsOFTZBIOr8Moy2n0fYckzLqtv
qK/7KtGvk4XEbTfjp5t8vKmODD9WtRDK2CWsjINa6r/yuzHnUgtAECXdMgoR9y7PMoDuAHHVgZpw
TJySowMoehn2OyZDoV13yGa4uf2J6iymKb5KZ4hdNgjyA7LWTkZU8zbpPOQOBflGH6hpH/KNVwLx
Aij0sIv6bz4+8sRudMTN/0LriCw9s4iFmMge/GbzBrUwxNOpJ3SrTiEmHrELM3VVx86BPRSXC9uJ
d1nRwOxWaip2bAfhIPQ0ab8RvhXjNUBRfpNfuAO4CinkMGu1VoxuklDONsGu7OkKJPzhQ/pNV2qy
JYRQXL+UBXROgZeFApl2guoXQsAqHARn8DXfVW9LuveF+i/JYsFocD/XRnHe5SWnDK97UqdOqdV1
NPY/9b7xvJlV+i2wMsSoWWxovXvyrXW5QyB+YRGSAgGkuSWnXHkmo06zlRXGtnldEuGLq9L5bBLC
mizICaAKaKR7b1I0SyTrW9chP/+/oyHJkGIuOfoK61lFgVjpa/m/+XxyodBenXkRgRFsdg4h0cL5
sKdDWYlS3EQ08gY1ZNtO5QlVOB6N6hlsuuAiE+KhZTJXq7y8/e/3/H5Oa6zJcGgj9mNnjfFHesEs
vnsPmrhjPdj0aIuS3jWp0rh3IS5fW/RmD/JbV6h4MPxpU1pTpB9WBKM8ugA46alJePHAtFmqDxGq
gh6TRqfFP2Z7jNh2HkUUlQD/UKU1LeEoOnsGnYdAKBYlGPJDgFyxZCU2JEH66BSojVidnprOvvZT
PizQJx4h2TY3GQY2v5x1K8yOqcwRNPRMS+kqFQrRqfs2Zo703Zc1lfHtDk8n9ziC8zi/zKXFFZ5t
7WVTS2QZ0MNdbU4IzYKjMv2XvhYaFYl6VM063lbgDuTdjwbj3Ujl78qvp8KIFMCLA451pTaPeDeB
6zjDJauT93JuymQYIgQxdjrcG9dQiu2sI4L2f5rC2rBDlMuvdIb4qxRNkYaxlrq8XTZdEispLv6m
ynfr1zlab3nvlC+6LNDGLi/OFEWdYq/KljZpBorHqEljvbnCBVu+LiGhcEFGURavirA22ahYoHhT
HNp9rzMjqDa1o8IYPHN/AKg8S4IzcEPhiBmG6GNybYgjceHzuWhFXsNge/jqinb52pAxbF6kmFM7
m0FPpr3tcn+xQPtp2nUOx6RW99z71f7rNMvVSbq4D+yM3OcTp9VSk+oMw/22BKmy7iH8u4gyWrRz
lxKWKYGedh8eXfDc3IhiDWepvveXKQwQShHYMZ4M6/qbBn/2mHRBaRnUdGbnNiUHWl0KeCGyFxxw
aQz9C3K2RK8CIqilA0kdpzLKIN1C3F4nEGBRCAsuZoWqRLZ983DhueaDKMBdOOn1bcgCYxA8X9OF
p1UFqAhBxYsnKrFvRKnlhjAWBJgeoFCkqi811GH6g2bFKeYMwrYLKWTcVUpkqq11ged8BIv8ovI3
aOObYBDl+ziDAdURgbBc0l1LHjA5P+jBhYouAweSHaxyR4BGda/QhBbCYEq7HhvVZUF4xiUcc+Qk
KoRm7jkppFvvms10Yrqx0MiPd2lbJNk3A/F/LxaVmftKEOoM5tQcleQn8flcPj+rh/Ls+obpx8Vg
Fw4bUwdLkhtpTDBIR78UqEs52XOVpy4BPJQo2PRF7SzsC36a4CAuzYKA7zmpgK8EdImhvExAZ59m
K3OJaVVZg3SLizixZp2A8DZIOZJdaMoHL6cfTiN0rcIyuzvTEpdfhfklqPWIZR8YMHpNoRwjNCXz
wA+ojVR/SZbgrDJ0rl4guHxci2Lm3K/69vXB91MmOLoe8aLFwRIGn2fz4qnr+HiiAZcHeV16ruRc
qEf2G/jqElGDi+rL2UvPb4MycppGWbNNG2nntozTs4QJ/nLlHodpLJpOXUD24SDlrLcEPQd8Fk0J
MZFGr1tw7z2Oe7rZCsGHMt+xu1gP4cvn4Zd0dWL+gnJTcirTtNlcP3pXa4TcpW92fQJ2lzFpRguX
7TdIq1UgWEVz9reFWvn3pv5VHW9HbpcnNijXvOWyORC9rXC4LQ57iSz+lOvou7o2gvAYvuEEwTaN
fr8yYVH9UPMhDp1wYjn0PpdFp3cfV8JdzYTos8L0O86tP80IJaocch31JcWT/nOIHAYwUYYKukrq
Grsah9XubEshePzmZBOoEKh3nenhASR3cr0/2VvfdZas3ub+8TGaGsd3IH4wphNfYxSF8sjmpVf0
V5hwtw4O6apqeaIPRX3Ijo77nVPrEkIIkWg91BBshyWXSvCg/WXdOdgaWB/Uox+Bah/zc18HFx73
jYZKqOE4XADuXVMxTNSxjfhpojLDcHQc7y1FE4r3IGuP1frgPJ2BfFlN942weXpENgpOo0cQqBkh
hfABHbQGWG68f8n6ylNxcPoyxhq2H+9ISs1J9DMzUJ8JSFnv6cKL8CZMzyM6yBFPS4aVmwBAmmPl
HHCBYUvzVd1qWNf57mrtl7VDCZI3R58uZdaXTjpiSnCpdxzd7UzraYTOjfxE9gqLljdy6DCbeakL
AdKeE5z4X5LiLAI7R+5svhmrG0Ksyc+aTqbmTB5UaGaN0KF/C+RT0IHKVzaBSzjNg3VGcFmGPuHy
IpO3FvoPFlyt43f92bRfaKITBrbuXBq/GZntyzkqtn48lxkUPX3whtVE5to2AENWwJXAZ3LmlhzR
CGi9OXeBetTsktNeR2nGX2vsZzo7vrkP5W3dAikcnPjVYfRuOsyUW9j0okoR3JjiDi42XnnUt5BD
pVBir+L/vy9sxakp5XyVmo+lPKlQJmbvoaiToRWu0iK6x59SYO/m1Kz3uLq6nmxsDJdK8AvEzDd4
9dEreCqP9S6ZYS5ZSWXFpXaRWX+cEMTuLokN2SDWsxdPhtCw0jc/RwDo/gBEYGnx8pseoEDwfR+D
W26HcCwmBnVrHVhcZJHn3MKu2K0FdSfxibeoD5Q16Xzm2nmXwTW/xBY+9I58hJyicw5yjD7rqH0C
0Imvqd0GqKneM0VpOY4B4qnUt/ZSEedfhgvpkfXrLQUraLHie2RbJcBfh1KfTymIBgfDPn/T0nGF
zUPX5uOeFsUGt10OkHkhuWG7ZeIWFJ0mnfICeNx2si/fvyZ/3H54ByMABaQd65/Nl3aDcaPPovKp
5j6iY2QsOB/4n/Ry418ewkyTNb1IjTY9+BXXk0oPyvQo4jFQwngE9rJkfD3g7qUWHsjO8HhVpxGJ
WxRlK71KN1RLbf4DK/GnY+MWC21L6ElEjYw9+8PVkW1fEU3/Yu5bX/StWLK+oQIZTZkOOE9S8OHb
74WN8/5X+HGQiyLtpGMnV0f1ckJ4PxMVCDg/MJwTWE46EyNxl14L53XR3l+BOKheOuEyhEhwr5Gp
Z5xhVzpB+/zBfmgWdM8+w/6AgXEgUAlbfzwao7M4KYAxZCBVdCqdERaf+c++TEN2LP8g8XtTGJHq
7LBgi1WDRCI+4kdrwW5aGv/Kxo0+Ve7YqOvVNNMrbzebRip8XteNVvTp9bg6YO+0x9uPolXmRtlG
PmC7J4fIDoRMQIhyWqGJmhee2KG1AFpKTlqtUC/5xu912mzi1kVaxW0z0/IgSPgSLkTeA59gO/sp
zPlhj4J9kCEjL3aeur+GwzS081wlEjCWQNuK49gyJpiOxaKQBdv48Zfdy/Om0VIreLTxJd+cwT6k
V6y1Lw0ymcYHQYxVA3y9Zqbkp3ElPBXGSpNeRQKpcxf8R0RWVkw7LutBHSar/29BXde/HMXsucRN
IM1ih6xJ1Vz/CfSn7gMQZW8H7zyIhXcgH/xrj0bpMLywo0vVOJNqxzscArD0zvDeEfhAwrdRx9FY
yA5rj4/ARJKPFAjXYTmVp0AtZ9OPn5t7COyJiaC0r8dWUvq9haf6Id954fUPWl6QNtn1ITCJRAHm
ouDNrBLN6dVJz4IGFxBqhCxafbJv/qxqyz8ZJ5HFp5lAxJvS0D40ediykW6ed7bUUrM3ls9bqRDS
JsI0qcFCWWh9djvCasQxAvvxOZHoDRteMCO7hb6DFUwhMj/+9xXPm1HSYAYO4rUp9ea3bHQfed89
ZbWtA93+LrosiHXAaKWaKpWYWQ22tCCU0NRtz3n5uRSLm0cvpferE5hGzcenx9iUPw7zV7PqVyGj
iIKKf/EQBhm1oIEOpRWETROMKNEkuRaULzC692PFEHKx0Xw9YpzN1rlRWToLHu+KY4N3WuTJAuwO
tzv+o6lNOKucGuH8k60UnC0Qq6M/drYB4V3lnPfzZImk32izAconf2+u5qXOSdlT5C775dG1ghTn
AG5CTm1bp6PAIquwBNkibbxr18vEjfhU5sijLvVs4JFarEJ+ieutJloEFjK6KO7F1czFiBI1kliM
a8QGCnF1vsJp10igiHba3MyAAK//yTWaQx+m7m2RosfZyhWfboBe/fYlk0VRI5y8TJG9FIvGTlls
IzJecY5mR3CBapQt2ngjVf3QZI+xj8Uuxn05wNBmANl/cseQM8znnosUykCwV52CmkvlOc4qvUSZ
NxtkALfZzqtH9IHF59BYiM4oOKJ4oKAKpjfHapjsaeaJ0tWkRQD3+7BPBiwV4eKuqmWp5VOuf6uK
QN23kibee1RZ5NUyXH0m60RlJND79FmPFYTxRj3vyfmFMxRSm3fKOL/z1ZFtgt1kYH/lo+sICUnC
VeLLoUW4E6YsxaRS6FJm1JG+xf98/ztbamk62AjQi7gA+zd7YAoaTO4fY18v3XzL0TIPL/2J7ZSV
ZLUzP42h0jZF3kBiIEOV/9h3Uzp83X2kjU+7m4VCRGocF6zv7+JssdzMEAB2Oa+YVFXv6oTOZMF8
9RL7SkwlcMeVmSC/sLksBLTuhNgC+PkWS2X+6KJYwujF6tda87Og4fghPZbEuipUstOXphEBc7Nm
cd7pIT7c5KMv3igkBKl9DhWr6ZeFjosaUh7vmXfH+OPPZ/JgEUjWmCoxoJays75EDtaDRdEPIYvO
FlNYv9R2IGI4MOuw8YtCWm1Wy9IU8GaRgR9HgL9or9YzPW/b1spNwHUrfHWWwt601eIdLpyjnLrA
yYeUHf/NQCr3bj9BOtIXB7LkxZ1BmyXCS1/HHwzEPpCS7FlFD/PT1OyjfJtF0Bg0ymRMp+/ZXJbG
SuqvhNlgPpUIXxH6Wr1heBollfrh++dKn7COalZ39t0SgbGR2Mc2wbW4JLe9xtDhwuShWnlp4NLT
LrwV1xZ0MVAInh4QBNUrJ2idwf96nu/yimmDTT+MkJNv8fYi1RaozGNdWY4XbvM2Fp4Wkx/xgrC5
o5nwyMpeTl3JsLIwcoj5tDM9qAU8bzDDv3CykI+Rt+rcCSXefn2TbUkV7+46mhPKGQYYB+VsyE7u
fFoTt7tbz+NOvMu0VTh2NriY8oGQ4z9n6fsJ85RFodOa99MM/42GEOVHQPfzdt6N7t2K7XTvYd83
kPVg9IevEIGW2w4iQyB9LhtW7ZqiDzbQw1I2PIta8s+9Gad1qpzKQmV+PRptPYa69XJiQ1YEbWsW
YhpHivUShZonrx5Vd0aMCltF09zPAvx5gToJWQxtlq3As6BCS54bd3OPfb9AdKOwRY3aWTUilfm4
xFeZTdDPvC0OvPeXLxMwgeKQtkekwh3PNEfi91dWJi5+nkmBZ1xUHWHbDuV7cFOd9vDxFtofrM25
LSYGdZwgxr4l6it1ocwK4MfNGNMSgcE1UGBTuY6o8P6mMBngBZBzsL0cn1crSCB1kXiPYz/s4mZV
8vlt3hrTzW3Kiemn5HE1pZF0NUk8XLVCE12obSPIOdndmGnPhD6KJemspVrlIvjw0DPowABFlg9r
X2vmd5mnAXR6td9vc7Qx+wgxYrwlaJmPOFrsfKMlk6L/mY2Oo2qZz6EsPg7RPXJNgiZBPW7wvex2
5AgkLeqxz/7KZN4VTnkppSe0MBATY5HHINUEl7NGb54a53eC6+Nca8bMbk9pSRgwQ+8lX298UQra
OeFK4f908XmSCKBsep74pFYG1hCPxdVp4E5nbTHzb9UEhEeUxCplgMiDxp2b9VVnzrH7uRMxYAC2
itJWYgHhQyyD7ktMaO6/jA3VHFmJPxmfhNlmeVMVVRpdGmkT2Q1ilPWhKAXFpv3pdei2mUW01nkP
ge/ITPMoOgC+71l72aLiBIa5Q6Ts7dt4gvi0RhJlANe5RQ0+ItgdQ9cwwz4x6CffIZr7X87MS0O8
LbeO5T2KhOAJaoDhacKyISWyXvLaEmy22ix/hBhIp0naetbHraxDRf2W8LYjedXAi7Iv4qsmHrfB
h1Yi/8l/RnNORWoez2vou9wJsR16BLvM59VX/050DJjYHMwdRBXNhHgJo6FGWwVdImHBfHgDOniA
MiAtByOcCnQkI72oYN79HbcHTLRhowDqUWgS9OdgtnOu7s0Hhc5MXwhGo7cX94AbB+pR+3+DuJv5
ncjQtO9c/wxL/zzE0+mZsSSZpvPjMtNMWXlAswZAzEcTIXgizwXeP+47oL93jIIAOvPjGSnY5eJe
E6QB8Rt0Maydj0X6d92+Mflg3aFNtCdSLP5jKC1cGJS+lOTUpWUqpVNNzAFyLHXzKyRKF8i6Zr8X
vLCK8qATefrR6x/QV3nTgG9Qzrt2czr/7fMrnE5zqrefG0mcFRbeRWXVBjJoHfilShS04kcJ9yhW
3tnrSql5NbvIWdZ4wy/D4i6v2gGF7pecpSNZR2qsod04Ebjjm+oWMRtTnYOp7YKhSzND28WTz0Qc
pbD5axpNrV1FA+18nGw0qgl3GZ8sdwjoZroGTiClu1qWYpwuifNo0+1Wfbvm95euyGPrO74CmMjk
PYddlUUEHV7flVp1ZcNjJYbLhpsrSxV8oLKyTnq49mCb+JTQcMfuYVI+p7oCeE6RF3Tbk67+GEEb
uD60IHsYggkbO1vPTIJ5RX0UJBjeJ5nIo9IrNU0pLJvS35ijiawedc/G8Kg02n00+ydgKj3FIdjO
eDfg59lVOVxzax+Sk3DylxnE17WKQe8kI0/1CZI5hQ68IhsyGZiJA4ekbUxma+ODatSqWwRLS6dS
Vcsx3CQs4w4Km3GL9RpKQ6asqa/DZ8R8cyXW+KKrBQ4VJVaw6B7uCJTPk6sdlkTmHgl/tGE+QZCp
Nc78kgcX/gDPX3jurDLBjD2mbjnVbzFIvlgSWkeRzKhuoS7KPppdNKoxsURb5o0a5ijKlyMifdP3
xfZB1ycSdzmrNQW+LOjYU6qrKObfHN98a3dlsD+jIUpEFeCqybWr3Q/8iquPCdmKxHLaSGQVaEWc
pv+7cCNeRDMNcqdGThPwwmkrxNfot67mtnmwRaurUhOW2EUBfXOE15yCXDJsogvVQcLIlqjf8XSB
phd1mLPgsl9TOkaLWfr18+OpuunMxhZ+JFy+0U8VxR0sIirNxwCgiSYJoRHO4JBAEAd7tsrgI8aN
En9opC6B6jogd4PLrdXxjkzLHvLa+z1zJPvAPC+CagDlPe3lOvBGLKRWfGZnu9tBcLDTaDc4d5f7
x42zYrzB88yeHL81vNQmEbBFf9tWp4Flwf4p82XWBqLJoAvNi1X1SItzcNR1uPkGZkygza4hm1ra
5Rew7HJwcAhNjP4UyLk5UXatDLpk8FETOxkN8qI0HNbn7Ewou4X0R4jGsbz1ffcFkPkzQ7B9FOof
PddhE4blAvTF5bLEaang9MzUgq04CfTNESIkyukrU4M+8vwIBwC++42G+w1DuLMZ503gBq0YyZev
/ZKzQCBBcisw/PhH2TE63VZTQYJWjp6Aie6nkbObIX7Uz+I2CW+fLOx3uIE1LoVabpMVi4xy27Ft
0lyf9nN24fJf18DwjGvuFqaj49q6oJAdSiiUKZvCuR50sS4Ajr0PjxOPBGbnSmnPXVcbaqqBLeG3
k7ao74+0Y+yivkFm91lZb+0Pkeyhwzu9H3hgU4MibB/tH2ytsghVhZPRhNbAjTSgi+BS7TdndHhF
Krin3H/xe5ttUAGvxm2H8esPPBzbxFwSaQGQUJzV1opdfKf+dhqdLyGaS68bRxMltNcnzZfemG6I
vDWzx8XxwFKAaUJpkw5EnifcMhSc3ROYBppSBdgy4bgJw/XPTpzHwCVloQT1PQ2GC7a+69wE98vp
J/7WJKaEzdY0lkMlSIMOfTWvqKUP1KORDnFw/78SkKWkp1NQ2+uOJoj69aZRzFpnHZCPQxeOCRLS
9TK3ByGidlH9xjIHiOYiw4pmd3GDxlC0OHZmBpYfg3E+XAKEXbaE1//5TTF8ldcHGDYBqyTy2oND
rULUpJ+2TbsnqSs4PEwXYYg5h2XnW3k1/W+UW0EHfPdtBOVnEXNDQ7pYlwu1+6Qg0lDiWMGHpB3P
6jpFk4W/OP46xV84gDqTiX+esBtF17yiUAFbtCbPnInPQgmtQAh9F5eoo4nx0xVjKWsSWv0vfUd1
20GnyF6sxILm8zpBiSeyS4OqTtnlRqt4dWFmRbc9PALadocDaOKBIfbeVRctIGGmSVgxot2sWGd6
9SJf7KzYWeMoHCsGAoDHphh+qSTBfQHHK9nVcHv2iOEQD6aK3J7PIBXukJsM4onSoXyzSy3+Thzw
pxTilVoqb5i1Wqk9Tfobho0HkckPcIS1XM77XsnmM9pISD92+S4i/sFDqkEi8QsUrvHWmqyMeoLZ
U42xGhD3uDJYa8MT//twdJyDZ/CTNhACuOxRVRJzYMv2ctKhkOx7QADn8larPaePtWGGNwVNyRX5
ySEMufXWw6YxR7ws/AUmxixxNb4LyJPqP0FpR1ioMZaxu8dv1ZvmxecPaHwk58AYCyhvIy2zlkT2
jjPHweJJUDbm6QWhMBkQF/p9G+1GlBMQhITSZgyxLEaXrGiXy5RFm3JnEK0v+hKdf2AvpyYKTnva
9dE6HlSFsrzB0nfcbA3uKWrqi3woeVdrQrrt6xsO4nOOq/YoyL6XS/1ip+jPAI+1vhmDilQBtku3
k4IHW3+PpU5N7KgqjXVgnhCyrXdzlnlMr2UcbgwvCSrsYt9qEtv0zwEnKWwp3zFGzXKpLsOIL81x
TO6+fGjyasr6F0Z5wZ5oY90KFwS9aVx3gFj8/buO8eEyHWTKY59gmFYWRY1jVb4QN/4vo5xozG90
7MH9o10ywwla/SfAEltpEXSh9++9bLz4Lw1GkpXv4S4W64+Lnk51cwlBkmqBcg10+NG1a229ouq3
o+BOcoK68gXtLz+HEndZ0VnzC0e1ppHlTEMscw0c6lJnxD0ub71EemByjDiYM9jyaJXLIjVHdDVr
aWEZbiSilaIYhDpV11LvSfqwjQolXX6i5vYqCuJizLMLkXnhqc5JCPRwwVqg02WMCdPrAYkvgcLL
1p3wWsw7A78AdS8T2+yY5ukXfCgXhI5Ui5LQwrcXK3HrzTj3agMv6F1lV7SxJCidEannbVCJ7Aox
vajvro2Qr6E5cz2wgak4j5bf/hQ6LmbRRGZrbYfTLRb89sAUSkvezVIBaP2ByYlfFBgYrUokP/fy
2wzHlh6e40zJ2Gw3MTgQtzHrNrfmGOC2vlZQSvF4TBqU/1JghsHjdtrmY34Ramva5gY9TieRtjLD
zUYYnr578VdzPEp0wwEcQnfIjT3pg4NRrt58HRUUkU41LDT0KelINdnAP4bDLU4JJ2GAHWHS8GSI
a1BoJf5r2cvlEnI+ljdl5xookNW9iI+N1HXLUkUhZA9kqODeJzes5iUhYvdNByCbpGWGHLRExivf
QntOCZruJhpCRXNHUZuOhCsZWijE35hZV1tj0wxi0K5Gp411cwajqfECvZDXTbrIGr/eL2sR0ejy
RMnZJh8QiUBbyrWMP0lJmt+uiNF6GRSHcfvPEBWDpBe3ZuzAt1FtpdczNS9UOSuZ3V4eGgWfv9fF
uSXI8RvtGiDDe7MsF/qtq0dVmU7Drk8uhxD32oy5KYeIY4aFEZ146f19I21jp+UTvwIibU0NAQDe
2FSXrlUsFe8IajAA/19mwxIs3Zxgo2Yi2CwxEV9866/vgtYlLAVDP2Iqlp6MscQKUkNVSbx/+xLC
mVHMfCVVLQNAWoZsmu0HluBAiz/TKDKXOKRGynumze63OfqAeaJTAPE4VUZp9ygBtla+rLZg8ONy
kIAuhznJf4c1IOM0ws6AB4+IMf7LwnLST90kUEUSIHIBvpNVRPwYYGwH9yqC9yVxJzK/8CJZuRX9
hAs0NVBCeY8TlrbJXe8t0ucBS79wk6p6EdZEbkPw9dOrOAfbbhUA41ip2kHVf+qL44SIxjuX608P
lYCVvhHZmeh7xiZ1gjqMk2oI/LCzV4iLgU+eyQiUpLhHNuig1ZyyEB1kRLj2QGxCzeGBc89YpDEZ
UaVAgXZr9YYlZ1+0x9Om6wpkmJNrjjWfiwwBDEu740/AmRVqACQKPK7gBrRecKeDVM/opLhQz8My
gl/mjtseCbKqyM7RJupKICraq+XvLlAYZd0xSxAlLmfeoZrqDgEjG5QBi+0u4lnVgMKnbPmXGpLs
hhGglOEeU3S+mswXAeCR8UzxH25OcYjOKX7LguKXaw0LOf0g+Oor/AISxyw6PYxe7tytHLgEx/2N
j3KSuTB08j3dRgkFyfNYw17GfKDWVxag1SwHZkkN83cTSg7ZsrD5cVODTitCB4bKdUJLitO5vZEj
XNyJjsZntn19x3RW2e9/VguOSvqHUqUWd3nqzeiDTpvPMKXYDwISIxyVG5bMEAJ2Fkbc2gfdOxLv
DP2t4IeEnG7+gCYW3WEX1ZCDaGOIW1Ssz8F8LoGHhxYmNL2vLH5k+Dm6E8wIeoCVTl7OeGIaDgPh
2vI9wFcOqjr/Ve5k2E1g8AzOZxc+rTnb2qKrBZkYPvs7jN4Kxd/wSHM8yL8U70maK/5kMUHVssDK
ko9pxvAHBGLhEDkC91AUSkaJ9vnMFW4Qday5uyLPMYcapLvMLOt14B2Ytd7jGdZ3QN+8XCnJnctn
j2HDZC1cmeFkUgEJf2h28KuJyIAz81cu+1lM+sdu669XIiBp4KZl3afO8KgJim2uROZ9tcy9ako8
LSg2uiHg/34AS8EK2p243UxcDtqyH2+UM7yA+QMxJcayZg8XGDcHHX5k45jXKJ3NDoh53mqu1Cy6
wDu8rpkpZoViMB10ue3WlTMHIE6QGpbGd0kgrsgJvhMlgtsIeG8OnxOHofNwqNtBnDqngBZYichi
UakUqkYkmb9UUPNxJ5n87B+vkNh/8irFuwW/j//ZF6a5Zut+mmJ3u+HhGEdaniElNpgi8LB3Wkcs
5gi6v1TXe5F9FjN1FfKg3XmZnywbNCnnHnSdD3mEUUSnZSlOJJRW4Wz/UMrTx69b96E7WROPkGto
9AS6RJW9nttPi2PVOyLEzCyrFCSSs+QeZKgAae2jL72eTVfpAwfW/ab1m4jevYebIcn8zyXlbTKw
RnOW1xXkeYqwwenGQhSgFkzMI7R+gE1CKt+7Ts+0CaXpyHB7oEtXF9QDAl3vl1OLEkjAe+p37wWm
Rxz3M6A2mZ7YvhucCZvJdQrVIUbO5QwkjgoPfWRKkJl9hHNjFbamvOuLWxbEzEL3JGXh9voVfdgp
ZYSHs2nPJqINnPa34In5WwozR9JOO9+3YnCp42VD2hP26XwYp6aBAMcTX3lYtaQx63LpCcJr0v+a
y/+AcL1V2yivoft7CvLEEdbovQwm95wSQF+uXF7Wvcn/qTN8EGr6VdSICfVs1K/jngETqgOvifTO
JPMI3kHwxL/IVGyysRriLstuHm87Hb3k446ETdgs6Q9yihGfghrN52yYF4DcqRRgNtvAdvVrWLth
BygD+uEoJKZyP5H7rX5FfnivoIcCD9jWAazQOE+IDhcxMC5oy6ucLxSPlUcqXYjHQ3/NrI8NLIJt
ZUpprIUBKdnMYtANeBZFeGJfUqXnoCyY8McQ7RnSSHLD0ANlPLUF+IHcqPOZkTn1DUG1GQ8HF0P7
GlfRuY0cd4o9zpMNYPSvnwfW8BLmVxDwfpHKNOOAAVtmnSG1HLhEOixq4oNmLV8duuhuCSdNRH1P
GojrNc656aeqaPyj8UToj82X6zzTturKaKYl/iKjikcFwlG/S2lQuJDQx68Q2DIuJbsMk4uSCUPc
eN+opcj7NEI1gzHcmA8Sd9ArQ0P+N6x2VNtEc443X1m+AtbjaNV19B5Km5HCmbmRx+NW6RxtUY+9
KjQk2bEu4qt+oYNFKDvONpCfOFuxc/0R6BeEsUyKkk4ppBAnM3aoxFZIaYDKYcEHqdFte+3MShUs
zJdyWaZvZL9nCz7hEDUEJylSAWKwNhwC+Zsxl1Co/bbRalFrwp+15M+CuwTvD8jDyxigiVtVCaXU
7Ul2A0Z02lspEEBP3cCCqbhVycuQtFQwbUVvvZF+pmQ/Y2xSUaKqOvQh262ohJ43ag9Z+c4yYJ08
IJ948JUQwhuoCTPh8FaSvGh9UUsNbFUHLCZQEz4zfEpn+Cx084mbtI7NOKpMLaO+aqei4ghZSJ0O
lZcYbDIIHtLpCqcbcCz+/4yGa7N3DXEzicDDYE+LpSSELDvRfB9nMqDyuiCdFPWVc46q+H/SEqNW
AOz+OeA//bWjR/wsP2Pk5rypNfRVzq3/QlhAJrTckKUUtTnZNMGEjcoxOU4FVytnrngDFJ9gUAUv
jYsmTnS4JjylvubloaOHJ5l1OEjirMZqNfYHnh/gXW/E4yPLO44e9IPBkaHhgbwA/6iR/jC5YT4U
y759z5WdxC2GqWUygHjhuWW52YtCtlEqfokDa9g/xB5FHw0aWu49Iry8doqvGEzl/tM36YbsEgIO
fF5USDld7zQpm5gouayqLJtT+YXPJcfnSvHN2tbyAB8xE7XUXQztNNXEhol3LZ2tUtBevVNnjx+e
aLsmRqiT8qy24Bd4bZMsp0xCWF1xWK71aT3cuBFqOn+fKUvZ1LC/3gi7C2dKn7qFTx+3D78xeqVd
o+sTtSo3fH2KbBcOxoDGiR7bqkh/cncHqTRIFtXcT/oJTspB2w+YTD6fPCm0sqhAJuIn8m1huQUr
dKdY+M/K6/tNKFqTtzKx8CTVg8KU16X2n5pKxl255U93VpaUp2DP658G+G8zaAde3LJ3vP2SPV8L
AGtWZUjYkf9Tyi+QRqffXxnvOUKMLi4f/Knpzmpy8P9C+TzWa5uRXYt2rwAp5ppLOlTdVSLG0Jfy
iahPRmCd3XRpexmxyqnBNkdGyA+f9EHW3V/PM5kVklZEEzM0BJnwfQCqW2qX+6ltE1MJ1fQDjqFk
VN98ziimF5dTtLLVjslgNF7pD4mRQ4bCo/g7lr8/koeXilUS3/4qd+cVRMavcrZ1na0+5iuETOL3
VGKHm7C3E//+W2lK21sNm91mygWi6NjA5fJkSTQyKyuPaqW2QxKs237WxvJ2oFGem2RaMASJ1Hkg
5ifu58UuizNpY9Km0Rz9Ekx3ksvqZHAg3m6Ogi9wXQr8A6xte4P1vy6F+Qum9RcXrGyhdBqWHe9k
ooXmEHaVlR4kfr5W/ZjynIYam2RFuUhEYkzGdw2cn7rZBXNtG48b/A1wK7aFNsMS+Z8/ssNAZcVS
l3cFkBE0dINMbq3n1Q3QsRGW0jse1fx+hKsXNR8tHa4/PFpcRgRO5+e3U2Pj1sZ0HLwPqY8W+iC2
5vmOXsudca+TDZH3E/6FXFysB8yayHAfkj3Xd12VuAgq3osalIEbUVvPP1no5PmuNfUdnkcvGjzK
Uv6Nlziy6MTQ0lwUTuw/wXIdzwG/tlWgrzdHH6cF4s/j+pHnfqx9+Hv6U+tqNzBpqh55rP/WrHVk
0ITTiDGUdYg7bN13wzjEK9RMlhI4rcUKy/dnzZfJpouniSxcU4vtfszvSbosF/E1oNijagjX+NR5
2H6jCWU1s01kfWi7Gdnel5pTA2dcyQyI2m+Ifx89spMgJETRlYcKIZlB/F1w0vG2M4h3DD/Qyloj
wTAifVUlrZmsvPtPfiVXK+NhUbfvKp/EjeWBccjNL4pI7EEW7t/oF9sWVef/l/nmyhFWcGOR15iG
xgEf6E+BsfkDkGn9SZQ+Lc6A+QmcSqwGqvJb5ujOK1BJCf6YUwA0yA1AqPe9EF7ICEaUlkTgT927
8/3LoSCvhPQQt2cI1HdNn5gXlXy6ck8NdUn9O4n6h2eK2NYIE+xZ5m4vT+oshh2h6IFCjpXSPWNv
ukIehFlMPVMlzaJw+oOt4wHLgO/RdogybZ9oPsz5hazs4rnjrCAyumbN34b1QKdSCCdiSMVQbFlm
AaDu3X6+hCmKg1/fGnqJFrdvHSQ+b6EHFu30aE3IqbliREOO1XXT7ZCcBS5vjavUnWHhe244hQYp
OeFCFHROOhNDKdQsa6UlLeVzynJzXFKi8Gh3Z27a8xRD2U2IpO5kfeimYp3s3gn/v4/WLo7gdQTv
iSBRef83cKcnjz90zer47TDzp/jsLVAlUMCrn4xWoANNo3JNtCvQD75+vH9EUwDqKCFHb+mseCs3
cFsc3A4I0bJIa2jpIkv+0ck/OyuetIFgv2HXqPTiRSe0ENLpz6Bew/dJi+jMHIhGhEDU3ZhTRLLe
mFDh18gFNKSkawfXx65Y2kisczNUX6UvHNG7tQod7hJMWcc2KzyQsZ3WJyRQQ1QeP4jb2XjDid5z
7iI1K0PtIMdI+jVE69jMgNfxB/FPfPPWPsVA2PtuG+q8Z0dap2DP+kd7hf/hPKI1rq4oQZxZotp+
rdMeFP5csbNH02A2Pnb/yU7HQpsCLD2B0+S7O9sOIrwMTDvAnRM5xdYjoje5q9KdsVraKADBBSVm
sr2lMga68w2gOdZUAwNXdqGWZfDA/MtzMZU23pt4kE9c0Tn1p6dJW0zJsIrfPgemOSm9FCwS9VsW
cBxTuGOCYoEx31FLAXvRZnYwHuX348DtpXyKIuuZRAhaVag8o9Dss6foi0/NiMQ4idcyr1iZWXhT
GS3EqTleG05D+GRFaGSFjenODsaDq/xRJcx5WyLth94Hf+YbJ1TfrjKWfuDg0CaGeNYOsJGK+EP7
osQiCp2tcFv4Xl9vrBPduv5TCLyQ14CoHHDqAuBE2xWBfXPraVJ8OrnYXeCneW0N53VrNsH1dbe8
8iiPYoq9MTOLDsAbRMZUEm02Zeo84B3le15UG8IrsXIcW0Bvg8RkhJN51C7h++Z/iyfIiGkqVPn4
ei+mcuA2CLRTyATU4WYQoSxJ+CuhEO1EmlkLf+UyMC3Z+Qo+wnkNzy1fid0Go5rhR39iTaL7LGFT
yB2tAhWLFFUpvGN/AwMkUJr5g7eSfMKc4BgvhrSd6Zw6kUfokF0yw6RE18tuHZuT8fW/8StUirS9
Xn/TbTpU/VuwnVGo6NhuHbkwlB1RghIjesTYnfljsRKjVPGKt3sdBYGDh2hFQYKb95ttwuWSfOFa
aEbLexm6ETEqKjIKwJZJ6NAT8zijtM93i5inkjT0gYzqaoz5fkeZC8DKufdsyu9f/MImb1fetvfl
JelQnsUdllBWIcdQaThSDTPF05UFXYhjZZkbZpN5hx05MpHvYJDZQLwxllHhkmDneECMWvLl2Zd7
KcPAaVOUfFEAS6vKwbbhtJpd01dydtec8FBB/eFWGfYPqf/xlAteWkiAclAv7KhV/rusQchpUHwX
oZv3MZbb5lBIohPquthLA4WsEHLo3Wo+ulwQXDPqHyF/sL2ul7fmtPWVghOzOypjHc8Qo0vaEY7g
quF3bo2N9VpUpEbwg5x6FLkSs2eU8bcYvHhjpC/Um1SSNJsqaALUhIJmAvAvlcglQB0H9XGmNQSs
iDuz5yXzXmfusy8+d3t0efPd1bdlINSage6PikhrAE/mvshJfnstRZAEp5qseeBm3Fmb22tTCCG1
X+xERFs8W9qb1wK+K6nqm3fv2EtfbeERhzRyIFjdj7HECgvzpDXNqzVXYRqyD4v4VIqESz7v6RB1
1Y9yn+3Z6Ez0uGX+A1QPaQOwtkz3oVP+RkZXx7o3DKRd0fRqORZdtv1IlifwbJZYXKDmqCCx9Aba
/8czPassMKW7nSivdjFf/ELw1UkmzKj0b3t3rLzLB5sDlMyQxDH7jtM+FZDDhTAtbGr0jWTP1kHQ
soGxZ8jfISGqWHrOzuEzOzhvoioatLM1oV5DIgPjMgHIlLWCSWrrsjMpTLqiyjkB8hUGCdvLw283
++kSc7nRHE9YJXNCNNKno86F1R/8LY3lZJ8GinnxXCVR4RFnxyP6XPtU333h97Y2371RrSWwZe3Y
IdyVwC/tCR8EpjYnBKDkVHTrG1JgeHoSMGrmy7UoHWZEBiX1OJ4/LvWl6DBv6Ysj91LfSOKBNkIM
7elI7Y0091HundfrJDgTTkU0WCTk32CnoG3aXT+da3nCD3im0wLt18QbTxWV2t/AtHUep6gGvv/f
NCsn5okOj7h1Zv3os2k6/8jee/VrsCygJWV1goKLuEXdtPjsl0E+LL6YSozcZddWEgk1IjOlJXLA
qdv3xOI7zZ7Vq+AZQHFQDXZZGZf+z0UcGGLMS6DNsi99VcrEXeXe5cQ7Rz/WTLo/9XrQ8D4+snXW
X968BaMGUw73phePTgf/hEVAQXCb7Gv88BbW0zWwqWFQe0AGht0xPqyg7L0U9Xh72LeMVG2W/DHJ
//+IxBxyCO6Brl6gFiyJ+5FfcQrJ3S+qspKeudFwkobP7ry+7UUD+1GMcUvcMYYLLvj2rtUwhDC9
xIBnpZUhWA/iLWm9U0WKKC57iERQwlXC8ha6SrhK4docajM2OWrKbfZNVPyrfPSOKmQ/OX+I+B+c
KRx4MiZrlSFSKwG7lDqDbcxlK3NndE//QA4jCk/c5Kzq4wEuOve4dv5oQaID8DWMz1/ZGv0GIDMv
3Cam8snxbgi6BvGU002EJGhWa/JZ6I/rZACPn+Scl5HFqT/1Q81hzsnldKYoQ6qwav8HQ8ldBKa9
+qXNhQ2R59v4u2wHwiVw2Fvd4P2Y/GrT/SsC7w+RSDm/XCXComMyeEQBYlXzoEpbhZgftvb5ChTR
xqnTPngbgOpaRCuPepmSCe6qcNN79okdxU0LkPHtbYvOwxderO06C8mVcH3CfKqfQ7+8k+V4IE4R
zsAO9YlJLlPGIrMDGygNAK3hngJpE4eg6h9QIG10/3Ltiiu/EnVTzpRE75I/S2kY6TrrCsgkyFI+
Fc86OXMyfmlpEkH5Pw4quy7ftCXlKv4v49ECk9bc/BcC+A15yq+e0v6XFB3m/Loj9sHBuuoH8FdN
HWvrazpMfR0iGgmcrNng6cNzylONBppU2smZEWLYuL4w4mdK9hRcYwpXB3M+TxduiFwSeQT6YKyQ
zJ1g8eYbVQ5aH5UU4kXimqGmDPlQhAiV+qqQjS84tJGpVgF30Mt/gZ7dmrDn6ZCTs7aLWgUxAYCB
Arg7W8cul0+a8t5DGDeb0Mla7N7dHIGZJFuLEnEhf0jfMilutcZhVkt4TcVL+oK5cLAFWIrFnEeL
vp0AwuTnMdr1quzs7mqZPmkeT3zXWtv/e8gxs69pU3UPy/euNjrqV8uScsf/RBWV2EScEpr4yN99
Ts6Jy84MjWWX4RdlQ5tNXKJfxO21GIl2jHMaHsEh58AwwJKNpnV2ygCaeXcq66OlnniI7IpxcY+V
dwfx/F4mx0aDzANj9RgHAtsnpj9wfP5Ly2XQJsU4bnjkGSLC/U1FBWygBN2vrQFTd9viDyhHPj55
j9qFLYimIgYqNCeVR1X831Zhl150H856uFIBB0j7uLQS4TfZ0jbamqPqqDcOAUAvvNEvHaDo/Oku
QSkLO+P1Gnr5Y9MmPCy+d5o4IZL7LmZ7SbYvaBDWel3rWbhAJiVXgHEZLsRf5oWc9Ih46mOuiCel
ZEAyeWjJXSm74pIok1qo/+t0wzM89OO5pRrWG+VoLV7WbeK8rGq+xUj+sDIhzBzBCMFqNkdHlePd
0MWE2n+gkDf9WF7knZ936yvlq6GAXsYgWiSzA86wnpr6HR5oYbiCbPNeuXUBI/qwvThGEAmZ0pzv
ieeiWz0bNjRXynVC2U1SMCbWwjikt0iULIoYfh1aIicLVSy6LvgVpuZvnITAFenb8cP1Ii/se6an
lEZ0sXxXJ0A75ZQZmGzgXfDHOWbUKnYht2KL61wkFsahXArEO1hLsGELDXWwmOdP77l/OmT3Rv0r
sP0kqMB2nv3OusNh5iP6ls5y5mVCDj3gZBxKrJjNBxBkEQgIBy4/CmoCWb6vHdFSqJwZbhjUz3C0
FNKDD/Dl923MSpqFO4XhqQ0gbE5+l/XV742w29pvOq1SOiJsoaLiKXL15jZyuTHBQ5N2+Btuu6Bi
nwCcFmXzxTsXFZN9f+u3AthPABCl+7oK5jT6OrwCHvM8hBAx2fGin1FmirfG8AJwZbsG6IycWeXl
70IHxDE9lQa7ktHQw7hdYXQ5HebPNxljbDwG74/PeFPNSvSITg4Y7IfhabpdtjRY02Ce9ZgLLNkl
mPzVOdleLpb/AzWLxevuhJABashwiXEj1XrVJelZhA1diPnatLYca63WrHfe7bvJ1YTmalaVU+uN
FGtPBtv4QzTBEVOb1RKf8/grEm7djRFkDPlvKxb3tjGVVtT2mWgIRcnLFqr21PY37eHPSdvNW5cl
umCj5r6FdNfBSGf0VFKTHas9sKo/5C6rtzIGIBTXaIhx2WSCd01zhHU0MSP/g5b/nuL4pjwdHoNQ
hW8WSaJgwThuUCBcd5kKP+ypLJoWYoo3zHhkXF9mkGrkifGF6DsPq3PrFItZaCxg+5fzF6uwptb3
yfJp02l3zDe4ablTIBHwuh5fVe22kd1jCcZP0GngZOgQrSAQ+XefHlutmQ7lVu1ElpIKZuDIxu2W
KQhbRt7ouhhYjgLA96DCuWSS9VpQYDGmA2+EjqAAtaZy04O6BjaHjKDEIvAOHDHCH6rz8BJakH0t
9emnGmcsX+6Rm3dswOBB5mbJzw9AojyifBuMAUCmfsOMskzpNAe5NFIpDe0k+CGMjrc/CZkdRLXj
Z+h+nGt3qBukIORcKdXbMRU4eFBa0i3135I8ZVCFWGrUkXZelNRbzrba5KPSrOCmwLghLAPmES5y
6OzmzZvi7qoym/vIIXLb8NScv2wsrvGeswMC3+6vqlg5ygSt401i1SJKKsjNDkISzOrsSg/xAreS
ntsvKCZc/cPqA6iFieKfMoqJiyoPLujWNiGvp69d0uobgkzpFLtIKtp52vSQG9fdoT5rmFpPwLDt
oTO2Q+an/R7VU1gVP4Eluac1PH/g1bINREdpKlSLAhMHbd8EhMPu39gLE28HAcdfuo0Y114F7b02
uJUd9b4iKO/jfRrORKM2G7W7lbfkRr/Yzv7NDIfGEThw4brciBeMABh0tsO05muI0JJW2gF5i3zl
+ZXJwYLMQ5Cq33xd9YKMECgqJlsWYRxDGdUEx/uLey/modlTf2iw+lqz6cMsYJBJ0iWMr9+viPVb
tE3cqKqhK8tCCscZ447g50d9At/bR03rye+2dax464fQ81UBD7HwTaaebfWd1zyKy+E7jdy0uJRR
e1qP0RBdAtZi3LK6oQK39LrCK/+JY5T9X7xpjKUtzLUqDQJEtJkyNpb+/7qkiKt7RLiH2tJCpc8D
VX4yyEOFPKX7u6shFYoRP/fXB1cD+qaRMSHVNFUXqj0CU365CNpNleuB4pS0DN67b/db54J7WGLW
n/q8za3g7Ev7/Ipf+aWGQRdlKab+xZq3OyZ+V690Yvfe6cn/Qrq6rRxRniIddzzbLmEON6tV9KQf
QUOqreSRM9csgCQQlAmSavEY3OeLFJNkTWgcigvp8CPxHzKgZiac5jq2wfDDUeOL4AnGWOCVqXtq
7rhQNjSP80NVcxpZEFNYh/QuQRVBa2r5pLkw7mL0kRA4cvMCyH8wcnYWrUCrTViW+J6gIn2zNAv/
70+I0+WnNTZTJyOaL210yPXSlY9PFAFHxJ/HPkGZ72gYJRRWUrU2pmzaZD1XChTLzEmn5tsOpQMI
pgME6PbLd0aZ2ktClZKZU8GTg0n0FPGMo/NTEPKcwvKEXPYqRCnRdbhlcpfQl8sLyG4ySE7JNXXo
QXAR5A0F/RcXhYuLRTOGO3StCLwaCgmj3WznZHi9s5Kz1GApjCFkcfWDL8C7NVqwsz8sHXVF7K3N
g2ybwA0oQBb7S4YEk5PhQW5W9PsHO/PSOoWAl7VXexzrOcAb4zracQyehPj+Kq+tkjD4WwpNLNqb
BrSt4CRQBuvJqAI34jBSi/mBNYSBGpj1XXl0ssZKO+tBqpLSES3ZcLptEApXibKmxrN0cuzpNaE9
74G+BlE7780f7Q8JXPtMOKe4DVEB+a0hHuHGG8+8B0NB90sWOQMMBr1PHCJnbUHqz6oodNW522sm
utgUpDqS6w0rfCwCWqEfBsnbyL5FjVd1t6tSe9X8KIYTKvsTJ+CVnDCE7z5XYftim707rmQePrW8
zJoRXtJZOGZl/bXA6b8jkd5lUtLba3fGikPJ7BJhAVL3Ua5sunquBPoWtJYCe5klqdvHCD8/BR9/
nElILNhq2fyrYLRD5rLXpXVaN28lOLclSy1kLW6f4gGs9dnp2O7U7bPwT8nzOJfdlHyqLgLfFkAh
UBf0BDPdAT+VANkaAMvlhXruCL2Sz+P4OvIgi39+i+aA9Xa1vRAVls/xtzVrATfmYdWAYwtRTYNP
qWTbnC9vxru6hNDc/n9kU7BrurUp7DmlUWCGgNjiwrFgpDyKupyEwPkYRBjFt1wLKa0mbPwnvZg3
VB7U3Umi0yYbJJLY1MhjOgt5IlPqDfPBceWuMDLry4jGNsyNX9zxL3KwUUptwjOzrxtRmiI6lhXf
r+uOkV9LlAY9XxV3v47TZx/xG1a+HKakshZCSmXlFLfcestc6ZYK0/d0mguPQl39F276ZDufLY9W
weV3lWfVRv/mVhpfe7D7Z6kj3wgIHQeftQp2RUC523q9UlW8q3qapotHLxcb9ryNCNDZaO5sF3Ez
6T4AJB3X4agMvU+kQSbinxSMC21zfScnsi6l/myUR7bJJYfuX5vxrYJ2GVEzCmOjBIZyZxt/nf0C
SJUSatBG1THCV+f+vtvGNtVsyYz8E87QJbbkkv/drj13EMEx0ab5fcUW/nofJgZuIuVAkTpyamIH
cTiW2LqwwBd4/bs9hlZ194A12Kseu/P8FyIjLx3vXWukEPD9s1jE1vHEXTBrmJ4mIvALxGS8c84k
bETSWo7OStN0Menh+e+cwOP5+wherKXtcCMdr2p5EF55/D6PUNWGZVI76vS+TpUlNiBJP+MVl1pE
Ur4+T2UQwitz51gb9hBj9gHWQJ5rlGlg69cRgz1/HaVTh1kJIkksV41HhiBJGsErgxpN07m0mK51
CY/6IkrKK6ejiWtpRVzv07/qzvs7YvzdHTVmbZN/ZMWYx35JZVP5Bc2rAybX3r6d9C0INFopIu36
3Ed9BNx67MI3PKoQ231N7eHjZxw2DaiYjTxBfPJC/K1rNKAkDlTkhH1k/C+8/CNXN/jJo+y3B/bR
zalcGXJEA18NADoRrdfknt+q5OUJbQ40fP+wRud0cxxIhJJFqvQtoIEWViW8A9FmhanUEFBR18nZ
HJeX8O6s7LN+vRQ4J/Tk9WAvBiLjja7ZTof1ooZ3jkw1G0yfxQIG9RDvUnFGvHLuAoe00k3CodeQ
OovxtZ5HVcdQn0QlwC+O/lqHYaCzJ/zxUA+R+aqLPkF5JQYRNxIvk5RAJbM1z8GfX4lF8fLMWWI8
qbTp//5/ugOq/Qw4O6KnqtqKvOLisimBBpu7kje2qXOc9bnqi2ndSJLYjHUdtkPqu2RTlq8HloUs
p8UBJ+n6GYDM6ZjNJVhNumvutyrvtvHy74ddhRdVEUH70Nq1wS6iP2R9R6vIAXOCee5zgGJ/bY+a
RjBudLcxAUwPrilzx79tH8ci6Au6CUy0tdB7LiwCTpGWJ9Y83ljSP0YTmLHyRp5lXzyesjq5BGMm
08ScnIMxgn4CKttDtWkkmOc1q5fRF4/6Kxc5/bcmvN0/JB2w4Ijmo/JomMXlyxYuWgTdxUJQYbt1
htfDZ6i8/qIuTmRN3s3HbkOX2S+8ZYdQ19Bl2DxQKeIcaS5n3NC67wRNdm/g3CkA+Zi/jC+1wcXO
SnDB4hyQSEd4Mkc1u1ODUpF7mRSZq5kYxJkwOq4HofClHPq2aBgIBugN7pyqsgLL5GxoWBUQtfR3
H7OFksgSFMz4yEVmKaZ/WrLFtqAdfvVzvAp88wrdPJMUYcTAPAOAjGkZRlhkPM48Fo4uMGnWc3tx
Xvq4YQJkZXjWMTO1RsaMoxJirV0zXivihCulIT0k6qoOFes0qbHpEHNVEVOJDzZnLmnlEvt/lB7J
oxs9PEiNye8Gm4OtUBcD+Yi7itNHAXbghGEB1iOmocT+9YuTBbyu8d0Jyd2RznQDBeYeOQF3xd2f
cmUMQsfuk4sqDgV3fGvN+ck+/qsG7jgdpxn8cBaiMAeFlptqWrFafwumBWNxzh+8VeuAUuSMzglY
hv5wNv4lqdIKkFDeZ9KNgdYguBiQ/3Oz5Z4oJ26yz3xvp9+Sxz1/aaLI2CINwu3fzZM9c3WcUwVt
Pik705gSuyrWk1uq2jeRZSPwzzqtXfnQgLCloICjOCjNRLfZZWrj2zdSswcsN157uHkYxEU6S9hZ
7UCLI859AH2Ma/16xbr+nvpFd958kQQ3V0X+KNunOSUq5xqVzaPNYKLMUQuSf6ziCK4zfh+Ho1fD
921Xl93+1b2E/8AyxZ3OFqzgTCB0aDEtmofd90d8gWQgGt0tAzqgafv2NDcte4sOxtCGvcVK4S6X
n+LFD+CAU6wfiCCdVtNkTdgwF25V25iB36poc/VFz7L7KVVWpv/vl5PC/scCx2aTHiiuXoLSD81B
Igg2DAwTtpdcbILbsajLp5A3ErkTnqLKryIpm3ZCDZkL3LNSGDmUqMiByQikuJaVt5RTq0yLIGCS
5hH68v9bG8XnUz8OHlOQDvQD29fomggX9UbAUomnbXrs7Q+r780jFLUApY4Al3cBuoVrsGRsXxdT
wQ2gkoxXAFRspTlsR9bgTXl526cStsFUV1Mpk+imtNBo2fdsi2iZK1F/wpkn8Cqf378FZTgHbsVL
X3dv9hp24xpXPrshxvj+Sd9BxYbRTbQ0H0ZthgcRWjvybz0ie3xGH/L+TFAahHveriFXdDeCuCeq
EJXxFu6ep0+Cud8TtH80anDwFdVoCILADELA18+oAa4uD+rTFxFMxN19Tj95WSstF+GhwEGI+lP9
o2E6TBuzNXRII+qqxLGHiHwIgqiru4CLTzbKIrTi4mVkyszzwu9FejjdZ7Ge75pbBd72o1S5V2VJ
D3ScBvGmN98P1TXONPAIuwCB7pRnetNPzKk7BPkssEpR6ZfCcwfeiCvJRUhKAdA2Luj/VVpKVWBl
ENvmatPhnsJxbfGlcQw0png8RYfkNeLZ65y+f9tlUSq6FeScef0m2X8s1tbZfc6NKjKroNDK0lKr
OWgjZEjdNldqCvAdJ4Y3FjKG/wIzGvmLN1hRcsbBJTpfcFi3kLG5zQNp15LVcatYW1JKMl3vouuH
ew5HoC43UbLkLHV+afGGtL8TpJ0NbZFFoSua5pw/XrmG0pP32oH1bIrumJnll9l62wIIXuBCP9BY
WleZLRw4wjAeVkxD81vkHdyIQdXek5G40qBqldUPoFF3klcVcirQvQMOF/SyOBaHcL3DSc+IALS/
0JBVgyp6SC+KQj9cReHe0nXybnKPVOdwwuno/6ptfwY/bJjdUA8UrdmQZDefd8TBCMGnxWDXNykw
hmGtKBflK15ojYE1AlAasCuUUErSYMTnG2yRUvJh2NGBJlEVXCngWVd3T0EZzWRafqkMlCR64b/z
fQ7B/oOzvb8MWnImZSLm/ECOa9VQPjK5HyGNiTUQAGwUXsqcMUAmW+qYZVYpUEG4U1j07a9JnNA6
PEUgOgW+iXlWnSD1UbQfR74Tnqj9zv8dxWav8unkcDHz3w+6aEhbkjLVtw5CZ2Dq7fRxon7NWx30
v/rxlsCZCDSGvybGDn8uaz4KTFKkxgUiree/JPqg/ZQXntxc7Hd821r1AAbNckDnEvU+x2P090Xl
LOYovjo3PxqUF5EQsrIpLzOGk35zukBVmRFdTUy3MRY4MUURMY9VIxQYMa6ts5rUdAWMzT2iRoXf
pvTNQPtgD2lECGlu5O2LwPQxOo5I3i5Agzio1RYyaQEQLBN4JE7EFToAU3J1/BQvO8g0KE6nkvf6
uBqJpL1R6hEhpwO78OepxmS+41qrAzEanN1Vc4Hhg7U8dsrYqOFeS67Sj++GG/SW20XroAeYgmSR
1Xah+f+QLat6sAMm61j9nSrsS+/wZ8QWviP4By189HefSMYYsiEIqpTgQdsjeYRdDbeK4NlUhJ7o
xAQYadhcfZn8uPc47DfbVPvPyJX1wzl//wLZiBrSsw9FqEKHZRq+qzICXjUaOvFdvL6lpQ7jbPbO
SGt7hKfBGDUelmOuqo7IXJCTzr4t04pwF/ZsoLnQFhLrQo9frrqA3eR3JdizMMnD2ez3uH5XoCyT
UWH2sV+d7FcEA+xMMMrFfAl9YgWslHoQP/17T6PMw5HR3FItKRczOVA3e3DTWYNbcVotjr+L1j6S
OHtqI+clKAoEReyHap/qFW+SU32AUP3pzq2IgPpg0bmOORka06gIcEYngmwgz94DVzCp3cawJCAn
YG7N9TcQzi6o/rAEigbhZI9S0JAPm1yWodrC23YdnVG+p2tD7KBzmy4CHjb6vBAXqGP2jazm7920
V0D9E2uL2wsLpe9WVhAMKA+kTiYaKalvTpMw8Aq+qKBAkUIdGyAmlkVVLzAVbWUXOEcDFaIVWmSy
PaRTcvAr0Axj/xWn43uEpXYHBo3Ju7hWm7K6bWhvtwkf2YdBekWlPJJMxzqt2HRDnT/FfubMgBqZ
oy/kNEC9clUrWfmcswEWKzAVrxD0Up8kmm4qYM/jRaWyTopc+gV0YgzYc0D23ASsVaFGsQmPlgce
CCmMeFSRzP2V67ymKawJXaAcYHQhgV+11ob/23HQ68FYPpcTiFL8wFc57YcTurZB5cCXL/1hH3qG
vKwKx2vY9WEiwl0s58Ag8TmwoSXlvHq1v025qXdeKrCr3H7VC0ZeGFMp5p5oYppvXnd3zD+o+UFi
j6WpBli8oTCUm1rV/ywA71SdqcueU9wgXtaPTGOvPbIQc8sqDPeGl+Cknh7ssBOgSWs7YORWFbw1
kidcNUULYnan5y9tXmBkeQzg6NzfMJXKUHWTogI4FOYsAKD3ALAYIVC3f3TK8RFOtMkdNDd3n1nw
OoiT0ry1Awm4SABFu9aHjJNTyKu4NHcLIEqVKtlobcvvSce9JM1gsVX18bjnlrZtomF+OM9hiauA
Zk59lY+u1IhZ+RegPoQE2LwCHGwpP/FQr9zfm2M5ipCthtbVqGYohBdM6bEOUCHojh6expgfoNY2
PJZVGfy1vAOIsOAe8iHKfzw+6woLS3zTS2iIJu7asVl90cLKK+cg2w9B0VBZYmk0AgkiWgZfP86E
Njf9W73TDnTcPlAkBnlr0HWgetMrIObpeXXhHgCPWxkUMhJVafw1lS1Sys4iyKbv0XYRrQJ8JDEm
6Zkm42jC42XQ5GyIpgynX19lkFsk8jPRSxvKfZynVLD/tR9ZolVfXwNudIjMrk50TBrudUVNxll1
nLfyyOx/WciVkLsnASeZDFSZGWkNe7mV+oKbqExquZvfxJIyB96JFi9nXk1gmQUa3tKwVo6aJ73i
oVhg5f8V0NEbZjN1xDsirrSIm+ELSUt7J8abY0kPSuGGfMz4p4ChNCji+xmQBH7oZczT5XcUIHnX
o0Mi84995p2DXcQ0Dpd6FMVYk7CZhpQs/MlKvpoyxNwNdEnJoBjMPjGxVI6leh5zKjtO+CdBOFp1
kXajbWpgWhZv0JkfdFCvekTXkckzSSL+/dWzhuxTP1e3ZNyn2naJWdhHtWMGhuz1IogXz+wIgX01
edXBHO0IPLOfcF6L2bFsaOzNEJu1nAc4vTfXaJnzhNAjh4hi3yBHOQLOpMchK0dKtwgI6qdv169S
0Glvwl2+2WmSQwekv/JX92wUlQE4CidnwWVg8ZVwjdTtGGTJ+9wEnnnScik4S6sQf9ajWUi27dM+
KT89btiWg+GIH7R2ScQRB8EeBLMM0STbgHcY/d5rISibDOS+RcdYQOxPGhbYUrfHbsdMjW+edc+6
EKgTkmBIZsIefm8Yp+pkpdj0WUQiK36007U6Lqc7mdsLbkRzgRdakXBpxZyGSLEy1py9C+c+5zOw
80UioW1cLqxA7IyJtX8x0abUMFlo/TZr5BKp/YmyeUF2aG4UNdTrZXST0IEn6fCA9GaEDtjXZ7Sb
1loVmhESgJMtJIGaesQ33hEkBM8ozSrN+jR1hQ0O9liqI6Q/khAqCgvYeZqf410Q/zcnyCctDyXp
MrVjBAcP6QaWRAlFPeBSpKMuOOtxW6D5QjcBbGz6iMqaEAgjh0UCF8yr7dTnRxfm5eUQL7acJ6xP
DPnbcND2VBsULNHA2dB0Nc+73INo8wxKehBuHkCYSsag9YJxWHXy4Sz/KoeNHkz2b9FH/YpWxNG3
qI5Umc3+49+sR0EZ6pZ6P4rKCkfGk7I43GXCqLCCSpMcPOUBHj2WdRBoNCIbXwxqzSQ6KU4FLzam
XR9EC6Yxz2vUULg2fnraEjh07lsYHK0mxKdMo4i+7zvzipIM75z4SXFIvhtlSTZL12C2qsGuYVmc
WpoQttsFpHMtRUPzp9wKCo4Y4JAMcKE8uQKhoqVGRcESZOJ7acpXcDrfTpSEYjLiOfZ8Roqs1VCZ
GDkjnScZqAsFEqPfXR4nWVxXvNoKctt+JHzk0KA1AKqsQSX+6YoaRsMKV64SZ9QaJ7K0Spo8IV4k
QYKbtzZVL7FlbiMo7PuTRQDX/xuvAoQMf/u9cSSmirLP/UBvyjdbAQWbm9yztZvSbpV6Gs9qpKNk
6hWWNtu5FT1FOGUn9zKxTUnK0g0Eqt5Dzu3FsQ1sVu1gjV0nxLn4po/KjOb0BtbR31qphByqVGFD
VwJg3cdhNXR9LpB2nMROWaJTs4AhzcFsckCziiHZ3NYgzmFBzyEAi+T67dGxWbQ3mDlC+Au93kWa
Ai4uXStvUrGBLdJmWjVvo4gPXIdcHwgzDDFRNDMEja+xflbm/SEuNBCARmpZB0QPbmLbVc7xraRN
GSHlMKG5aQZPWEMuJhAd/VU8O1w6nyJB/e6y9LZuzjffvlAF6rOmrHEOU8aBowGpt/I8BiTUTQVn
SJjTHz4MX65btgY3flEJSs2wHs+SW5dDBE9LXSW4Am2nN68nRiiA+c6lKPgSnQkXM+jPpvJ3kCic
NJB9DXWp+cc+E2mvCXkZJepitBHIj4/0ocbmIOEg4ZES+LQ2YoG9e+yg3LPMV2Gg+V0gMAGSvPFg
Z2qmIVaL6VPDFpw7NQXQ7zGTsmWC0vnRky30/1Ppsn1X4r/W9n95ZTXBa9UVidQjZfgk+Itgtqdq
AqO8CRUXRBaJj+KpbxWPIFVIKiY7PrDyPyTvnDmWymdJdJO71jji36lRil5n1yYEfQJXMc2IZ2fV
g98gZPVGn+fcxLOl/sp57tOZUTzcZ9AQ5LEJ1rUjOrnt0z9YUbBehm0hECDqLFdbjWSjgRv73/oO
xSFpZXKEwx0iciYvgFhqfhDQcGqU6WkhMHADS1dXXCPxJr8Oh84hr8Q1SFnn9g9H4GXso1UJ0my2
FvovEdRYvL141NXtCXV+7F85C3KyxwXmqIzE0Zl0ea1UEjODESsbzbIiyL5jL/6+1mNdAHs3t1IC
o63VfKMOkCUf6Dwqfqf1te2phPacPT7hOwOc8emaKrStRXqz6A27VyJsPKbYIZGNXhujIEF+MKnp
UY55l0YccDdsjzdIOtq7gVWeZDsFZaxELxazeObvWIR2m77aSTGZXQjehaG+FmF5qtMVNpo7V6VC
oBFaF7y/Mx30VvKF4BCunJgf0+dICdCW4MNf2v7hL13sW4ftivGmnvb3Q4gH1jacqs2F3ZO5wDXa
qZCZJxEXdTvKuyIoHoyY/Ut5Kxnzhtzw8FgIMOBCsbCAk1/oInnoCbEPYL6ldx3vaSU7D4XGOwYq
tPD5hpPWTWaKXKr71VyfqAOKX811t/hnG5vCZnAY3Jb2WC96MAoTHkhM6yzlrk88/dcJ6QoRt1xc
nx76ArSVq1g2s4wRjJ/4ZzekGTdlU6uvfmeHu8/f9YK/D2WNyRP8lWEiQvXUpxixsJyL/b+LfoVB
oy7v5vUCZTwyVag+cR5e2KEtkC030V+8P162phR6PWh4xjNrG2owjX0+MjlIvgDGU2dg/OrFLla+
rnmTl+qrC7SQ7KiFx+18g+8Kyxb6dKU5z54cB3q6fTDeRX7zoZByXkXuIzFSUgAa6YLzaWwnlk9v
eZyCOpDAkMFI8gzX2zApr0CQ53vTj+tGrEzN120j6SPBiB6we6A8HRbyEnoS/mv3NY/fIcNUrcB+
j7pLBlolInFUW4xO6j3hq0pdf68odOxJrHvGQ17pKL/jp6KvbIqnFCprr7bv85mrwTRPx92m9GOi
8QpxykfvEYwhe6z+ImCrFN42n5SMuH4/7yrhjaXtLbjpFOtE6D20N3K7TTXWo09RuVmn3LgeR7J9
Ymd2GY3xYIK0CYxGP+EZLXmiU8InH8pZXUoT/I5ESODeWa7AWYR2fwRq8C7EfJDu3dEzpeG9uavy
mkvgIORaA35Turr/Ca+32XsILPDBOYlmZC8c9nTQ+DqTU70h5Wy3yu+NOChDFcK/w+ueSvdrgstD
xBPyyvR1E2FhsUbv4L6SKZ7vBs3vWoE/g74Pw4R/VTrNxWvLWLBu74ALP3LkasxAHag6RL2TGp0A
zuSUg+1UD0p90d/1NVv1PpcpZqW9/QumVFpKwN6RMEnW9k8+Bs/re9Ocys8XmLSX6dvjE5/1kLxi
LvsYga9y6fB2AU2RIGIChxgHYAWdLonX13zSr+cm01K47yJUK8NXBj3GwWA6l/JI08XSZ3N/06Nl
xdCkecpMy8jZB12QSJpLAva0TYGGYdJeTMvYXeZijYMKBm/DP3fOJsOBXvY5nsOftF93LcAKoZKm
I3lTYJAw1fY0riRj9OwJI4LgV6SQ9Hh+aC3pi9PixEZwFTmhdjBFKfp8joZJ1mw6+/0ojlWlDZEg
DAAtY1T1CdgK0RYw0UM7V9/kmDVCVX3YLxvVcmBpcI+P6UiKHN8OPy2Hbb6bmz0h54oFSuc72q35
ntaW0lmVfuk4MjHvk0I0tyddmKWWKoM3Xj5ekdtNJTmjixxPwoqsa9mK2OnXctF8Bzhz7uH37FgI
r6El0Y2P3Onumccle417kgqXIqXSn2885g4Vfnl7kqRIRjA27hzLgEQoIwNB+IpF3iAeJVRwGPw9
90owQpCwj8FKna2KCC52UuE3kNBmTTQSaH2SkIq23rBFWwZSTfjReEAs02mj0XkyxmUflIx6foDy
yiF+uv12VgRQuqlK92qAWKqsTomxUWfBD2q7OwllYeSnh6pK0iVGQxSDLmyF0yDfnt/qvnimyu4s
dxzTqEquAVHtEMjD29FwZ9+PWerd889md2O0pDYgQULpjAWQUogQZOaovlZk8E7GheSFyUnRixfb
cjvEwp/Nq1y//6cA4wuV5AyPYB8oN+vc05qRxeV4xdDkUewjSoXnzG+uH2sDzHmOaUpwkPIzcjws
V8LqK9yJ3eRIN4uBOAdvtLqWp9/zEiHV1zuhSK9V2j2irfyXNfVK4vr654G1kd/Jg+1qQCUZHti+
OEwttZ22fPHU1DFgppdVd13O2WoVNp7si4eBz172hBB9Jolpa5u+6JOoJNTNrVTLVbo7dCYTa+8X
M7wCvuwKFLPJKW1nhZ8wKtKEJc1VtQK+DL2nOHyiZZovSdek3yuAmmPsDlZBTvCyE13OZp/gYK+J
+03tx6uvTtfviHdCFo02dPPX3DRdYJzhhoHuqwtc+K9Y/ivTu+0cnllX0JmIhR3T4iEYPb7MCpBr
cr2LJD0epxT/I3toxc5wrT6D9ELfYqGYN1OxjkQpEEq4P8vuf2ZRO2fcZOirOARD9CGBkRqO6SMi
Y6eI29wej0owGP2yEypucMxKRxxNayYtgUvSMGmG3+tdcTGXl4m/RsA67BH7ZjQLAnjsPsqBYp+E
XMAQ1ERPTTOlrFExIL8PiX5dC0JwkofXwBsIBFwS+9ftmvgyM9sfFKdUpwaLjmI9s4dAPnP0cB7+
6TAjDoPkOBG9yD27xXocSmwD3gZhGnGbHHYiFUfeSx/2ftJfPxMNgWsOpRv0OvxLYLP2T0eZbSbd
V3yoLPe5vpydwe32zSWfNShlGSKWPy+jV7mnFhhuWJmI17xMpk/+x+SjU350lQjiC9bGL4hXlYGv
I5ltHxiZqE1TbVEpa5wQejZkQPc4IuZwyIXl1wVrMSXDEIimdekG1m0ATq9XVUqBP1py3en0J2JE
mpNu3+aHX5qCwRPaqGJ9GzbHr0qFQY9N5iAwvy4DC57bEeGPHw6J2YlYydiIwggkDC3WMm3CMHsd
v+1/7dV4ioXWfV+eO4+9Y9fLeYt9IYYvVxAHGYCpyM5cJNatQlYWiBKY7Q3xyKGX1R7W/If80MwO
IRRYSFTHW2Ay3PkBVHWeArm/Fn0uVhO0msGJJvsfSXlkz+K0tnkX2CbBKNhUuHnJsrlh6TInsZVf
k84FatcKLvd610Z67ISQdqun8lf3lByoEUEkDThiEqKFCRl5wU1TcF4ePviM1css37hz5fIgJWIZ
Zt+NBQ3NRwjQpEQ7CjzhJ1IMK2KzK/julxzCpjrIWNpNuhJYtbcghE8kUGNQou45b7hKPjGk+kbV
XSKyv8kFbAZB2s514JAnIKWz7syV6b7H0/8U9Qn+tdMPQnXKsw3JxZO7I7OrpX55/+GQfdmYslWr
5abzsWknKZgoLv1bt51R0TmF+lPmSO/yHwI4Kklh0jAtA0d78yA1gTWAYmsRRqIAXncs5QBleUL5
W0zusCBjdmKH6Dcb+JL2CAiaieonGQVdlyEaPKpfrELgsWJ0Idm3rWZBT9oEgj5j87JePeTJf6lZ
bYog6urODQgV0oIxmnOC7Ndh+B2lvsf/HQgsg3/xV0gDdaRoTidNDXL5EPQPpdnxYcQlbb8Hoz/f
85sfQBLLEi8cfY+rk5/dlIzQx9bMfYhO8EXWexAfRsze8pgLaxwy0egGfysKSt7vAI2Esrhp6orx
uam8u8qFWSUj4QiIl36kdlyB3jUQnYMRkOA+G2pfmS+tNIv7dwoGOfgY9gU+rzHJM//zyC+UZZCV
P8l10GE7vE0KQM69BqrBEjqqHNPFHAofxIXqfiB9sG3RM1r7mB4iafEQeZ5AJJZjXecQtZK21bud
2HHsA7Dzw7LkxUheJBfAm5QpS7VeSvfEfYhsn/ZeYAp6zsaJXAcVd46TT2fR+2am1NbxOuVUG2s/
rPlDKNOzklbVrA4Av1RbIUXgerR/8JBFP1i/Eejky4glHDHHgFs86X6FEBBj2ZWasuPMVCU1BW+G
Xogx6qQ2gDZfdYJfvS63edUvNbhykOS1bpb/eEWpASVHyebHIIkm8IuTsnjDrbcEXboNJqs2GDpM
wbRWZzupwaOhYkyLo7MZquJ7co4+PgtiPXPMvqMlU63YTknrpd+qRnO0zsHS8/3hK48hoUbaKOFe
PziQcScbgqshrBQNlvEYMs/kIli3nIAslJXzirz2CyBJw27QkgZpthXh1MuIDFq0IxXxvOUHHYNp
ohOdyl6IfX4ST0cHgTvtmP0JZMGHIj/XQZHGVYnfKhF+CLrFUXK+iV8KuXI+iIrjwVWx4D+Zg1nT
fAg5w7IT7ZDCZbxYMW+5SO0EN0xUgsWypkO+WPDEd7Pr1FzowBT9dtYHMWf1QHGF6rE1W2jqwCVk
22Qc0JHpTVRO1aDzLpJeafoyOIDWMJcz9wHzJPbMQfVyIynfgcKozXyS00lr2F6WWocUGcUKmaUK
Fc1R1EdgidjUu4Y29BCWZoTnjUx5YW8lQZOdAO4ggsS3RiKptiS7vhRBg1dkvn+YtIYApqyboTxu
Tp3fdI5Gf/VJWGZDbjoLreQHCJ4F7+2HgqDmrk0ndLLxXcrCiUjXebVexbgaIRtz+tmYfYCfmBit
FgQdNnhot3luyQcoRis+rah4k+RBM+Q36FkT9G2OBJQdJ5B8urada06Nn44opoJwvGPoZXGlYV9+
aWD4zNIs9Wnk4LpD7+pYHhBmo44pCXGZ5cpwhSXJCOy+M/VWjKkpdqBOsSwtSpPf0xkdsfiHImgr
xGjVHC6WdCl0tU1vBspfoxxqU4rbHsKO6J6IokrRNb4+zg8LAJZ5iML31D91c+gjDJ+MscpycVmM
1on035VJLr4IxQk1hjiXbInBPgbBMgCqWE8w8t/z+LT/lVP5pvwYNEF8CIEycINDNUpWkSX+apnJ
nFwaTVrYi1LfPxz86QddcIbwaAO8Jcq758X4uLbC78el/oT+ypj4UbQhMHoE5SyAZeVjYp30oHrV
b/ger0aWvMmkxKqsEOssCpcKQbLv3UdMdTi+vCJFaplBg9hdDbToRuDzarIJRO1FjvosqjvXFRJr
ufb602MxxivheZ8zTZ5yZx2nkc53rGIIV1MiwHX8iHlY4aK22GUYh14ZE8o3NZgqmA369pWe1aJa
AVNl3XpO+JS5kE/Y8AlPq9PFQYwpluUm1X7Nb67Flz9+D+gN8h7IvwxwIbbtB4H0Kz2Mi30cUY1L
g6uFG1/VD7wyhxwHcDikC1gyHWEW1KuGtZdeEYVq/tJyJ5VLXJH68Hj3jYjBvK7vLxHYZplFsqvg
jM29TftlrsvNhXv+bmiOOd5mjGf0HW6V5T/UC9tbwjepoEK/ImAHm+SG5T/YNfXA5vVj1YstmH+g
uGe0ica8emG4PdJ+5y+WBmXJiFik1powUUQ/IRVFLTOP4tj3qEezxq2koMNHRutIn0WWCZNgkUKD
yU5Wcg7Ska9Y2K4B3dIIM4T86Yo94/+KdFSg8VuTiWVoi/deV4CiTDBbRmV2phCXoQLwsR0VFOq7
Wq1zw/Fq3iaYUdWxOpQHDOBlLl0fjiJsJ5oOEm7+QzttZAgty6XahUlTHfO/1gHlOlfk5ieXjPrY
ejEfBoG7V8LSfFAssFrxo43dVgckpg4iJxQUlxooa4vukJfoA8YaarjDZj0W3Dc+H4hbhb9e2yHa
wTGEgKPSHXN4yYybH0qXMb2qK7jKCztdxnKquD7rgjTTWBTOBKFOEkM/QCBttuEdmqZjQQufN7Eq
gh/HZS9hZ1YcI9O7QKWr5XQXBcYncCWwH+PZJfjBnBSWTjkaWUY3ZZc5g4GzMk4zq7pnaQKLE9NF
PvuGltiMDCtHewxuTQ79ydWhzuKLF5W6lfLUPDneH1w5BR84iLT/MhZM8z+IoR209jVFsQeefc6y
1BGGxP7lWrKREp0yZl4ZASk3Z0XOkucnn+Ke/jYmijYFsk9Go++FGDc1LgF8z4eP0Dog34CLoEig
bRmv9QXwaU42/rhvF1XUI7jPGtdr7j6cVvFEB5fQ3ZanpqdjfQyzGrHaaswJeldWjBInNzlOdVeJ
Y/gEjK3IQwpIh/yxedz7GyxSfJ3QBtTbFjL+yjeQTpZEvFwa5H+9IAcZSmunSwR9+XItbxHfSJl9
LCLjP4VYzpBn2snFFgtCATqR1RKJwoAC6YNYsX5oN1mLEwC5OAomMM/WZSQk8Hbk42HV9bdLh0V9
p6UVonDAbY8SrjAkKapVG73HLZacRUqYMvcy4Cl2wLrfj3ror7XS7FBe4RjLrGa2EcLMQJqm/a7i
oACu1jXykd8Bbvzai07mhFmjCk4t/BHTkgkaChuC4EBX+0TdYlLJsMJrd989XVdQ/lFEdcY+XWdv
SpU+UkFgn//D2ddQnZvMwxtOpWcIcKeMwT4GFcNA5YZcg09uffao01bs1IwDhfCF/dgf7QCzN1W5
8B56RxZr6GpPpvYjcbjEvJL9Z9dLe46Q822icp8EoAg3ibYRFtLBlgbq2Sed4I8mEHZvu4SY29U1
oixWWnQ+PXwgMzv7MH/rPS/dcF74pvDWV/zXD4mtSdgbwUq9oX3Ug7NlfmsqP2y2EAuccuvDefPW
ZlbNDUm1pAL41DXnddhQFvKsB1+pxuhMz/mdF4XWnE9oFpsX7SQ1ZB5ndyjeBwiEHhA70pWXnXhA
HYzkc8JgR8pMO+NzmtfOkhoH/+0/3ctD+vQ2aW8re9xkn00CPZsS7mMMRXdV5LlQLtCcUg0CmghK
LnToMxQblP2ixdO2ncShG61gZqmJ4L6Ti08/LzN6iZ76cIswUPcY8dld7tn3IJVzbwDRZRsoAcby
AKcmf2A9mrOPtQqDo35LcXBZAL6qCasmJxDPgl6LsQVyWYaKLXtCnYbbLPD80RPC5e88hzyeHs3u
6E74V8+dJnE81F5CQNyMpJ/YXKio7TmTOTzq0zH4tR7KjVtG84dnMp1ffC3GYyZRz9IA/j1vVKpm
DmpbTLxVh6wUMCGLX/qO5vidRXIOlQf2wNqJ0BiM2d4Tm4JRTXKHgConulf8AbUQmLczuyCS8oid
aGUwS7gdHEEcFbZV25gw240iy3GQ1XyfPKm6vudSn7HR4Dtr1D0jkVpc01EujA+vMtN2EZ4CjZr+
0NKwH47jv/8ha7MI+mts4RbhcaJ786r7tMEFFPy1gnEU+5ASZH4IGwYL0RO6+n1W3HW+XA9BNE3G
V+6bs9rcZscNa/LpRKVel8cgiPqawgIGtpZFzZaUzRv+LobeVPfhU0uL/Wi3ZR3eb/vO/o8sVa4Q
YYgVuW9P3i18Z1hPjE0wIcVErKAOB3/snzkmUbYVBxKbIuDKT6HDIqBR4FE6OpQfq8onS6M7zlXj
LEB6EmdL/mjpdhHS7hCwmEN8QTRoMOBCI8pQye36kRGE7tErYVJGCNfOo/3BSzfWe9Sn+2ZhWx1e
s9IJ1Fiv9FYdf7JhNs1aRb2y8yb9KdaF1VDPa8ROJl6ZACegbX6idYYKcg0x0dhfTnL1eK9YS5wQ
lCLCGx/7eN4iebxS5z+oUkiZDHTd+eGe/zxbSWBnqVy5ZYR+wHutjK8hmHq1pM1PmFV81N01z8iv
eBhOZQm1Oy+9v3znmhRwSdxBPrxEoLzj/WM2ttUv5pGX7Th1RunWEcdkDUFqSyRRyMh1XOmCOu5o
DPIFcc/fiQf7fhHCZtV8f2kvxc0s+ch2ylTeWvcLY1T9phterQOQMGO5MZ0+l4cRfedBkE4OdN6j
7ux0hE23/ZIY+kTD/dZC59rzEg3adCWZjEGgBj8/hS7/iowIz6R5eOB75nKjBWiHQv0Cqc5c65OI
gpXapZvSmdXA8TaHHZHFgq1RvwZ/bTr+IhQlmxpAc5u7GyOwupMKKjo34ATFdfuMncYmtSYwvQCW
rNwvHH5V9oU6gBq8f2O8eAnUOt8xtdlcdrDCHjIVx7iy9+yZJ4jAv69m74WoCYCn+4txFXdjx222
ZoEv8t08/dewAL40uxh9IkWsl+FOyZXULqn2m06Qh96eUalkLlUtjtmTwAEkvUloWAMUeBhpAKup
Z6W+TA0dk2GGOY7n928m7Eoe4Oq+RsSsEYrX8VQFs7NRDCT3018QtfFO4fyWfFskBr5GbdDRTp4F
2YOIOlQlsRuS63BbwU65mhJty8TotVO4BymXKuPmRu566KBlpZsFKvncr9M8pGhUcjGV+sFOcPSc
4eJpSuOY70LNw51Lxi2oefygnnbF8SgQO+tFavphsl6RaI1QD3wa5ioipwz4nWBo3XEVZHvVHo3n
M0U/+WQg0P+5ypflPiCZ3nFL2WsTqP5p+ScTQ0w1JPcPvkEbV39toefI64QEP+CwPOn8Auj+lPtX
JdxLLQH1nmdOLqwKEunUP5j5ree3E7AJNQ8oaIrReRXeOr/8wX36lXMXmaA99I2CSlYgDhtkK77b
td/S8GKNQ5vn6fxOJspKqFePbcgkdZu1plffdyOw9yIyW35fUvMTv0yxsdgCclfjTYc6IZpss7x6
yizBxdRcDxMqTqQSUE20Q6KKFHl2VAujpmiJFm9ZeROdQiu83eTX5iwXn+w7UKckapoA25/OvBFo
2d7FMuuFNA/3X1Cl59/tevyJN+0uLHeG7hX0MfWukYKntH1iP5gd9EQA10Xa+8ezUnjfESpOX4w9
4zklC2UqkdsAD4qAUU3x57C8V+1JbfCrRdk2v/n8RcCjSFYMzu0yZDsX66dNWweSpAMTz+XDzBWb
OvFGi8jh/bDoixEURxbDnVtiF/+Omq7eZxgVGo94UQDCNAwuZA+3AXisMBNLoHVOcL7oWiKEpNnn
8TzGWoQjib6Z8iAHkcKQKKbHkCFt5eWjXgVhVqmd9KO9lU8sS5PH6mDzl2/dOcvtKoGzf4jxvqrT
sdgbNrTYPjKCdCTVnaE50dhyntKZz/vgApJDDZYpPwZflCsCPQuLX/dDGA6nEaOQk+uLBqKF+O8o
gQ+8HzRX7mmgh6GJLMFoPmOMk0Fau3h/TDSvHtPE4Ex+f/asRVPWG9+6SRCq4HoMRdUQY1egKuCL
bFlgqOgK109KkVFOWhU4qK1dN9M40C9hSPjM4UB/ctLKKFFPdN10u4pHRqVbpgIo6pd8vGi4qMzL
A1TV8HyYCcI5OmoG2NIzYyDV2x/5laB1112vIRwoSh0sanV6kG9d86WQsOwCodEvMB+JlVogFisu
euSJdH6exRyLaeLQxiIeh1zfiTi3w7T1HtnnfvooplVFHF/Z/hGM1aZ7H/fC8ahrKRnTU2k51AKq
Ge/78daq2fXVyPi1Zehb+uN434rxytMvrDrYZ6Lh5fl8zrx7b+yAfby3xvmfIa72yV9p4h7XGJeu
0R3FUEx2HhxuV71CLd1mE9n0z55jsPelJEe36ESCTM7Wq3V0wswWis+IisXpbdWo4fJ29gMBt8NB
iGtuaEveQQ5672VaO2dZoUqNmBgPKRbol7YkhZot4A0oK0HzGSp5uAafaLAs+EbK9iXw/ITK4M5R
rH87OesvtzEJn9EbVrRqNVWoCLVM4ucXeNRgddQXrDIBQ17Ent89DSOGzgYITPTxId5MHHMGy17e
9Ikw9N8HldFFi3vr/dIkRfn7uO4I9hhu2c2IizRlk0obdT0tqGuLbyeccejt3WNyY5vj5HN2r0Az
knpdT51Aw9IhR6rAjRkT1d3eMZPwN2C1v1e8uPj6K/kMwwCrhn7rHLwlafbKi+NdaIKi+T1lvCMo
5hpiRaTRHqeRwzSZCYJXcaqmOqtDFEFR1IHMjVb0hQPz0jb0L13Y1fcGUDjy9fo9UOlPHhG9F7dU
cTbkwOs7/n/DLDlg+JnYEm5NrxzNIkX5QrQXgSXLLXibKu4mnsVLh2q9X5l/sYHHd2Hh636HCDVF
rUg7kRXU/4cjlTna3szBO0yOXnfA7eQS1Bol001W7IJ8GU2WzxpaA6quHAiD+HY7t2GV+pLOYr9y
78jTg58gyGbnJ8Ttw2Ga0gbnNS25W6uyKVVU9Ct+CrQ0hpOnW+mgiO01p8742cVhbG9HyM81uXXD
juwKs5JmAp7NywkoROGdlxcPqm0PAR81fdB83rICfm6qDeT04JNKxGLnqcPe+ejtLa4fxIMB6F/W
yg/pdHuch350h3z3hvOrPA/T3RSIYBXv7/VH294Alpi9PjVOZu9JHZncWWV1riRg8Bw3YyStCAF/
xX5amM7WWEJUl4aNWbe8tQ9yBum2xVAd/v7armytJLJgGUDINB5drL2DiTUZdazpX8xelN4uuRV2
2Eu7qPMNROO6uM+dYmqdCPNdWDnLfFQ9hdA/DgiqcOgZPEOVRc+ak0OW3s447X7nGdt+2y4oP+/X
5LX7Xk/vmBSxSGRigi6cNjhpfT3/+sJMeDwbIfFI4CRQtQPqRk0GoJwe5FhvvqckFPTmbemmX3wu
B54/QdgaaK5lc5u8qFYstKbJl1d02ZZCn44kf5xeSdHVyplARWaYHPO7diQM22OekA9CM3Eu79Cp
+Xjg6QyTt0icarAROo0+qJhOZMsSaLfdYKhNIqF8xSNApuqWm0myIon9ER1ZT8genHcuAG/Gqe9Z
frhKwVsg5Lw0mITmkzJ3Obadz1rIhrrT9BtgzJgsX7/lBpsVEew7zEeji60Ybh23d/j68eHKj4SZ
jmMNbHfZzugDztErmduRFubbNHuAM7Se1AZVoJyaIW1nmpqQxU+lnB3FCmzc+fFIVB+J9ASvMcf8
AynbqYYxr7ZTxwtkiphxmUOCO1XBddfscAi2Ac+YFqP6WUfrwEqwAumGEeiY+/zL9NwoWNbt84b4
Hxe/RHQiYFKevd3jUPHwB9HZ2QWlYeBVHxen2F9GlcvLa4mNgsl5Lv6D2Usi9mmLZ6bWG9bw5Ma9
hI+dG3dvm6Ztf91uZ6bhNXW8CEB61j1LRj88r1tCClWKfmrcD7XdwEG+5tNfWkMDb3GmUOTD+MdB
YaqfiScYBGvWs3a/7GgjJh8eZYj47tYx0AxyJ0AZvYgQXaft1bdTtHVNuI8d7hIm6Vh5tc8rPTOc
tBWjvTVbqxLHXdiJ72/EkqvEANDWARYfu/7zApQ2rOLyUDp5+6cZjsjp8bl2+9PhSp737JcSr4ir
pPpAb6bpCgpDCma6K5BtBcjRbBgt8dmhXV3+5tE1vy3tyilLzE7innSL13ojeRT3sqPtzwiZcm4g
YLN1/JlZSnRp64unrZZorIIJig1WFdGAc5K1BY6brV+DIbLTT2GkrJtBzN2/2k97QBFw1nIvUi7y
6duxfc3ruFfYdGFJ16AVvJxTf+MA/PDOcVbAFKqoohZ4z2ZWLv9KXoZ58KmlcIT8jsjFodNj8VDT
w9XfebGE3Wog/qP4zIi3ZujK6HCdM3bXiMgJqRVG2ViSreNvHN2QWy23Tgrll7qx+POalLhw0YpW
aho7h9xnwYTlYe2YOzgjHXpUopJaD3x8bls7jAwNeEA6fWHUUVY+6NeN07/sMhwBvEdnqd20AjxD
HBmvykawGfburJR2gPLvh+7XewKwUNToiCtkai8Oggn8/SBhYloYPVYQVV4Rx6x9lka9oPxNnBpL
3zerH9jabIwuTChAJIfG2/f7gTjL9IM0LGecxvbA/4bWrVHMnuGI5ue94GomProeqWzsNm2lUteT
8YboQRTcr1/pR9HsrWSkd+S9sHXKzT9RFntfuov91M+fxLS+N1y3LWXkGAYgSKskgZxYga7pbCeK
EFyYNi5AQ8vwI+I38ReRkWAC/ovq2kpxVd5vtWleF0lS51uTOhJrBsak0zrDsg2NoRgmCek4WJK7
Y5XhbQk+tW/ikUadCK1YCHSfHHrLnNFCMW9CnbOkBrQucIep0TTwQO6MB7uijmNO3LxTzp/9Oq3h
Ph9xYIjJaMsw1595ZLs7siwtvhzRVfkiV0r5slakBWlsutQh8e0AxXIwxziTdeAY6WFrctWbPA5T
sw+2gEFGLWSZ0VNVbmxdhcnuRl5IgocDCTbsptMntspJPqcLtjpA4/tXpcPRcTob8q4hTdv0sdYS
QqeQbfOqrSTfRv8w5MILoPqXRjT2fuBwpuN5trqrWEtvwomontX0hvFJRmn6Y3/iUjHoSFN45Vng
e0yFSFF/W8V75Uc1sX6bCjFyyRKl43hJmw2vepArWRRuuzVRKSFV4crlpbl1LNgsFm03vR1ZaYtI
RxW6ehxEIFHZGegpExJlyG+H65N/aNcCK95wRtnfLWPC5IK6528z2CIJYa8UEYOAjdgeV44HTDT4
72qofeM+b9fyBZOPtnMB+a5Kg9485I9TFl7Mnl+T9BX9NfgdG62uibKjnB2IP+kgzGxxoA8O/ZMT
K6t4JfpoD8mYKz3EjpeUbPa92NjOAcBNYjGCWNJV51u0dcch8qYlIzKAC0bJCxR1pFY1/zmWe3rF
nowc2Sf3JwyQm4RkkZXB7lrDVw5Vje7a19W+CV/XIReOZYSLMVj15/4h0xZqYJ2c66rxYcbFKHcj
Xw25SSY9AdQNzM7VVZm8Mn2fpNA0/ZFtjr57Ve5yA/WyPS+NAQgwNvkltSNxbnjMqBxWAIp2seN3
Fd1D606t/enokSs6NG7NXuW63oxFJ5ch711AYV7lxtNolupGItPvXuzwDr9/B6IpP//JmuVQQBsG
HeVcPq5JI50IF+qhvsQrwe2qIimTCPhbDQndFkzaPHOL1n7HX+mquYkpHkb1DROMaXEJjZt55Fmr
pxP6cZyFp6ZOHhk71wJxsFX4nWIiX5pAt28HQzDzi7h4FsxGJCiU+OnIjWYykzcSPx9wxGoftBxL
XnDWergG7KjUTG3qYfJkWLq6PLcsL5hp+kvs/dKqdIrKBVqFqrf7BhhC103Sv+utXHLi6M4VCO9g
lW3+cepYhp5kdtzWTt7W4EVQnKjUbHyWkS88baCpgLw/Ss67/jlIBWSd5rQbJWeote1tWeBtKv2m
Q8j6xpmaLOkFXGERotyJsPpIxrgTJBIxxa6VI8JfzeV6xD/b/e0oSDl0VxSap4RJHPASTV2g+mDN
fW5dS0troKX1juImMVEww4pnLsElUObWDD7KlMrKQFB5mv2DggU2kpbHiiAUuBtC9Av6N2JDUA7B
qkaRTmN3uXsufU+vszriVOKunA6fo9VHqB2LtNvr2Xn4R4BJohopnXoZTgozdSBtcbOiBOuwKmW+
Kv88TpnGjV36kWsCEbyv5i0pC2ZL+Wp9w7TGtD0MlessOsXiu9R3sSDqXpf5VUYUeYfT4/7b/MmK
x1AVYsRw2ZbNDYIy4vID8yTzI5MI0ohT2PxTn4jrxwOGjJcwH42j8JZ4Wq99XUW5h4oKQTkpYBmO
yeqPOR12Nk6fHlGM9ITs7EgnmTTfrEWnJgg305uTiWVbdKoUBwHMJp0ueC2jwbTlUSHFMAgylP+H
gYCDiy1FhSxKqDgKQjgc9ICehutolSbpVYftwLcyMS/nY+3xqwdx2NGU3JujQA8ppqEVkeJPSMm3
m+taB6n0fN0d17OzAbWCgMYZHANAkAhc2t7avx9r94ev8N0hS9AGpyy9QvXxeG8vw6ckhuBck4XJ
Khj6kLg3lCObKmxJ4tb60DX0TDNwrVTegUan1WB/Y1JCY0lWEnJsigytg7CppSkjgA2f/2+6OBFv
iHvW5kSlUYOISYYRmQs9Gbhwzh7sJgF0lfpVG5rOQqDciOQvtlvbLm1ysRnklWdjMMOJz+X4H0jx
vZwu2JRrxxLY1LKCKJ8+5dgX6NScSV3cCW+7RhqQDd3sAfQKpYygCSr70dsnWvlwU9k/7iAunPpu
473PdBinI/JC0V3lIlkWzV8lqKpUU2KO53QmU3X2xLorSNytYhu3VE4C8/ecGxGM0ZiaydszA64G
z9goA4tJw5k3ndHBdqCfGuO7tpm72TqZhvgh/Kk1CHhk3hbbtoZ+PGWTCnAjF2sBZcGB4RLu3ttx
K7Eagecz57N7yKnn9dv6C9p2gZhFYFIVw7NmLm+SuGUhLF56J8DddbA06mS5qdDM3hoju8NtL7Yl
1RgatIm2b72CFJwskwTQ5bGYv5Gbfop6GKSGdOeJqk1siXVVFslBM816aH6djn0lAAtnN5rfPFwk
k5NSatgN4uePzpNJLxcyBj1zX23ayN4PVtYIoxoMzoG45fXBqAnpdIJxc73ls4OKMeGeKGjIIsPn
IHp4VMzrmhK5I+UBbGhiVDCSejwKX+Q8ORgWLP4BT0h994JtfQQUEamZhUFxN4Ipbjd3H8GWJk3m
QSlOfSUqXGsjA+jU2jTj0EFjE2Spisq2pR3S/FQDubljBso6OP3JPwRmjU2vCwZtUlYmmYexAFCf
Azr+NLg1ZQsR2ugkQ8sa8Uh3by4bknFw3IZv7/sRmoanVCK1LLrjJeOzAbQVZSiWbY29+z5XxnQG
g5fVfu7yAsIEL+EkCuwOOBKLWjlKrVid7F2Ogi7OqddRm2mdy1LJLtgLz04BIC4ndNwVKlkR8pSf
xFa4b6Ohyf+fIpm+SE9/DYe3TEijCmihZwTPOY8Zm84s3Se2qX7b/2TICT1h9puNzeo35vilXYw9
m7p6ucCSoKwslON1KjvbcBusJVgJvC9ZZzZwxQrnUKnr9FX+8QrmihhcGOtOwcyY60AkeGMXwsC8
g67yuRDDPRX2gMrM7E2RnQPoj1d9mhHkhZVWjqxWwwCmZ1E/AWO7iqA9CtSPbqXwNWOnfFKurHoC
6Ic25IsF6+16xrgreGmPA6wTKYiOoGXzsMrEPrQ5v32tC+hMeFQlrF1Rs07Cmfq1Wis8Ndi91wbx
IJhWeQwn9hJqeTCK9dENQfiChRthphiHzK8yrbPlZcGfI2rUp1VDMJyJTW2oyWHBs3BiqamoKf/e
cKjRXXdd46BPatOemAC3RoMdghDJp3TdIr/JGqgjsLN4AQOkaa8qXVqNaHRFgINndW/hhZ3QaCyC
OM8AyB8FbhR0nYh4xalJm3DUVGfhsGQSsBhXwS1YFPlcX+1SX3bWngaaH31m3Yjc2v2KlG9jiGxo
Uvw19WeW2TRVk2SZKU4MJxQaviIZr+UY2g9ErRLxycibVwsHZV3hpfPT3Fn+glGGpY3VZDYESp7f
0g9ugpcaVt5qXx+/rYXmGFMO6+SC2w9kBhZfjAjvvE1KQt1JhEirUWHz2CNDl7+S8gdHiy5MN1Jj
/ZvlC4TOiiDkD0MRZ1adLDyGPMRQxsWUTOO+hSo6IKTDK8mSMVQafAZTRJFeldJtjdHCA0zAk2dF
XUzygYqRgR2RqgZfrITFF6TFYV5uoDv3Zeq4WYrYISCcoCKBbPJh/O0vLWnI8RgyvJkKEDmZjseJ
ED97TDji+4+uQQdPxYpllN4ElcZ+WLNNwvdKQ56Sea3oZ66AGVbhTABHAzsU6yq3yY6VTQIVBsJ4
5tTAqQnIDzG5gQow5J+svD0OkRiaz4XJiyxFLzh8e/9IRUpbn/VTfvY04SzSyJWWmKQUzb1NO3gR
LvMYCGoRi9b4hEi4vMVeuLC5iK3IQpebPk0bnvt9hGsKV6HB36kSZ+V/NtQtb4TsNx8SWW0725wf
4F2uzPr6/hP2EH8603yAY5WDxGATSZOtqnwEhlURLkSNCwA+OTet5AMEoXYIz0updXy13wFVvwYS
rya9SdoUKjUFE9oMVLXcPIcButabOn3CTJmsu/otpmbKSe0WrYHypblIc/+4dD8i2LfW2d6HqHSi
Oe34hFBUg4sDqnm07f+oWYMCU2S6ac9fMDImCUuFeF1Q2VYFNGmAoJj+qKtUB/9lHNNteODmq5lH
RsyUH8clmWozQdGqHLMZDrXrAfGNsNtyjuOT/8/3UgmldVHwvyIpVPJpDkzBTZuMLNBK/HWwTzP5
1WeN0XHjxdRR2bfm86g8uoMipT6rTtIIVUEY5L6r6oLHEaN5ZP8gzxTlHno0k5YbBE6n2WO7U5qc
uWKyMQIsSX2qfn/lcrjvOPgr3bobJfP6CId6x1qFP3Aj90/eW4pXorb765CzX1N//gdVQNr6qJ8O
NL9/NFEo/nABQTnNLq3EDkeRTS1B4HUNbgp2LO7/QqVIngGxYjo320+N6sFm1xoPwC1Uv0h5iY6s
lJR/y1rueBAHGcnw1Ud0ayrpGweJaZNHCpumV6Nw/q1idLHjozKe19ET+Mw4IhQ6umi68BVRVnnD
OEMOJ6MpStTYAdaDgp2Yw6H70WleZ2dSUgRpYBbvm8/cw+Op0FYQ8Oed0OiuUeM/vbH99tUXtfTt
HeUfVIillgo/Bk9kqrw9XSeQsJu3ITU2Ro8r0dkuk5t9hPIpDd2EqhKqQywPp/UJk4mxgHqsAunv
G1cQucd6Z/Xgnn1rrbFGVMrPfF8sFiLL3iSDzo45i5IiLublR1zSZcrsFKirIrVG/zwtiM1d4IZ3
Yk3POvll3Avw1lQGCRnRsEjO+4xZgI1mzsPnAhcRBy5no58kQVyUbixLrEr/HI9i2olL4Q8t9JCP
lVJ5IcMFhx+ZTT8z73UOE0X0mRjk8wzsRbyhMSC6ZDBdYP3rylrTE18vA6e3yDYSUStZzU0FK6g1
R//Qm3j+J7N7U70jtiMl3lrVLK3EwS4VCyjWRoWB+adpO50IbQvTsQfCgLBZchi2l9MXn4lLGAOa
tjOJt9TXG9FroYzChIqBmzU9fWkV679ioLBZNaKadm6ch2Kp02H09ZOIgyJddJCP3ro1BftFjyIk
PDER8ANf9XzLX0hdDM9V1OSSfgUgvA8j96oFPXwIQFQHsvPKVy50N6niT/9iLS+JvCbaP2/Ywy3m
VaqtbTNWWTb1VCmripeinmt5ZyohODwaqgoe6PFfgUljzmyMfqtjY/LfKW0McfvBpg9Ot2r3gScJ
he4pH9ExpyUenBFloXzmF/QnydOwGKoLdGmzysmcVnF8BamPmoYUkK5wr22Vw1Yuh17F31n/gEwN
PDT7iL+xx+bEcMCOus9l0mMUx3s6etisX6nkIfre8GCakeTCox3n6Ek69saBMToigdQGgYrSmmFR
oVn7dK0z6g0kwS3ipV0p5tXoXpvawMJ943F2utyQ2MNrmL05W6BU62QQ0QczykVv5Q7xKbFyQ50/
dR9CLKESbxC0wgM7jdcMNbRLPbCB9U+KgXLFOxOoGtb2Ry3KidFlZPzo9NXomf/quC5xvab3iyMU
m0k6FuSfUoOsDxFlneMgP90lo2l3WI1ZRWUnAreH5KVFAGqdUUxJ3wOb04SrcPLNiSlHtbchDw07
vNexKZW2tSNHpirP11BuxhN6wxCEL7Acj3OHowPtgzx66limwfwMqwtmq36y17byJuRBZ5h74QQB
xJyyZdtYgAY1t5pW/AoMAWjEpTc72TCCB+LscXZYuPoqOiSFO+czAQYzHYVNAj0Wz834Dkmgbzwt
4WMYd5p3FSMWRL4gev2ZoiTX/vqfGCjS+a2c97ErDjdjZ5ul6KrU6ky+DGNYFzTqlrwhmqgE4b18
DUL43tSreVKitDbUCmabgiZ1YsjpTjSG2pM/vqYz2xTQtPMrsd/YE2iIgGVDF0cHvo3jhZRsLDjO
dOXGvzlFwMpTPsq4MG4Mo2EGUawz1HuD66CbJ1usuaTcyH7ONMCtyfNR0P1JzFmf+bqHcVjvc9sP
uV8r2tvnfFQpPWZ9zw0jy7qAIZpLH1AMinItKf6xxHpBkmcfFQorPpEowNBpBimQ9Fg/U0XePKv0
PNb6fhHU75Y5o2RWOHjy0kYmQzFDgR16Kdq0MnAUNviiJFKEmKHyTI+hkiVTsfgAzHT6+u4nU2Ne
yuxXRUw24/lhqQmbvWmg8A7Uyhu2DKhy65zR5PVJRo69zzNJaKLHnxUuRURuWhJrvv2UXUd3cdBf
MKcHC+y6lJYXQBSSgMYLQawKsR6ERFWu8Whej7EcWzbazZkJVuD2yPlCIf53WW5om3IIM94OyqJ2
75SXRYc9twaLGhJstXz5TIrVWRHgFmmxvp+pw31ozEf/71RmRJQnDi5pnxFQN/k7pcNEvXmB1KG+
GDwkteCQ8AQbDQODZ6dRMWbtJItZforAq/r/XpgEG1cCSlOdRp6P8Ipbzn4zVegZkAWr/aJY5KAD
qHpjzF62aximNeyi83fZl9tZVJ13oV8Mswrs6CkLvDQe4msJjxVltJ+rLbzbkLc/IJvtVqLczLOh
DwzaiAoo916+BwovLFa1ei++Sn6g2L4OZ6DcO2XeUZkEF98LeeOWfBJAqRfi3b2BH1Aw2PbC1MId
/m6XifSjP7xiRxeegC3D0y4V5WicMBmRZ1agvMZuSjYDm+bNjHEBjf7OsJQm6T9Bb6gLZE3AK4lk
7ScU+vAPc+H+bCEAAomS9w1lyIuZlxtAj8I3CK9DHxkReECqgiN3w1MkjindgCrursa7c8Q5+58T
MRqeDtJO+L2Leqssj/PEpATipW4VkN8oZcT/D7Lstl5ZF1t6NThZWAfB5q+dPZ+tbu/JpSn3cFSM
lFE8bUQPBmIfW35yHsFgEeU7fF0F2PpmyEv9yjRVWtWULq0dMdnuPBnkTN3tICcqAkM18AMqQeeF
VWRrZ2NexUqcJvdtne+c0O78jpF1H1B+NQ8/cPk1NkSt6HoEvLOUu7jUquAIDPeXVrsL8h6F6Di8
g70o3iYXhARZDUrPqI497xor72QIg2lR94U5naL5s8+7uZR94iDuVKwtz+0VpuNdKXpCtZ0GrjET
p3PshYJHiP+4bg0p2Dpjr1EzUoWaawGOQmNKgCoQwu0I4+wQ3/5nEsM4z1KkDnRxlje70FZiD3Jq
ygvL5rmRDEBCMgLFmIL91yXnRcpyMahRYdl3cEIsXP8lNwyOXNnpMP1YyOvQvZM+ox6mmUau+cit
2V7NIBpy5Fd0/eiYTv/6T0p8COvUNbJnrJGcJ7dysOJ+RaMLn2X7Nn5hw8WUADlrhP0oricdbjd3
fXpJ6tqn98OkZnQOSwyt1sqa02mqqrWDOPycU5aFmO04Rz0PSgGCWXyWjUqzDFtqO+IbaFqI1FS7
R3lwDG395k3EUQG1jDpjJlxEXzsBGR5dMp+U+hXPg11LgxbQQSO3RFEyRqRwRw3po1JhvOLej0SP
PQ68KMD5AMqLsorucuUIFBnIK/b1o0JUjsjYDmvv5z+85gYZgjEv2Ia7Mqd0T7TcZWZ5OAJT9+sl
/invAn+XaVNpbzf89G02UkW1EbrUprQOwihn8gPwzlVXSfroDGvXDq+8bjmat57zZ7GyICat2Rds
6sJujkYu4ZriFTkGZRC0SWAqBtwg5w2Bm3sQOkFQ+i6NeU558t7A6iVn3ACfXMc1MU9kBNXoarrB
QNY2H4P4NfMUgTFT79F3PgATnMmQJbdEG81TBCRfJ8ukLe92qW40HxWYM/lRd5g+kYZQ9DdyLtMq
r46692Yak3kXxoViSZpFdaRJOqQ1fx6E+7FHjVKHfjpdIYgdcqA25ZbEU36W5lnQyTgNxiklfJZ6
7xhazOzCe4KQA1mdQbCEmGBGYeLAzgDvFpHjjPfzULBIb9zMwHXsQEyUsdCD7HxC6hBw3B6akGDV
GrxEbVkZIBZF9E4IV/Ze/8rQz/2mjOcoRb/tNyJb1Sek268SWdam6/cd0AEyolpKP1THmK/F3EiD
GCChAGMtkmRXgOSozCkeMxveU9a+yiruQ/lfWPAZ3+g9P9ObU618NkduPvvzXqbj372uioMiMScr
hmfWjrOFk4yilcH2NcXTYoDN1TwqrAx3T0l1ePuPyiwqNAr8Rh1gCIqM3hzJnGIPFWiOzNDb8VTe
7QLlyBhToQ13M+dXRQa5GImuuITow3qLl5cktjbsiXpnz6Jq8k1hqAyJbGueYfy5J7HiLYZny+sP
Yld6WLLE73jNPwO7J4d9iwo+AQ2ZZIeaIthQlcyC8WidOGv6dlemLR9FRvEhLkfbJnnN8kvKshEW
+iH9UOlmlPZGYRsaGsh/sGyW5daKKNrXtI/QWJVIxR/yzKv58c2g5ZTk4eVD6iL0Yx0QC2vNIWHL
dY1IfpL7N7zCpvkPvxSZu/GrLBAKYqK+x8jBQsXWdS33nA3FmQw4lTeum25HZaEq77K5N5efL3TR
g2S4OkUSt8/pZFEcT5dKtp0Tmc7KxyS8LnYxnkXvGqiMfsZJ0+P9JIpWEYVr0FcgjZMKw53g6R/B
Svm+4sHg61pyCJ23QDsKG36Vo3iYvBB4d1t8nElQcWuduOhhjBxEWliA81C/a4jffkj0CiD5YiZR
egTYysLRjkaOeMN5fXPxwbd7l/M2GFQ8uaAKTmDyCDwyHUdy+1P+ACSQgjd0LuSDbLL84j7Q0/jP
zD9/LwHDR/02slLw1YWAwyIK5y5ZqtHNKIy8GZ+PewHth6hGKjlzUgTrQPl/MVDd1mShjA3Qvl4z
PhUOfD0RLX4pwg16BS9i4gwPgN/U0NZhtP39+EpHmQH6z8k/xWbYSnVfPmiBruJlOrvLIGXkTgMU
wm5Ttb9CrnTNVz0zbbcU7krcDqOdWVTVUcRXx1T5EI5armKNuTPcfv0bN0uqOux/Bbhif5ZrGyQU
bN9dLfV6h/brqZ1/ZakRqZydcWDRKku71GarohdjaaTrGe33ekIdnLSbnHWg0JPdx0JBC1Z40jAR
Ti232YGmm0IUW1YD2xsaXFjzodxahYlxPd6vEAhCJtHNT56MiQgB1NNLueZJNYJnUe8D71NSj7NW
+Klngq7D/aZyDptRCTrvT3aZV2vLUNJM6FUm5M9ZPP0I8ETKbe8NmUWPRFX5dDH24J/U2vUeaE+9
PTSplct7ncyJUI5OUIz8tgcF2/fbRFDu3XCfzUI1sPU5Ce1He8l44UyP/PxqI681aypd1ztk6EA/
YH53DV713Qo1nwlsOhN3IFm1LoAtGLxw8Y90ittkCKl3woPVYiDWda5qTpSnthj/iVhzI3pD8l1F
5JB0bnEFp2xIAYYSRy5CcH7WYqrAFU+1xLqN0FqgnOdqH15gtwv8hvKDlhsNyG0ccRgf7GdG50E1
YQe+p0r2yOKCulPlzaDZBxu6/60f7yZ8qPHHc4QUXrmh4l0ZI1fSTagU/+74dO2St7CL4NpK44zI
Qdsm91E6oJdFSwHEEZdZxvElro0xAW+2ES7+vyk2PXD65lZNLsvBkRZem0CikCuhm7ly3co9Iup/
X5UjTm5qBocij4pl+IcAqZmeTRQWrxmqzcLquX6BupkeqLWOAQRywoclUgRN2JZ+d4JEJfUTCc5l
yHrPoCbaABVd9n1NSp/hpooUQCYCIr5GyoHpm6e23PmFK0SNAHvx6xM/RQoshi4HNHwjF0EnWJIA
lN+HgSrbalRoxY/k3nDG5/xEKyKBbw9sUGBKKKux+5xfPIylk1iwNL92ql36qKzMEcRL4Y4p/zkP
EPzUMHtROtj7cfyO5Be4+Ai+IA+MH9z8nYr0sLbDWlczEos/P93IDFIaUq8JyOBJRTN+K6bC6qQR
WrkNv+vd+GruVHOkifKuebB2dFKT0P6Fq9+FQXIHl7MeEoNWACMx6tw6pNSPIHTawq2kwRVWOZ+Y
3GCzSN2476U6TZlGGy9//FsBG75P5wojqNGUDRnC4ROe6ALA3ZnUlQd4dg0mZF+eqD5/2gMbzMk/
klKehonE784POPJDuN66cbqtp36/3ZOCwdIIUijKRjI9MMykdJ0rxtvEnsIWkFz/KsD4eavnoD3/
L/zo4aSTa72J+WZmYIVGqL5OVRa+xLSdQyr5rQqfA+2mmDaye0yd0h0r7p80SHiXOxy6NZC6H3Dc
bdrubbPeJ/Nq+lx1PSnn+8TIousETu6GT91rJbi4Q73VJNke/x6evNAnk3n6nmfXqtCAWp0mDoyg
kg9uRBL/CNgne8hXSCEx6myphGLwzy0q346BgmZO37FNivWyS5y+7ZJKTuw736aNWdyAtfKD5hPe
tW/4/GvAynxkhCojACAn6hTpYqmpTEk+AUAPo6dvPyiSzObngNkP/jOsUh8Y4wyjtRh14P1ACaJ7
iDwXx6r6gLIm7bvPAz2bnLkhC7CBpQZlE3dbMf3wcPh/LA0uubfL7XQ1pTEQ6yjP2HIr0FTROb0S
A2fZDNzyzbUZUPRfShSPFVEcUzkvH6ldt++dJaRNoqg5y5h9i+NpisoXs5dU9Tv5yRLcKUr9IErV
Md9H43xXvYq8iciTfmx5JhNhHNzwngrNvrRbpSGn6Pb8gl3xNi/+c2NLA6gV2PAMpZdaJpRLygh1
JlkGulLuxmXZMdLL5EQN6UZSaBMk4KAlRD47OmDzKbSFZ+YSDHUxM57U0OMRNet2t0qANYFjVrLi
3yymWuB6eL22/E5eH7+8YJhqG2x1Fa5Ehl5O4rTfAcXR8sjSh2KRVIMXqM2YWwPvILxKFaueC+pM
ePWCPj5t6JJn3DiCoWz9bfynclzWgiPX4W5cdixWen7RlLCzwC629zhlM5zh79LN/7hlcIxycXCa
/o2NK6XPN/Yg2QKbbX/89b5F++x6mATRXNR+anJAxY6RVLKPtYHMaDFFk8qXJjhaJUXmqky5rUPN
uEA+NYJczKEcejZb+KHJqSEY9a6I2oKo2i6Uev+pzCazgvlJDWQxFFSJQo01tNCLHFGuP7yPPLIB
ZxIoGfq/D3CFE4T8xP7wnIlBb9EjNeCL9btmEzx7z5LkTwkBbX/uPwK8F7Fgwcbf8Cs4hCdjmdgK
z21PGHk2Bl6w4UrwXRvDFbeyXVi/8W5J6qyXqb1d2V/Yc5PKJ977J6It/X5YG4KOtbGZc2ubf2f7
PoavONFGSS/sf2BVfuMpAVgZG3reFUXn/ZzNq5URj6H8EZDmaMB41RmxxwIXAxmuo4N8LVUzLQxA
pY6tDGqL2G7l+JzNTP9mv/49Qil92daDrX6oxLZYaGYvWeLOF6j8/9UPEl9TQ3HFnFODpjKQj8wm
goG5bUaqewPL5r8FKqROSzidjF5DqABuNvyKPSNKq8OavKRrcf/13CzBi2nAtFDP9T8bDuGZSgk/
VRgFZrEFoOK8kQJshXQy03AX5uJv3JeCXYUaBugdEYx0TkKaFA6v+hfERHLysCuBJxo0TgWp40T5
2hwC/Ip5KoapctQYpjKMDl2jo9PS4I3dRw5elK53JjdtZAxxzp9BilRzrMULCbOVlKZ0Hk5GO09O
qczczQk/7HlF9XMASSVzbnGI7GCG1p9uh4iNHZj9Uf5v4LckP2WXbo+L2wWqzYWbji2f9sWvZ7xC
hipvg/+WBfeknNpZlX/VkObrKvjicJswjWsNoWekc7FiNQysvzuZXJMl6xyAu6r+DX5rSpad0bma
s1B8F0/5YWjWVMtQ3UhP045stfDSIiYXHSvE834VVDlzYpr9J57VyQBVIwqQTR5POneUvBksqT20
j8s254KeRh+eNhJh1EoiDeVbB3HvpmNmTj8TT0A/L7mK3asDODjVQFx6XSY71+h/6VJzqRwpvHkH
jegFnrzrCni4BWN1X8gRYKYs9OUtJrXIVUoNfQlMJ6f2FJwCn0Tdkj0TLQt/abakrJtMrdNofNNC
3GKZAfAYP+N7DNU5Kaikm27dGnUSBY7zeApaQ5mAy/X11akB4C9/B/R5V7xx+PrUH7P3ucCKIk2s
e9gnmx5kgJ+VWmzqpgLXUVut0TSdBEPtPGmTRvsHY9hptLo+qHdwH6/FmOG1yYAiuwY1MpYPMex2
LZT00YgOa5WO+1Ka/jUB5UZMwplub9CTsa47kCRk/IiWV0P1jeryFyxV0fmYto6ZbyE33h8rFsG+
QBomnb2v6pN040HMFAT6ergjh5JbFboGDOcGxmELCnqVSrCC0BUoPhxs0klSklq/XxjEsnz4ZlaT
LdpfOCWjfprILdhG5Rtpyd42+rfiRBeno7C6xlALfQjWQqHE0RC6f3kpMmXQrq89K5B+sA4LyWT4
W3+fTccuQZ7fNlKS3GHtplHOw9/DvC8KS5Ykovp6B8C0UkDiqLbqOPpTqLRh24mxTJZvZtw7kbir
VVfuUWHcJBVwv/lB3IefEv8wiMyAojuTPZaSPvPNMoGR6x0tMje5iCEvS6TjqsGzFmQ2L3Say4Z9
4eRe61FgPbcxTueKOAXto9wqoQWIDGRYYTI2IbWmf3Y2Rs4j3XKOWAONkfZuQBY0NbgURWeg1a9t
V0+8F/v5XtT/GsBwL+wN11Iy3KFuphzwe9e65SK6vWjKyFPzxzo/+fw98BgxcDGwzaXHsApJRF/9
Jyu0Xw2xQZZEpCfYOq9sbpqBJQK9SZY1YAXpy44LxBVDbTb6zrgKXY+xK0YcPyNtNI8j5rA1JkIN
aGvlmZvbShrocjvCAefwhwV1tZJ+GzAWgcTD2P2cddAk6Pt1WfsbX1YfW2KmNMIFGXZSGlJOgcn4
A14GZ2Y5W/LslmZbdTwLoLKcxn8UgtwRxTHWrUfq2Yor7FfW51SRx48BeQfLw1anUOcaUrH1RfeQ
uwBfXxAcNZyNy++Y4vAGy72EMWgUawCgSy3C/JwGKvkLGKAIudkB+bGWew4zEPdgAY/7ujEyXfpv
sdBzOWDwakWRFFVZylxdptj162ii2Xl+Va5c31XO2yya8JWDdm/r8936UwH3rq58HPgsbaZS8fMj
BSjT7uYEpfXnUMd6C2vRkTs06SCPhET655aNWweGz1tWlbjfp/jGBuFMkXPGTjpJYdUu5iOTr3HH
X3s9mLgri1umw2ZEQBgQ2weeyeZTYvi7sXmBEBFJkarjiAfi1asROk1e9clDZobMcUyRgyzo2Y22
lK/D3nD8L4LjD9bEaY9G344RdyIiTNXDrpnnmI1Y5jbF8y1kReTM+lQrJUcMjfA+A10cS/0LXyHV
tAiFGzkjV3oN47ss1HMdl6Zru7CE80YxizY4OzZfQgobtR7XUVqt3FRWpY7prURMUTML9yNhnM1A
fVWA/RhCIbcD3dPR33hwQmd811gCptR5cTLwIoepGRGvHQSM7xZCPTOjSS7+AfNlMLXAcdltk7JS
2c7y0h82WsZ5Ci+j1Z75HzvUHf/+obxsWCfJ9V8a2h8avDlB/troPHmnbq8ym8qV6cz+AGkic6Vg
CSf/K3X5AIbW5RWmS3yLRUDf7TJ7o3WUH32RYwp7Vtjjnc4DiBZR1xZ/IsI8i0h+5OaBcW+9QUfz
Te5AMpu5txb6VQg1/i0fZAHs3BiDYOEPJJXfxdvyHgExiQ1ryKSdZzuw7nQEIdpmkOfNjLFBoYJO
IpmcidwFD9aGXsqIUgR+b//qgohnRB4J1YB+bbzqnzi3ifUVyoU2vTb9D1iWtOxN/DemhauXX1qE
vv9CaJ4dSQIr7t7oKCzoUb2zCpzEx2LPgCpBN7vsG7Yx9mgfR5VVpHFEwtdW57QwAm0BTpShu88R
ACC1oQAqGYOzCCgKmPmSeuBr30IiNEihkPBe5lbbrCOWJsXKQbZYBO35ug9TuIGNedc3ZpWpnWQi
YDH7Anxm4q1IGzEtevdW6LEngrKlJO1iMNyBIluuwjqI6RR4mra+yoQWzXZMLAVTsPcIhLG+JXsn
g/wNOYg95Z8ZWGnL8Cj/2dOlRD7Tre+jM3QrW9He1ijGVVGmdXq2LyT2JAVjx8KfUH8bCdaQ2UF5
KkrcAv+nLBMqSVRhhSVxYgD/0BDE+GZcyrTH0gX1FLtpqWMqffGFdFZx2ZNwNxSjguS8LOpT7mKv
uMiK6mtj+gsfMvrg8UuIAA9U31UnILDSiovaHDfMIWhPi1hAq4B1cnHTLDtPQgE3OdLoa99uqpHH
Q3FP9VZyBpy+ImmNo06FQGdcM60ucjv4xElomw58M9z6jl7SKnbxZNq/a64hbWEcoFRBV5quC57p
55zCKzIhVFPIJDYWwZQhbMcQlHHnVhoqEdgYKE2J0Ic5IUTSK7C2blCtq+Y2OjJlqkgQhtUbg81E
l37cE5Wb04y4vW6yaC2HhtjQUoCjtuTFi7S0UenhOSyMmEQhL4EMlp+feNTElg70CI0hEskKGlOU
mf84B43GUMpP+Db7Sy0SOMnGna1SGSbOrRgmI0tDGJ6TAZ93NKJnwjZs52BJ2asuVYVqPnTfTDco
ZIhNK4gbxNnsUOMm2saAGorlHYEsvhrFyppFBUTeybRL7uIX2gBv4Yz4E72fBop9ngdpXTWPZBYQ
KLJ/4WqHxn7plljJ23nfAe/wPrEt8TrNhavJMfQJ/f/oJuKiz7y9V9h3X8HSA/tygi7vs/CEsu0F
EYgIp4h9eF87eS8kZmyVhHcOfRra9FcRCF3TssM4vkd/H/q25aEevrY9l2eVZF3nK0/yjiX5mhvq
djz9rGzpv0/nPBmSVcQgQm+/LcO1veQBbC1XcTQE+zijauuXdkEx74OrDdG3CUU1kp/KmTh+9uup
Qe/nlH3g0im+q2GaudH36ZDf2K9X/vY0EIpwYcBYs+o/v3XCFtyh27tdLaukc15976rXDjCLt9r5
dF9FNLDaeX8O6E3v5VQkUaKtuCk2jaFK9LuOAL/F63siqeRvAP00Q7XZ9d+FNKmPsq7UrKsQ69CV
l92wH9MI8dJEPnMZnEsHnyMIc2riKIBrGrLOmlmdgymvAh597x/fOy4PzDIBr2WvtfB7O9l+bAns
mTxd8pFVe40iCbr6NtZ9b9o43nil2O6Eu3xrbrnuGT4HVy2qM3fygmEorKXgCK6KVLQztmf0z92a
uXsqLUxrBo2Rcr1TIvbpgIC0q5s714UDpYTLwiDVuKOmrdyvf6y94Spu43lepQro4VjLJi4w9Y2A
S/nwGn+qROzS3Ih5xlnm7Jd0rOqCb+keWGJBvHFMBOBhUt9hYMJ9FyXXobx1oJchdPXRDv2biBvd
PQ3uZgQ47ygfUkND8KqdkejX4Vmr5lhZRSGbvz9CqVXE80cGqfS7LEiK4ZkJO8pEKFHWFdpxM0pF
5Fbb9+DMNIN2X7ZWcGYrbpErUKu9C18WKXse3Stz+jXZ1+4QPI3hu5eryt1jaCR5qX4zH0OcWCKt
7hv9euAtcBb0QMIfLbKZXFDBp1AvMr+6I7JO/jqWX4GY1pJGK4zeUjxiyd/qMBAMD8M5qDqZF7qx
1Z2HvRRq3yX2EO6ONnXZb5bcMHahXC19SYDQKU7JjH/KMGIKcyRQ2IPouLZbdUBfbbYCt0FdtFGn
uJ5j2bbJTGro0fyeIUzzY+f0kfqsq5jOMoRl+w57xT97GvWc1XCYEBimx62JA8zdvwwue+HpSv1K
d9iM2TzBEOd6jy3dUfG3EgseyEqwev0Qeyb4JJohEqhDE1zb/JARwZe1uC7BTsCxuUz8FSuBHrs7
fFfW0tidh/up1n/sRFc0nVr6RfXwo7xMNalKwlXzjFeRvVTeGAjiMCh4FQ3AJTrNxiqTAk226d/9
sYB7hFQJro6ejlf9bQhp7ukRXDVfbSurFWRCl45M//1J7bfcK+7tLgWvK4Xy7WCQEbomLTpXbUMp
X6cn9Es19soCHyoy096wv1S85JaR1xf83n7yknyZUlSKV3eJz1vunF/manaq2n3G+2CLkhn0K8Z/
ioUwFRXqjpeCTGXTgW5Du6z7S5SMzLUpdprzvyEnayJGIyKFIqvVOfMoGZBDhVk4WgVEmvOLa6ok
2fHUcMhQUrFbr8RNkXjoLqVzE6jf0wIxHGScDbwhG3QNUGvCbVObx0K3NsivzbRaIVVPjIXzLlby
YHxUBpWrpHQBNuSZqXVu9NopyRM4nt9qjokyJQPH3d+OGXO+buKn5MkWFS6W0OHXENza4o6TEVMu
TqcXFiVr7UQnTdZicfEaR4SVq+oik+BKL3F/Qo+cS6Rh4KhLiJOTH28yimFtgxytmBn6UOfZ6jCS
Fp59Rbrt8pdMnP5bxoUMWzrq1LAa107sB8eSFtAXZ9Kg0t1881lNs8fgY1KWcTkpxe1BrtxA1eAw
Up6aDeFEpaZyBbVB3bm7/5xEBhYdFS9byLfqeJ/EEArq7T2TLB/7tKOEqkaT1L5LCMs7IgbzrASJ
gKk520rmHr3LKIUyuxybBdUksSubqzXGF0yU+C7npvb2Ga3o5RYnL/AbMybYRBBIlNaLibbxFA6X
ufVtkRVxC2FgL1gJH0NLgB/w4sYHuql6yMF3mXnD89bz6xDYQJWjYsRN7qkeafSqc6VfVT9c5bu6
k79YxPn0FF4Dp5T78lisIWJSE/B2YzounbsineFSkhPP7R5Xboyfl9QpeeBz1SAoWxSSHZMKl1z8
Hv7VB6ZfdXswVWusUYH7NOdyH7hl9hay9G7pIzcx3ddL0ejVs8+dg1Yq+LtOgdgQ59t5bwamK+up
yKDQ1Gaxd9xv7v8EDhHXY3kDdkf+1HY2Td/XkY9xWKzato/n3nPdNgWzYe8FTDWdY8z7L8G9ndg1
y0G0sjcJJgSWdZ7RB+1bN6BA6DVS14A4e+5Njqe2lyUImWKqzqly4p/Xq2eHg/UIL8zo7MxhfYiv
r4T9+NnsgoXe5rZ4PVPMHvP5EecCLh6tLyttJ1prDkIZe5H2Zmo+6mdQaZL3k559j26bf267TgeL
8R3VNxaXc4CrhdzXZLgAeVLGbNvaw2GJzCcSWk2FhRfPUK40fEiLsrOcST+bE9y1eU/wKVH+N87s
lJabJmFNiEeeosuf3uk2OUCp/AbwOHyxGzu5TXomXDSXghWSm9KrgV7zyakKwK+m066z/3q768y0
9pnslGVRoMB/OUDS2EtcsJ2DUD65OjEOFCUz6EUdlvOFJzmDnq/Qkdwwvi7ex+2PYpGMopT5s1cJ
wVmUvJe0a5lsrD/0DSXnBaY91ul8LDWnXYmRy45LVh+eW3qeQ8W8mh4ORUqjdsArugu3al9YURof
lLfyXVp2MroiEVBjV8SaPy7TnPgisSQ1CdnBAmpzynOBTHL3PHtldoKy3njPnlcy29pL9cCKiMTY
JiWmgBRKZghRa3hbCR9AMphUuvufgOuj8KGYScux5obiG8DgfyA2jO/LffBy559K4fN/y33mk+na
NV4FBSTWt/0KIq+ptOHc1uIg4Q+hIU9oOLHOM3V6oInhgLZCokLcjYw0ael06QO7H3o0Ak3bXj3A
HRw+FkLZnYNQPjm04jIX+NK6qybx4MIPjIw/t1B/zi3Iivok4o6oHHfKpfIJFEqx1dN9G/5fH15H
/t38a3CXCmcL1Y+CM5jyqXDe+QydgiCOTzUZRPC09qyclHavsom4EK5aOOlpz6u3X6zAvVVKCplO
gM4jeFbOFk/2xZCODFM6jnVTqwpMVYE0LcEhfm87euxIfFXwTKixi5ilLjE/Y/FPFPC1zvHubCdM
A0J1qe1ulsg9lpPUcQtLN3/njdZlAG0SZ+wc/XWEBLw/FrxLhAjUGyU9R0FVzu4E4Tffy03YeoJH
0dntWXGLjHmFsP4221llgDhtzIMsl2Lz3E+/Ft8REhl8bPcszFU3UCTW+A3JP+SzTNGnj/aJC0em
haR9kIo2LOsLAoKD4CFIn38kpSAHGNl5lR0x5StzXjH37c0okmyBhLFWVj1j0lwTwKRP7GJrKi90
CtEqaIJNoRyVhsGz2d2HMUfqZKaaaWwhLipOkydzsXnz2/+BIKiQxJGcAY92IyQm73FJMdq3GlOc
xpMcpiquFi48J2Lmmf+GLGr+FxHGHWpsTFu56oEptIfc0w3OxlhVgB0Zxz59sTLRccbeXrBw9Q86
IvpvQj1mIPL9+qoJg2xeKclpOX39mGcehGZDD3eoE7heMgbYI47F195ip02U1EJHKfnY7Eb7iWmI
RzzQ6dYXYTlsSjHGE/vCfBQ3MlVwMg4j1ZZY2UNqz6e//HhqFq/FChRwvlYuy6JRgnlWWAMgo+IO
frWyptOZHql+SCGiC4f4bsmET6WCZOCSz8C1h5cTl7t67RGeBcVyE0KrzX3WdDlzWvzCV1plrsyR
gZFkuUY/AUIc7N7JBB3c96tps0mtZYG3lJZjIwXi/h65bj7/yZFC/IdJ/pmRkrO06eo0nsa+MdKe
dWfckzSPYWM6X8XYC3H7xYhtzqsaqmd8WQLMm6XKL6KOWTQcl4TNGDxEek6Kc1ZBwGvgmFVo/Iem
abVkPdMNHKOJX6saeIzUmz8qYMKWHOCkN6OL38kg6mnsRkC8FylczDdP1CZWefe/J4U7pZDfVKnu
3W+DLEEKAp951M0V2bTA7ys2xiT3kX2JydjIgYwXYE17LdYQzo7kezP30k1qmYqAifGazGy1i7bA
keFITXq7XOKM81L6Ffb3RMnrGnDGEHi/tJU4hNos5+TsGqifaN02JGnyvph+Dj/PZm4ETMv04xyl
smpvZsTCFbRcLebcXrbxPk+7aIOT+kyJ+HjkSEm5Ot1eqsVbASZygyZk8wN4S0ogdDXKL1SZk1H3
1IAnOiW3bxjSVmLEIkpyMYG6CkPFiz5UWdyzw+DHGsxQobAygVvIFxqhgdoZx3Q1iKoBI9YE/1P9
zzPih1+59YhAVXy9J7fQWxFrElvWhMVrXijn9y8IDc2NZpVNs/4dgmPpJB8tlyDC/bfqzrrPAMVU
r/YXYkURl6Ju0on4JKFAqcFcmQMWdAM5wXT3GE/+1DCKW5kklcoZEMfgqSVgNuuJq8ysR9sLckQd
MxyIzlxnQnHCTUJ8Bze7n8bBm+tFvWgK/ebrn0Agy8sHrv2uzbZzwHvwvnqEj0NShuEAX7c42yPO
ov2+vI/9vLcGEdsqYIJ0oktQ1mqLYV26qlH+J+vrYjZ099QdAX6zpW8YAQtTFIf9v8szZoPAHB4l
Qp0R96ch5jLYG2xUgyJzMGPCmAjWI7g5U2P3m+ZAGgh1j/0DpVTXrRcLuxI0JGe0n8P4+0Rz+xcW
neOBiCN34xuyk4VRhBvzJixpuWQSEUtgQQmbD1TFPtabYNBEDsAZxckaQaLXMykNfubE/eQSh2Go
y7lv3pznzIQeUZCfoZgpTx9hYAL1heoJY4FhYuuAfjz4qHKn0mrc352UhLu7Qm7FO2pFx8jnQRQ6
tzu2aWN6NUoir8w8Y3iMpgGpx+yUrAX5IPQrvVF//Q1vMaOIRqOj23uK4vO5gr+V4Fc+XKeTtbi1
iDg+68ehew41upcU65BpbSmURXdXA74QiRiRUcJqRhz8b5GPCeVy/hvtWvYo+A7kw+vFT58D8JvG
9WXLvhvDW/AEAauAUOgFNWuRjvgfptaCg9MQxlnAUT7fok08xwaGzgr9sBi3mnV64CU2ZYqtKOB9
f1MD/Bkz1Gffa1dJTpzxTwRy/ikMLTN2rSVGhOLuYYD90IzkmdgsIQ7R3BLh7bDVmu4QSBu/YFXS
p329cY5XEu+w3WWXNM4DII6BnKFUOP3aWbVCfE7rkAmgiRK2dyK7jqrVj/C/4ygNj7+UfJTFKwa4
riqWX2VOVy+RcYJ7N+1MtwhE3O1Ja8E8K8ctqylCzSkfgeTU5j4YbwVBN+vhKA+jQUV+cuN7EmUF
Ed/HuNh9NKxYBN6ZuC+nyzNu30+ySCr+byVZXQTv3E9lt6CD0Vc2ocJ3lKEA4cRooJqcnV4JOaXn
Q2afsKiYxPmB64XW4l9jq7pUHzSZ8A66ERoxHY36/eWcr7A4q6/tWQdbg+ZIsbWsaANxhFZzTyB0
jN/SRSklUPsaaPs3boVOtCdzkcnTSmv2AAsYoVFe5iQp6SVZxYCdrxcTYu9SsBGrEyXTa6M+q5/3
z0XUkDvwQ3QpNoSRLS4ntoCE1agomVKuZR8rFFmqDJtRWmW5YBwr9Dgqd2NvncF7yyeEz3q9uPfi
HbRwNWft3D+vIutrPVL9MIcaS2icSXEyhxigfOqzht3qo2Dh3OnqAnFmEtkAZMlf54fBCEkBsuq6
IvAQRMozwSzHVTmkvyQJAkEEIloACW9ZH0+maHI2A06Y/yYUj8YUvp5wPChLIcPwVekL2/4yvaEU
+5xSW+OoKL93qO20iQjxyCNYO/Rwy43JmtsFxB0s8t1VSAkVkPwiY4ljsFJFcYEBiqb80MKV+/GX
M+p2nVp3n9xowYxtndLNGPzdLQq0f15+DZVVxCbcrX+nkUUMxw4P+mHTOvQIittlnQpHO5O06gUh
9DUWfAa/XHzsJ/orHGEByPcYDZzkfNXv7F10whXHOa73fm28Hex6m5P+plVSpOnpm+V3mfV0Hq79
zCLNEXyV5eOFSOh1UMGkJxoCmvPD5jgr8XZeCl198C8uTpNt6YGNUP2be+V16lh9MVTLNw0Ej50B
GfLczb8KPCtb3m9D7uw9knbGZz1/Fyj/ln3DXBMuN4t3MfucgNRY3ArlazjIijh0opGAZLPWkm/a
R1qf9tMjbaTahYfZ+rSti7EYSp3z70LgDqWN64UuNjZaxCUMX6hVviFMxVL4xS7fR/bwj7z0spk4
+FzDTzGjHLIZE+Bko+q9w/5OZL1XWFkWfs+/dxGZNR+GNiqeie97MR4O5xUVgKa/cQofg2MvPVPI
Gu6R2SesI19NUn1g42kNJ9ebdsCt2TjlZsiRf4rigwBFdictyASS1tYKQZSuy7iJiFucnPwZSWb7
23aFno3MVr08fqNijneuq5vYwYaLm/tLz6SXD159SCj3eyRt99UD9AEYtllCIYtAmh6plrxWLlNG
yUmEknvWTtnox+PjcZncR/BDqdQBnxBzyCV4QS0muzKXDwJYb88GXU8vQ6fBKbn3PpT3r16Tcd81
NK649bJ4tYDkVTpEJfNz3WG8avEknUAgvgCbz6Tz9BYqRZz6+6LlLm8cwNqRw0nmH0acG/gmtaXe
A4OQ9D4x2k0atCoSkenI1aI43tofD0lCgn3JJ7XOjNKGHqOxiw2g5V20eJDcwBs9YuNMXRZceAqs
B2xFOwRh/Z/Q/UAMdx2POwvStpoU6xq6MRf6LIAbVWj70zhqQAeCCO1X/9ossW+iC6iQQYTJupBX
Fim30rDZjGtrTe1cd1nQHsT5MDyXK/lq/uJPHoyXbkPdtt7928Q0fvrNnZ+Xi8uuvrQi+fmkQf6V
uJfrO1tJKu8JItVjuteQqxC2OMrSSfDJg9cULPm1GeacqWMVokUndQWKIPFE+iX72sWOzg+IoZjj
M0gSJ0Y5gCiRS+Ue3ieduasV9/Z40u/RSebgasxMLMpOQvr4FCzENzHAzP9mNAI/aZP9K8gfWbBh
KsP8OqEJxrAiRESocwwIiOSHq+VT0FB6u5YPAZO3J2hrwKisIdkQchvTOG5qtO0/S82FQJZ1mD+k
hTZVgtFrF0dBwZ9dZh6K7rbs4lY3OCxCXBckjZKOyBpzu99hLSJtgJRoaxWmddOg/RRwq1FD+GOD
09RTcphJfC1/n+/ulpA5oc9Ewzkz/jNRUx6SL/JyFVtCG9XAXk+iaddUB+u5EEWYj04GpzQFYJGS
GVO0vtglZGmJJjrgvRVNVbqC6UUjZHnR4IsSBxPSNukNJ6Am/Trb1XZxZHZ0imhhw73fSc3b+Grq
kkvXZ070/0tFyriSZu+a+4+vANcx0XmdbQHWjcs8Mkqqv9vhmGTebsFfPa5LdRybFFQnEgR77ie8
vPlPujbPqinvAuZ/01m9pergrzk0CLhfw+yXsuxkB1BfXbIDWGTjkyqTPAZHdqWwyf7ZCPdLIYQA
Dcc4V0x+yQIFXjsL/3BNHPRx1af4AKXRNdC8rgTljZopN0JH01wSMMmGlAO/70bT+T7otv/aArVT
2Iq9dZN71nikKtvEv0pXMBXO/77EEMQu9PUeXmOMstrterWo5F+nchLxF2cM96skNNi5CTaKriSy
hevtgkUU79y8xMdlQrhVWhEbXF8O2KkB18Abk74zuVA3VVrKo4IBXIaMNCwbdAYUmjvWTAsbbbML
irRdiPNoVfMBoOP/HRNFbxfTbfS/2NpCfw16gmxuv2dY8K5JKqzGbFoXr5UNC5xSGYgoXLrMZkAz
ul/9bVzz2BA9G5am1AGxiAaY0A8luePpStN9Q9F/AmxSfuZSsZoRM5HJ7Fkyj1d1LpvantPbZLv/
dtE2QY8iZDkfmJyVr9x6c5DH/cOkswmG3C+152pELKHlQgXfDZeB0H4vqxE1L5WpXe8sp9Tc/OcC
sE4zwNSQKefrw53a+79P8bQua1aokbSEz809tM5H/I3lGf134HGAprCeDrxp7ED9xp/28WAxvefY
DUWGbvCwNrx78hG/C69eNwOKLGwyCDFNV/kAwciHnTrz0l8gWP/KowfbK3jclk97vUdnUy1ojC4a
U3tX+9I4tKw2X2sx4bwCZPLYOyCbN1BzzeD5yywXwVz6USMsG9yfXW9pxvOUsb7wFb8JfPLmyosq
WlpxXDU2b0gT3/vxq+lwPpGC+jNnFh/iJIl1Jx79A2dHebK3gUU7PRIEtRJaicOCYTTE3SMfbYyz
PCnGEx3T7adgYDOKzMlEj5lnQyeCB8auQq3BGoMZ/SRSGvVsEKTBFtI0+c27/51KWeBmu6oHgSVp
rWKhATPyc1ECJ3nbLX8EU40jURbU/3dC9wUvX922QcRaO+B7+mHRUMPeT0MtMVRp22ACbUldWI0X
zvONaGrwzsGXds3+OrF2dbFlIy6a+kzKvlvx91m3PwkPNW5gavrvO/Kui73kH9Bz7te5telu9iLx
707Ul01O677W+twRygOpI6t7Qnq6x0FqKN/2ZwOntHPwPoYIuvH1Wjdxdfesczhxja3997lHxvOR
47lcGIOjJ4U0yW+g+RlTyzsUb/xL3D7AraeCF1Hjkco5cs9Q1k0jKLmQF+Ckm/bfWZdGNcAKn1zi
jee5em/pXj/0dIK+KtKIywunhHdUeXuTcRHGqmODA55KAp1Z9cZde7v1ysEl5KdC/qPzEeJjSBWk
7SYPEpYyo7qCKchq2PIbtRXTjbsmm7FchSz+gT1Jci85eC3Q5wigILDIE59HNjG7QpCCJobaWTB7
BfOL2FhANmxOuYO6RxjQyMRdV2vvs/fK4tXrQRF/ClrcALVJdb5zz/xecVB90hbUAHblqZ8r54a3
bOARx8VuWwMrq5TBl5ibOcjtsiOkX+zccBgCwl9cv4TbTJPpxEtm0EajtKOq8dLglcd1cSdzCiGz
7S2j+DLUOyYl876/9PNGeZkYC7xFx4X/1tTgZH+5NudqW/zQElolA8UY3ndfafDSPW5CI/59D7Zg
nfNWE1jMOqIfnV/yr+4PaAdsH+siI9A1LYARYjUJH1MX+RznE4SxAZO5aoW00fnEYP023CHvX/bu
brf9NgqJavkPJNF29S7O/PL7ugDU9jLlT3h6VmNex5t7LFjgj/UfuFGUjYhJT/TXvx6IlF8KXZrd
eyLVmnHoF/qSppiKY/WIXZAk34KZliD6Bv4iqzOs4XswBIIvv3rD13MI9gqpMHGHUV2HopHXkgrG
M3SHqARPx896Hqp+O/4bTNeMVtQWB7ZybKvVnH8lmcG1O+92iFqMy+M3qo4zazi+tPeJxkv84JHq
Hl3X55dBR9k6/cVfvXl5Zq/mah5EqrM7Z1fRpOPHnu2QXRJ1JOkDjr2anIXImBLYZPFq14B8AekB
YmymLhmUGDk1DpY9h1+z57IweCBj7t4oRlR2PFhKSj8Px0IT9XDuOaGgy1XlQhWZHXoKLyzMhHNW
j/cBfNP46D9ZMR2czsqaYbpOVq/c5FRFc4XDzCH7/eP7L82VjvOEbHk9WWE9oeQAQs7L/YUJWgVw
mCn2eiaQqe0S9nXjVbFxhZQzhgpP/5ERr3aU/VozfDadyCBTxR10/8vRBVvCqTP/WjWdAR0ZOLRe
fIpsY7R7PJ99WsQgBlX7geHGT33gdddfjeAkJDiV9Qad7KZi5AeQg7Q5JkOMEtOaSYZvCkHP8dum
w9enho7D+GD9hFwaagDwy/sg9oXw1o2kWPdHyyXaHpRC6/BZi6C4UR3J6nNexgciGj+GsjdBmCo7
jMsJfZAdQakjc0ziDbCZgYT5E8OqrbiyRpHy7sSxKi0fg/kDUnYVwPhwM4abQqQR2cpisXpvR15E
Tzd1Xs0fYYf8n+YUcX26rBPnejXNHRX4p5q2ZIffXtn+GFdnuEz6Xpvp1naB1wljfqNKE7QltsN3
e3ieJpWmG9AFlmySs71FAvcdE7KVx+BtD5U+9o2mAr4a6DR0KjnB9BaKRvCyaTR3bSxnKvpv8RP3
7NhpGgM4q3os50U6jy8UqF4zBOJLmv46Yw2+l4UzljTslFGbb7sLmXQTadX6OzLbsM2vusXJnfjO
E0QdrQtxyz/WK9goUvKZM5SSWcoZkIvfhAYshxLjouAsFax3bigFQur8pOVyOVKoXr5XfFjx29Tz
U+k1BgDm3gP0MJP4/W89SR12eDf33pwt0dmfoq6shKasPMQarjw7EQ3YkagKET9CVuiG0caZ3SM0
JxipAft682W/SnB+RDS6lk1ZUcguIUBp/psqX8Yzup9BTs6F8V6w9WLfUowq5h+GS1+hEmQhR0DM
dcxRdbvGpHqrhbBZhgZ7QcB9NsRCo4uAWg4pKeNnTBYhIBYFbAWHAOohmettokOW7uWfiBk54S/Y
V7jrKQBroPP0EZ3h5oM0MFp8Z+uT2D2Q74SCMyLsNXtrFs6qcMnLxyOVXCbPziW1KtgjRU7QVtbo
pb3dFZE4cLJJmlbhuxLfvMVzPBKXo456iBlth6T8bi+Sz/Ff0f4u9EZcR3BFQLxWB7/EOXXh+RDe
0dwwUjbLZYxH1l/lgmmxTUP4TeyhN1B7aF3H+hEHquXipYG63xdNG4S2l6rxb1dK36WSlxJEe5ns
azOnQy69RCFlYBL8LeSoXYfdwXhiKQc/DfNQQeaRD+vPbH84CdWAB7EmCWp0LSGuUNj3TlSXzEkh
iYKsQXe68w8mN79L5EdrcWQXRS3pYJAm+Wco4F5MMc/CunOLf7LDGBNzo2hRPriZVm2QQ4Vdu97O
iEwdhvA0aiS2cWGxZq4LoahLAUAqJbzGs6aWhU3vpU4nVqpJx1jBmV+lqyqTk1CKFN1WyAU4P5QK
cBGrK9jvZP9yyRW7GhflcK0Jn2/uhRmdwlsB+LUWHLp1t5FPzvnnV22gDQjU/c+29dmsuaSO/+ni
ac+IeQU6VwDW0cQnJaoa57yaOtpTvrsB5DOOVl/MIifbPK7FGbQYO/ZVZMDzdvX6ykkgPTruaZ1U
Jp9zRsXRClBgTWdxQWFzJIay6uEQvkXO2rj29VZxwvIDb6zvbnceebwJF1nLRE1gE0xQU7n1aHAU
xMj44AcMm7qscrgxqLPUiHBRc9rvJmrjAVYYyAuSPX89JoZoEdUIev8O9xYa4BuD7aNAaIsyDvQJ
LxXwo4ylzykhsAv2tDoT4NF4mXCghcbsmdx0hynjzPpyOPNYWRZIa8LfTPDUNbK/0FlOFMDvwlmx
i+Sh4EeICfVHChyOPV/EQLutJfBkeZpJCVu9GDKRmKv11AJTaDdRP5NuXPAB10lySVNLHpS+t8XD
vovcRhtweBwJC7GDKXBcZl4sGCAE865NW57dZLc6EhvVAdEwgOz31YJLcM4VIemuA7pR1V0Hkf43
nZiViW1lBVHq+HPt2OjRJsK1hvdzUu5E1xgZBABKAP9TQUE5PfMmOt/FnUysUtNObkqIJKgXMi6Y
JZOQiRjnSYoYgyecBsjZQT434aITLm9X97Ua1MhE0MUZHMsSSIlsaN4Yfv+eu05AECHb3w9L/VPy
iffVHUVlvqaT786pYNCjtoS2iLWM6sqk8A+ufYd7tAJlDjkWi2E2rfI7oa/mKxqT6cG9wViLKgbQ
CPH1+7oKS8Wp7I3Tl4iEaUGhU6FVipQC/A2wVgmh3UAGuB0HI4e+3C+hWz6BqwI5TRVSzvK4ot3P
nolEm8opwkfwginFcxoAiSRwEnN4uNCPmpIgDOGRhfq5OuzOw2zaa8+Hsb9PiQZdHGEP0ddH4qAK
q/3MqUG5VVjM3PbCAWblAgcaSWV0+0WfH0mw3pdAzr+Jm6sepLkh1Esof8lY/pYcLOe9cIs9VkEX
/GL24ajArCt7k+84p3FaPw8rxuK7fa4M+TwYs7TkKZU+30IqqTSHxkdlJ5dcAJmlVfIp2NPhB6TT
EPEzDy2RoSqvrDX9jfd56uZ5WGV7K1zhWDdDMxnQXwyMqLGjjpuoXiajAduavbaU3hp324x4Avrh
M9GjjizHb68UuGU2afe8elQ7hVG/AU8QWIijPs6jMV3m55XRZusGs1HxvF4CAYURL5F4fQDmOJCe
DVnHJfOb0xspZ/qFTq+qrYjc+fSY9kHzCiEGUNJSzTFgbBUoVEfmnnpWm4RRgvlSkj0eSxWvEedJ
YmPUomW9kQQQ9WQ5qjUEdQbDez1w8oC+EjiM5hzlxtQ6SJjELBH2xturAxvoADK3Ykx9A8SWqspO
pk0JztSEw/bVsZ8ylhbzInwozkcUI2+ZRlmLSnQ72sPdiNO5QevDyNJrJ/hzs5Gsl6JlyYUz2OOx
T4aiUssVpv8gjGMknFmMzki7XHfAafr4mklt96ukgReFupqnkN+4p2/TLArBc4tE0ZPdODCsqDaI
HHssW+xagXFmyeBKcipO+reKRVRJDIPj6jsHeCq56H3SbY6Vpo5e+kY2whZRJxHYFBMrmA8w4nty
AbnmIO6lSn4HW7zjL+73m6+gRc22ZMR8Hy2CPdvaMU/3mQnoQ6PmOCPcfLvnGoMUBh5zgvVLnpBZ
piIw3cwuBM7XrH3uCYfj+6CUIc7T4NN9rQ7b+LWLpUxfu3eM6HU7F8KnVt3tQpCHvic8alBgi6Uz
nH/xyIb2fHDbO1lxe5Btr2DaL+Ff5pF7NKP4y8fRtXiotJ3aH7+XlztYTiU9ZFy+45rvnxHVR2DN
7/u7a9DvHwKhqJff2FppJIq5pZ989I2ZMn7tj5i8r6w2ncaI18mAngKSK6a9vgDZ8PDdPG/QhMTJ
hiOJDX8gFn/gsQ1Coyklc8BwRpIFu3iXjFa7JQxwB7xKCO80pnIdU1oVErI6Yyc3PRrguQ/4zIxV
NTkjrTvoBFElXPtL8fywZ6L98Q2WGVvRn7QIM3VnZYf5O+gqTRkbKIY4FrVqjTTbVijlecG++Lu9
ILa54bn9pXpLNe8jJPoNlj9b0BiqhdJhlJIByfh6IP66b9EpTHFilsbaSa4D5eCzM/1JyeifdTBE
GcbNAbJKBbo7tTY5w1Vu8gG1aOWPYR/stw81/urHmQWnk6ZWKPj9nWpR7jGm4YdHP7jK1lMOsY+Q
8G0B9uJVLRtq6A3aGPgf/X40dlsTxvVYNEFLJo7ief5RNK93VnCPG4LI+WpcQfmXBCHOXjGH8Oyj
iAxu4rhB3IPYwmCwjXn7Q0n7hBLby0MytfZQkOwU9QGtGSeimTdioivZykQ8oM2fkwMNkjQIy1PH
3q0F4pMzS8pmSR4DstfSw+t2aWIIIs8jrZUHQgq5f7YR/nED/IJEwgY63rfi4anF44e8muhvX8+t
+/e98OVDNkP5izDq2VY7LDqUi1ama/3BcVWRwbHT4jRzsChu35ydM7/5+MS86Z+kyxcD2mBWMb3Z
BI/hl9/vtEjcdl7swQVqkvddllcOxek9Bg3X+46+wpwOGMy4prosNwonZjon/vl3WQzDmQEkQ42F
/IeCS+wufYBL7TVPGJXnqUwJmPCX+HDHqVbbt356XjjNIZ0I9u3CG+5JohNXeiDgfjsXcS5TGf3c
XepspB+6zLrBKtFdkwEN+8lQ6ZUBjFrDc5xAYqit5lUWhV9kBvayxWfZddzmjnarf8WQs6nWbBj5
/rI/hkkLEzXrOrA1q1dRrc6rakY5raKZTTil+zDlpp9imT7Lq4zpGiIj4sY//1C01bTzF8Bhqy6h
ujodyvP7Knm2V4t3QTQoIyWHWBWJeQLeGT3ET+hQGzqq7gF+s5Ry2ARgOd24NeYGwt27K4jZNO/o
vWBTvravNlt2lH7FsS+KfqGSQrzmjfEbOylu6IPHTQuYcdHPLBS+zKLa5zQA8hXFlokc9HtS8ook
0enkXsS4VWf6npLcFz++/EFtAQIvZrZTiqltbbaMRAsjkSyPnLuii9ne9VIixMl2fWwER9ivqfjU
pE42sxAyCtwwIk+1+R6bOVVq1f5hVQX9JpFYrApYOTivc6nMRKw0wn6YY06WZwPp8r5wZ/nsGJSN
ScpptPg1YSAnRdKLqkWs9YrLadp9W2+GVPzHp9pSmNEtrWlsFjB2HozXOnVOqdVF7AmvN8MLml5C
DOYrXyktnhns64vTw/5Bn/MX6GW1K/xZTPbpZsnsdeob0HA0tLdVwEAVNjYrQHCAf+eW9V5UkbOP
oicUUReJJG73aLymwoeP3/JSYUPh3HwbiW7PviVLtt1NXFmdmhaJfOh2VhGqZftV+diMIF4N5OdK
MqCRWi/1JPov5oCpPdgIScU8cQSc1rNGaee1LS3fMkH9KrboQmH0DzQBvqs8vHZObnMk157enkyx
bPrO8Cq8VXil6Gyd5f4ohzsxtUOvQGc3MHR7dqTDmixR424v6CfRHUienq+gMzExTfwZkCelEewR
fhVfWYuN/ldmHyACJzammohUSXCk/f4bWT35X7yurE9tLiDEQfY5qqMpyVPRcW2D51j+cBYv1lQl
VUG7Ac4PtWkBvKRlS3329F6bKTtHGZjU8zhoCAKVk6ZHLD+GC1LHzR+XgmH/locQnnN60YZkvHV9
ckVqeHQG5zSug0yWigJT1oTiYk/pzS7tjrPW9lQ9WSsHuDZ9mw+PK1ddI8whVu4VlB/JXh/wjIOZ
2/URhmUji2TSX7bGijbXz11YRXvEeyJ3L+vELeNdT/OwtdI2ZIatZ35RzpySTcPV2LG2SHMsLCUZ
xjCdT+J9kkDPcbEu5n0TQiAvOvjczFqd7Hh/QVWlcX+GE0A9GNTxbx92fqov/0nhPLBXRnQpF7e0
bGF3HOsbGh06FOoUR7kugxtlu765N9OeEA16LI5kh+RAtkq4GOnrwtgjF1uH+Y1kN7bdpj0aNeSb
eWyiqOzTw5pTxVxduJef0rTSyofVwlhZ2Zb4X0qi1qXs8xtjgCEmlS5j7H2mWq0VHaTU1A7GLcEs
hOXIPsQyTeZgSd2t0cOxLdpA1XQ0d/xGcY8Dhuwt4fCjYOLVFx5nVsI3hHrpXsiNL2slr3Djae89
ycIuEXMpM1vPjNYUW9+plKvKFuooPV64MPWHpcHvobUcwqNXT8lFgqf/UPElElrY6F/qh9QRFQyr
Ad/h39KJSnGUekVucHwcegymiqOT1QLoZMwLjKE9ldL0b03xSOjESFeqO3BEQKkeSH7eOMl/6MK4
QCwG23sb29J0HGucGPXWFcEi3A4mB4G/OKsOnALUerALLvLF1rYRJ9BwmnNKyqSSVO6ZBz7XQx57
NHkTd5g0VWDLDsExuM1pDXB0mJE14LBpRaYVuNnjzO6pN//nELeAydp7mrDvEhQSVivM6QKe3VDV
EEo3TAB0ZYf1Z3rczyI7+lQEN0ChiiwXYesS/lWsr0ZfU1RW+BFv3fK3O00xMTfWfYw99nSyCGtn
Z+93uVSbzUdWXT3eKOMwJFB1k422ybT5Bu4NJW9daOmMIaAdDKKJ5azgGNKrtI5onnGsHLeANb9E
WNGGUcEPJLpiq0yK2iBXjFwznMdov9zspjYGl9k5onn3BI3IpUGK1NrrgI1UMkWTiavQ4ZP2vxC4
CXegG1tWUoll52uwYl/FoHqRtrtnqUFwdM2Y5ejpNFP02beA03ubDI5aWivbOSteWCfUpyZmmHsT
Ap2aWKtsicQne6XE33k7CncYNlSQiClo9X342zJ/23l9XCPfofq9aXxbUUgoX1T4/TfhH7YkkybC
HwZiwCEB6qn0/ibZ7pMJzUde1dbw3bxbdYePNi0fGNZWG1V3d1ICg/X3vDjnSKu1KpDnkDDR/27d
xkVSKm8Dk10auIaumagGBaO9fKbAxRpZTu0ZtamKl3LCJOov1o7SK1iLp2aPasr64GSJlLHNw/tR
4v9fgMCxhaDVZpGOXyVVFF4Hz4cb0WEVJP8qyu/wwnfWzLsaSSdKJVu1VbuhyMYOhYNTcxUihSnn
avkw9i76GCz43ek1bfLjzksNwJp5ceJc6UwJosPYqZpi/vYCZ23A/x+PC3VqLRwXQciOK5LNre7P
b48MnLMRvua2N9DdxjWwVRZB12VCx7UZZ5W9TZ5dRb1thsg70rJt4ELlKxSWJtMEX+w6cc2TBYkq
9m8ND5vakJGfoBhH/txoKLxqqMYsY3zavKlXixTSJXvrH7A82cmdTE5dCRXfXHqwbuEUJsoD/vLv
mtYK8f6YMdQZR92AXJh2g4bkFIFnm/E2xaarOGXdwg0aDMEN2yvBQUIppLkM811RlYZwwck86r5Y
7ZPC8Kjmwh6mAcxcbGtFLKbo0igUkokOniQVV413Cd4RFox4OZMrpkfa+4dnxrsF81GVvtvETpDQ
ywW0mB4lMbG+dzeAlUnd7GIPeYeFz0832UZ4vRWWKktQXqs/e9hLCTxE+3BK9tncKEfadxA4lse2
e/HwO90HUWQFaBKK6q2lL8czJdY8du8r5YaqDP3MvcPmMLg++7qjwqyk3cWiowkPdJtqsyaRnETX
AD5Hlejc8dna+LF2IaIcKOs1qi4WC/7Su1+wJEgrO88m4I8nfP0CGgi7iM13dczQd0rYLS92xos9
s1YOqOd6HjYsLwe0GUW2e9gAgOTI2QVQI76t+jJLaNs/2G1VKla8gSJFpvVDvJbxjQvKdVp+g16M
BoyMvWFRHQ+coAYc4vwNJCy59z+TdejFC8X7J59/3yj2UGQBiBXGcM8/Dz6KW1TfM/9kzbxSjfhk
J+zIKIFPCgOI6cJCbGsRIQxCnEM4ZHItkVytbauKm5n+XFOmvKiFbif6mQgFEjRzbQ8g8vsaKeFI
lxJ5juaeWRrL2hBPfttUHDaY7iDpVkd/XH4wvm6ifdbQz7sVbGPO7/ASunBayQmiYupkokPtFvGz
u0+Iez8VbJO4XFeWjLzTeSPpI1WKALJSP29TogHbZoTqpB0kqUFUwvBLHTLizXIB+03zrBN3R+Rw
/4kyydoWdYe4kCn8z7r7d+zSKdrO/tQcpLG2QJ6sCCRNR1sAPQSx3uGH2xSMRBQ0whfX6Xui7l0i
ZdH/8rcenhQglH1dhZo2/rQUrCWkNtnalHtpA843d0DQuXswSxvc2w6t4jtvOzpe28p3YyUvofqM
Jv0XMM6sRQz8nn6SZAAEs0nVgEG5Veex1rL0twUc1ryZp17ErB+/iLKZv+8VW7F+zzajZCJzFazg
dUTUfasKReFVDzHvfdzS5pCOMLMC9z7z/uJpRCFihAnvPFpJGa5QtzVRvumKMARG2LMZBjzEY40k
h9AyIqlcFSmoCsLN5izOVte8XoVrEkdHg+Y7q48GmVWL1VKOk1zQy/WvbKJ3l4/vDW5rhu6U3qFs
IVxYzLNXjgkfepGwqJB8AJBYCBKH3dCm4of5IU+/8mtKvHAB1WS61YIAQKTrUA6PhKpNTz3lTEKy
hzV7sH/ArMiI1jM1sq/xxChm90j1SxKJaPEa6iR+XamglUPks9xP4U8efoXhDwgkhQQqPURzj2bF
P/RtoLn4VDDlWtVUV2rjBGDZYT7HjN/76T16ypeiVwNAQXnVxIAg90QwbQYAzRjeewAdBz1clueL
Hlb/FJDty5+NaIRvBEFit4WMNPlZLd+uoys0ZmgoR9+LytFI01CbRSsQksfI0MQ/gx9TRrQA0WV4
HXluFbhNjFGICL1dlcdV+ShJ/Zyzs65cYi+/L/656G4rjr97BpSybOi2mjjInZF9rTN8zqxbyq5I
7osftjp+NQTi9UPi9NRSuPh//5W03JkmRXiHc1MgVrCACVnlUzf1lWRW4mTEqhIRha+K+QyKaXgx
Q4JbB8GuK88n/jOMBEq5iV3Lk7Jadeq0HgMx49+KWMda65dJgOEGksnb2Og+zq9y6BDZav2AIye1
11TfMs78nSZAhi2eyqfLGwNXmicGr8twWAYdVnf68pTGhgXfym+6rR2hDVxvvULuenrfizueKkU1
RYBMD+nQIQ2hbff0ONGKQTYa1AiwAe84LrQpf/IgwoXmhtNozLR5h5dQzLtMEtYX2bGhNyqWXK6k
qH779cQwjXYKLnDCdIhEcQUaIR3EbvCaFNx1nGaHN7QJhMu1Bye1eCVVQ9yDahu195dg0wy1/t8i
8QsBBegygInPobbMSizq7znacCgPWywFn+PJ/L+wcb+xO6KDnVpnFuHPxwEWxu6N4vI4DBmZcwGI
JnDKT9NymhUuy/Eu50UBxRe5EjRXoRtzi/je1ZIaUKnGy5ndFv4xtlSOmDdUxwnXavfObwK9Kutt
Glnxor+QX8Nk7HYuCz40nTwKZb+uqXU7x0SBSGEjP7yipeRflqYZ5kLRCgBYqMYAXXuwMVU9/s9o
bhgw6qgitkeViEG4XMUEf1Yjg++lhdsels+pmx24TiWgZAaDh6w39o5soaGWxlFy35ipnrNR1jEm
Ir8tV7qomSoUiV+U9l1i+HTSBEi9AWZXgKNUUJmjsDdZN4AN8WTAm6xPoG+l7lbbiw3APORPrDKk
kHaOrsnl0ZmXTtB2vZi25MnYx0WZEH6MeVe8y1Y5MlorGe2Nc+j4tl15OU0tWNIk2cFE0C8g3CYX
vPuDlioQJS9cfYM7R7Emsk3mi9bc+h8aIKKe0OOIOYQcXdsgC8ECs7YCTbHixEPIuchDkKRLhb2z
WZXYLg6GENzP0ZV8hvzChnlz1XYdcu01VMvvv+EcXgtSM1C1R1oW1QTpkfU/UYrH047YZapHWwZy
bC7HuvsWDrz439XnEA4afZ1qiva91YzclYvqKnnLBHu1oD8GZt72gOg8tncuxgqOSyxjOJf03lAq
NfUB1E3FY7Q3hzAoh9r9Bpi6xXlXImp62AUxeOsSC8sSO/jynN4UdSJrLOogtnoe7A5P/wSlg7Hm
zPa/Pbq5jtbIYMaoh+hIrSYwxnwoofvaRaHgwgL26Tb4LhgFbHSuUCDOps3SuY8QYjq9pp5dZf0R
xiQ/3AqgYs1crJ25NgBUNrps9b23X97EatRAdfcFXFNjRK7QmMeTaRmXHemLSXZCPfaF8eZoy+tW
hqMA2NuhD4efmPgYaTv57b5MJSiKL45+/GDCU5FeoEAiq19mf9/GMZwFdLnlCEnlNmS1wPY0W/76
7KptiAxK46hOBUJY2oKAzz0yqIGKVViWk6Th/bOHpVk9bMYDXO4pFMws0RgiLTT43uuLd73rzyRb
oR2gBWUyB7HEo6mh2m2kS1jg3h1j95ZB2GQFNj/UWSo3olX7o6G+yEIRdVZ02+UT0qSVyUyQ6Oj6
EUZ5xRwOG90mOy8oLPERv6ZuSBrVlM31Bfzp8iz0z2EjANWx23q6lJwiymwDJG0ohFtOhiYgY14T
WhgvRC0s2sq1EDpiGmL1sc0rYauL+31T3+eEZP95gj+SbyB4DAledoW8jxAh6UqA+XaA5lHf3UXH
duSHComBlsCLvLPS7DCRxQN0nKnGBpp7P7O8tdnz047bN8wLaXNVrExQbCLwpZGwaGeiYxZFFs2+
9SG3WxkgtxaAWys3hpoQ9fSgb5+bFtZAUVTIaG5lAXQxa7WAevcu/37kWooy6wZYBMnppdHV/W2k
x/00ozyrqFWONat4ZNKVgfRgEAgx5yC/C1bATw9dCONUfGeJ+2Tw4VXoNEqu49caXhMVX2QweGBx
UUf7rCoyfS2K4f9xu1vOTC7XbKSV25cOYTDJwdkgDNv8MjrdOuvcHd0iXE9qf7dbSfgOg8hLgf1v
Npi2P8R3EpeQJcoJxzN8CvmJJU4cuvCDGyULkGDGGSgRPOMr4u5dbxxAs6Cj0j6A81EihKTcy6H/
K2MjkC59h0t6wvqWl8hPGbpJjg2oPn5aepp2tGUbHYgz2NRUOm9ULaJtadAKwFXLXILzqqrAC/wU
+hPZahAvOvcP8WEjgCAAYP7KwaVOp5wE0oJCNpHcTqH68Oi+Eol9NXIv3AKbt7TeTMUbbefj9Hxj
Uxv5WwTEI3/7HACGyDl0RXcY1zILp72BBpM+pNpAGJeHjST5sxK17A4VOlkiHYU046Im3WBbodwi
LA+HEnnRftMuNnpDGmUwtQH/j3w14HNYuEQ7Lz2H87q+1YF8cJdh51H0V+L1mBN2xsTXydR4erh8
uzDyhRHuIf6IW/Yf5R6Ke16DgK0M7BScOkeeq9VZaIU9yLa14ea/Nag67gbHGioJKG/FmVPOSUT9
kUduoFCzJES05U8tLgDJp9qJ1fvEYI9PfoYQgff0bJcCT8nbLSgFZvVUU4a0jNnFc7ftxJEr3Cx3
wne9TXcilFqBT8Jk/7jAPB8O5pOyUKjAmoqdPTQOCdEtDdalS4jRacZ457TX56Izzc1PAzVC+LfL
5eYPz0LCmya6DJ3pHxPEv37q7ds64Rv5ejsjPDltU5aljw0Ihv70qFqYGIpnkdcEcI90fCNcbSXQ
4yJDj0BJjcrUoEwdr9hwdbB1525iP8YQtb4e/Hn4Ff/ZTJMqIWSRqP1v+4yGMifp/9oXwPCQ+NE0
napxr/hLZbbuQaeMGnUDLGw2rw3d7V7Re4v3Nd64zeNreKATLlE3kb40oWXrbDgixtm3JlNSwHf7
Rx1ndxeZtR3OEra9KYQiS3oM8Otfau9Ow0evtaETeapeXpU95ffBrnuaGDEp/kqU119LxKIR23Ki
izyALpIqfyKRiIrvRp1XKthi8RVmwurle+HpzKZV5Ui1oUA+FtC60f0TSOlBODA0qzInkeMIrfGV
R1cn7fyXRqoJTrgG6VuYfyb0wsr7Pg/+3Wx2pCy+iLLlF14rYFQSosI7gGtVhUhxSI80Dlbf5of+
9UmP8rKbyi0E4qBIws+OU5wfKExKi5E4qGlPrPQ4HkRVDb+f0u2FqK0r84qY5LeXH3I13UNlI9Lp
xv5Zy8zB4AU0jVruPIF8zUo6figF3hoWvMcvMM22C40/7PX7f59JnoxjVKq9i0aYCw6Q64Tqftlh
uakk2qS9SwQHbiw1sRFQWPmp3PX9iE/iVJ7dYt+RLADJgjF3kh2Uqg5zRMME0hFeMnTjZ49YjhvW
DYgv/oRCNNFCrZ+3KuvcBt4e6qG+C+tnV/q56siYRR+U+JMa8+CrBZCHRa1nAjwakLL2gz3HaVYC
rbgTM0Cmak5hFW5d4X2Sc/rv5sc5QNeX5ytORvmOYde1fi41AkvUceg0woSwqbqTlbZoeTmPqx4U
zVIUln/y8hb0GT0n/BFE/R9bI4BPbJLeO6tvm0xCkAN+4lBfV/SHY4lmt+3+wngi++lMLYjumEJK
3YVJ6ym9shsCWfITvaO4ShVn8mnpBvlwnRNNjvwTxLQIUQ+ORgfGMzNd/vozuQwm1+h6co2+HbHb
+7DbA1rl8qWJymxb67nqa+RXV2fQzj1dNrLqTCYdLLu0MyrakeLYyfwgBvDmv/zZZ3XUr9BL4zd2
bU77nAlNHsHJr5EWUgodkOXPSADaV+x2+j1El4X/HofMWzywQqw0iE4jwHS2h8FkCFv0OJtYgSqF
8+pQIk7yXQ28cDr1EfGZ8fhqgm0MNamK49eKXO0ROmjqsQw/dB1gJXnD9vfaUO8xquwmFhfy/Uxl
AcXvW95/bp+Be4nuz+Uqyn9CVz87drAfP0f9WaX0Oiat0EUaW1aVBfCxRbhZFjkJebx+F0NytYhx
2U4PHZn1uijSh4DR+AJF+FHKqp/YAPs5aU/XEU+CdOcBiqFyTSS2LY6rO+FfS3i0y9culKdHBv97
Sx7xbLhakbId9UtlJajcJ+VgMjjWzbQkk6F8ivSM2x/FVYe3l5Fmz5m83xhppVB/n+rdaDGYexm1
lRGfWoif3lZNPhTkQJy7NGIzU16IlEejiN3Zf7ykaLv/aMegVO2tlLg+JjAkt2HhrTT8vd9FCRab
AZi1r8vEyLdm/DdeWU+kByY/d+CJ4LW2hXGxRLXritUR96NtCnod41g8/Xd4Oh31153yoXRebmF3
ca4y653qvy35IzMteA/CB3SF9fBX6gf5Snk5VO6xwDc9bRFM56g3ZV/ihSu0fDWj6/NMdXsAdVfN
dfxpniMCM2H2jbVeA/PTyDiqQRI4kn60Mabhs0KzGeJHKOnB7GYgUz23QIA2/F29+y/wHYRqKEoF
t37LH3E6BTnoKErLiGrFgBvXz1lvXrNSekMkq4pUfqvUF+3Rfy1KMuemBYpbMFFqSdNBgfMa67iP
bTtQnilLpJvm55efqfYht2ZMZdP+tfjZ31gZCJQg4ojjRyigLrI57xXOzgZmR9Sr9yKmapxRIbeF
N6JaBabupeY/LBJ8X8lpIUAXVM3GE1dmsx+LOqbBSQWFyJF6bYOce38JP4N4zJ1P87DHw2y6F06t
MkV9YiBFm2RbHG89fb3wi3nPIbbNYn5FxW2iSwWFW702DT5y4rSsvQmkys1FN1be/c/2SXpZO6MR
rBc2SR306lTenDr9zCYHWLEkvjTARXi5p3XYhW4CUz7YGhtQMUFwMRSuZGLQST5sYfe6BAJdf+eg
VF03YI/TF3iqwzOJIIzdBTi7evzYMLiINuR4sAuOx7WMm3R68MBfe0J/gD33YVWnaDWV/+D9Rt9F
/yeJOTF2ua+4mEGKsgXFfac2oH0Jotm1HagnrRjZtbS5gUjCYYTLDweIHmjN+xYrFnCp9zElVzse
USPbDSCf5AnD4Qbl6eTgtJ3hrzdoRgtAcAtDaFMioIt5eCWLR8y2Pqt16EXI0lfa8d5/kiNJLFY3
oxwZ66hifBn+5DS97fygruxw+VAnSxLADB+7ZGI1dXqMWX1QJwyV4JxZQODwAqLkftf2CWdMP3i7
V/3dq8JtkGY0FJlJLxWV7MgsMKHe8K2U283SELzAbOIvkrQrCKTJxC0IfuEizm2H1N6+nz6Osx9s
F/ct7VdJ1HNcqW9wenPLuNDkuW4R/bl24rdyctw/N0OoSn+mb7nNpmxinRRJmO5CJE/6aKs9LN5t
tOG9Y8XvOl9yiQQ19jIZ9emCzM22kv5w4dvbEdbp3S9bI6cyUl3ym4kwYIq8fcx1tPDYIho0MePz
aJ91W7es4ZGGH7LKH9QCLy4E7h524Y9JVTiWoHkB91QRA+e/8HFWApB2DGNDGHaHlIsgeRuxQUW1
E+MLSIJ9OlTdKOeGMci6h9kevLHjUYvZArkH6qEaQ+9U+S4So0fpxg0p6VQkqaoF0kuvDc1VChvc
9YZeYNh1Kf+NqbXKyd/bywRdieTt7j8BdvXzD5f0XjXGh7slgzPZvwVJZaG0ehAx0wc1v22xTBqv
GQ2NHwNZCyn0G0QteO3oF1oTdRrHh/D/NwwyosAC8d5RdJptWYxMvj/G9kV16RtbLdhtLd3PVDu9
oXGr0eUZ3uWi65cVYNVbi15Mt5RW6fG1MhKqq+LeKeC6c0/EaghMNL/+EUpIBD998ueoobT9QLLJ
GUac5W4rcFAtksR156cyjuxTda8hD9jP/VqXOPysq67r98EFPTG8PKKxQpye0ZvIkpmwL+0IWEFR
sDLIIwSjeDlGJZLXuLb/wqVOhzrKb7x+l9JzWv2Int4oEb69MjtW0cLCbKfxGblnDOsc7ZBAMUg2
ZcQveEasV3k1uBBfNZqP7OlaQYUtM83whIaY9PuKS5Zifb036Sxk+Eu3hYzxRdCF0LVJWQzkFO9c
TNPlJzwfx3tsRDVDjN8XNJNADJ9Zs7yinlrDr1IjeMIp9VuibeL4blQoDyF2q52F7O6fnEBDUisQ
lm+VFpInUJ6cu/nZy9bhTWRj5Tyf+Wl4Itx7DFA059WbJ49jLZmernhm9x6WAe6+EKiHE7pqKX/D
MyD5Mk8Nk9zKIWUhRjbH+PmTH2JjrPpBAwSXGiEIVed0qmP7IihVswAxKlzlamfo9NZmwO5UoPZA
N83uaWI5HTrHG3wm0pL0PX51inHw2jQzBzSzs3fQxw412WaFxRuQ0IB9Bjmon5uNTeicjTLajf5O
H3ggmr8Jem4azsVV17sTvvEXft7Qu+nRGIykHK4Eaoyc1aS2aQEPp8e/NSaLlt6cNP+2D+8Uk9R6
jxSWrhzV74NwGXK5wMY5OcigL6JCl0FGasjZr1xgey5rcrXg+lGGJZQj2dvmZNbKN5erxD9Y24V4
svBTPXlJcVDhaX3E0xsggMVrLkc3FYGwFmnQGyYywkn6s+62pLF2GmfvkF6t8djWzpXRMMUkbfqz
fcsw0QwJG7pcq0fFt5ef5cF6mzuIwJJXrSTj53/spGULq/M5gtlPmYIclfmygvq/9Qey8ndWAQf/
pbxcpk/UYttT+V0jwHg5+Y9Buop0/D7FBQZ7W+PMgsqK5cDBH1OwKmjHv3NG/n3ULUXxNu5MLm/9
EtnEOF8zAM1rU79BQHXlPfa675qxDY6HOm1Arx8Lgmyi68mi0dwNCaP9M8SBgJ3ZKDB8sSS4+r9j
8ag9CrGuayDRerToIexVyDiOPPaIllBxf1KCSmaDdg59wlnNDUu0xWEbqusBdzB7AZpFCS6/JVFF
hlUpBoAJomdoK7pNf5ZQLJlmrYTYp3+cF4Cn4cio1plPG2hNZRVN5pnuEva8Yf7UMrNR1Ii0uUqe
5Wal0Fogi7TtBOHYmNoomRdJ14D+v5Mg+Eu0ubQav4eRHeueJkMaGTWe6jqz/d6fwnomsszDQRfQ
2s0Ua5ziPrvVq3NVmcLfpLgVN5fEOsJ2FVyKTkN/26wczfeu+W7AjeQpmm2KNMZqkuLCxx99vbDB
He+0CimTvaUQX6/TBacHGIUrdARhOxZMOBAYGT0CL8CpC1cPa7g/87arLtULKFI3qQGrUea5J706
50QO4sJPrmHPfhgvgS6m499m1Y9oOMTercQYeIfxnIJwrCI4ScDSAN3psSGccDOoSAjq0nw41lgK
iVyJt7tLP4IbTOk2lItRs4ek8QsW+vTZno8oAnce5QKDAGd7mBxljDVkQ68l2Lyb3CZFVqOsqk9/
R0lUF4h3J/ut+zPRTSsgJLY5gEWzOAFle5tcxVanjLZ4h4o+itaEn6KkQExmSx+IL6IBHeicS0m2
O3YBdG5x8MEuEnXRgxPTAX01mirGD6pSpILBc/MipuhjeMx8lYrpZDsxMMPTnrXSwGlJrdNtuesZ
ZkM/VnGg+AxmLz2/S/mUgHcZj7RilrUKiwHaIsc03wtZj7PD4diTZod6ltoKgnk3n8z7o362ctPj
1aPKlOyYUtUSAxwbLN/hBZvTxfPWOJPUpuu695a5DRD2e5e1L6TDEl5EPWE08TK7PRuzPlQ4KebE
7kBXfSADmgdVwGqeRbOkJTWjfJrKHCYSk32Y4COfwZT3iztewu8SoCirybpPXKghcviCkZQAIoIH
RkRDZs0NUy6lB5YK1SOd1CXNhUwBiOXP6XLYfzUI0L9XKuHRyAUyiBcsVK8Kr+2NZOWyJmc90Qh1
u9PzO4EpbRKCnp1U2pcWHX8IL2iXiQJly4UW+v7JTRTBxdhhM9k48n8OZgILd9TTfbXpEtg0DXND
pA2QWNRmpLLT+mp/5gn6CzmLVKeeFdgoYv7wNVaejF4qFA+CbhSVhY1Q+MzyoXKu+KXDwhZA74yT
WYAzVO7nP+blMa0GIXJT2R/UbyFfrb8JXWBb80xDZk8CQJ5XtAUSTjf5n0EYVi6/BwaMxCNi9kk9
SkaHMwC+9vPOoDz3TuKZLVuIWphveB+ed1GPwhUgVJ8eOy7Pe6yjo+EsFjiTc5+DEbTYkqGSr2hH
RNcNZBVtB6bsEJ7AQyS+O8cmwqw2QBXJrJdwqOF1klZtTxGsxpuTHv8bP4BUKZAh16fhNOya7u5H
A/e4mY7JvpDF4xGDeF/rq+mlqyZhrM0SH1JLRE66DBnZJD08T6O76xSEod3QuKr0MzEcHnWCC2ib
iQ8dpvf2Rd/eNQnVWMSoH1Iuqe84j2KoJ2yt3HuVFkhAUT4sw95s1cTmhLgrVXJsJJIMOcvdHwhe
fZbW89zDaHDE/alZPsbJG2DkD30K1fSSinfTTU0jo6LP9oDt4e03BtuRgEJ0zc7LFBg9JYfpJ2kY
PCDRNZXuOfsZXxbggO8DhMsNV/jJfCb4nM5PLVZX4K+K2UxlpUn+DR/05MH8J27yH2Yh21EAhh3Y
VHyA6jaRlWE2HcoSHe2ScTBKvoMFCEQmdq2+OcUv/Fo3Vgygs0qQc8S38h/ierZwhCL1O9SeY5sn
QceT/fEUzbOvXkjrNL+WehmE+ICX4DUgHwla4BWWPQH2CELycpIRO2ie0TB3ZX7LUXGYjJ7LehHi
6zjWz2WmAWmhvhawwFardhJZEroWa3Y3F944fDxiOAVOafoc6kt33V4d1vhh9PqdWG3eK6VcVDD0
BxNIO2n4AcPy49LF+C/7ExkxZyqP3Xdwj+M8QIIzIMdXtHwRue0q00vDWeCyF88h7PWQ+QtPGz5U
yJdRYyLy7B45zaRaFcyuDsw6EaugLQN2XMy5IYwMLASgjoAK1Z4NAJsRC7XPKUu1I+S4mDTxbv2E
726x6N5MO96QBGNHxqV+qd7qRHK8RJKK74iAlTFaNGEjkTKu7rp4EsY1LsV5rGtQotebKBx43WU6
uCkIRELBr7TS+2DMMtksyx/HIudzx76IusA6EfoH32gMDf6Zg+XQmyhnp1ihYZdDDk65sboHUBfx
ixIjKQOXew5J8VKiIFkv79IYTfxG1LCHeIGWWa4ggKqyJlWNQCW5QiZIuKsjeRkUJQkEK9s3UYVA
Hibsb3jJY+xGRwScTyfwqhUv78vUgD4DxujWze1Um5jUUKws0KJhUJrer9C8PrSoT81moieVYKxR
TIWAs4M0cXfBWJms3NXdx4gHzh2H2fRQlq5rFh72OtsLgRWLHfi1QJ6rHe+s37XLk0tTCxwDKnKB
4kUkL5IykyZN1zQiiUK4DSk1lrzD1aVGuCSoUOvtqN+/TRnSItU7JbVuQ+HkCq+4SBYujOB3X8OU
89JahdNUQ+b2lzhIyo2lSHdPnPADMdmAQkqTfWdNpcGOQjew46x/CHij450VncIYd2GGrndZQSeb
MJ8ZBMJRCp5/gBqZXalJVshTwzqShHQ1FfdGtMCuoVmccfB6x11qouk8zCDqD0laru9fNyh7zROY
BFXQGfFZe9YQ8iSHBckt0iS37I4mxSAruiGD6d0IQuOIa5dmz/QwafwmJlvgiAguMXg+bCEtjXSi
0LT3j8qsAcJNzuZFY6ksQ028mlst1IGrHIkCjkUjBTLah187KQ26jyIgAldvFH1gNov/UgEzOGMS
ITOMfCYvp9ds4oSTjkvDWKfa8o/GedD8ZT8pYXnqwcodzNerfuAfRDZ/bzdG9csSdVn/wHwOsvt6
yZ0ANfSjUTJiO97HaV1aU0LxSodlCwbIQXxZFkvORimACF1SG4UNwAd2uGdoCBEaMVbDQGW4mpI2
QOS3nnotfIoV+LYDdsd8sqshoZZuEEPUR2D+xCzPPYITFkIrCo1ngVlyHeZM+A4/RoNNS76GhaYs
EAlT7qVdG1Aa4FshsNJayfM85pQC+LrWFzbLgYwgsmCUZHGWeBC3IjYP0iFZiwm/qXIbCpb7pBmm
mYZskr4qMHvWBDGX1fCnOsfOW8lstiE37nYRfpEzJUfoZQS73OR56tvkGztieefe5hKEZbjSfbvn
5h/ws0Hq5/0YZdBOCNiQ0sYZflcbOv4Gj5GGKLWg8a37oCgzepiVqjDnxClc3kZEfeuZJJtR5ACJ
CmyGnQ9lM/WUDYlpbLbsE0JCD1meWxYjunvPRmmVgUBLaIOmxITUzMFzQBEswtWIBzG9s/SX8WfF
s9cfdv50eT9A/31U5U5wG9LNqzPZIXkNoM2NjFz564JoVE2V4C3r/FHCG6SoQpIue7AGqsMHC4gB
XxY3yw2eCif+OORzV19h+qxCFYqDkVFp8G6HW8dBC6oCNJX6aQq/nv/x4J/UbrPfgYnhYA1pOx8k
NbjMiqAkLK/M7ha66IWsTbgG07j5whmVIvfw6v83cbfx8LqkUns5jhfsVc4XNg9Tl1vt6HKzG5nD
J9ZPaCyUSI0308ypWCXXLThEoZlkAdmgBxzrfBEzxw/1+dsre4oqCKgB1qyDAVTHj/QjcRNHyAzf
xhbm8PK06BAPIdK1nyypD2h+5JsmYqAmynxl8gGthm6j4nB7dC9xEEk8pGj+I8aNmqRxr19YCdf6
aVLA/blKc/x5a6p3R8JWvVkfxO4rOCCPVKbKjI7jawmKiTrITB1ExH8a55mjysXEFmCmbSi/Yyik
WjOFzbI+s2rs+AHm7f/hp01NCjZYiSo87tOR0eRAkvPGS9y6rcCzh9VIKo1zZMCtsrfplTsVxK//
IzzbaRnqenAFl6496MXzX/TcFSQ9QrkXFbDvVJwB5g1Y59tPSio7twMPM/QD8jfICCsxbKJzIcFw
jUg9/O0s6pof7eRGlAqCIuWTl54ohUFPFuDvxGbSF0YT2jbuzX0ItDKXKvH96GO2o8dsPL5uXhIz
bMkvibHWGME6YVra20OAed4EIDVDhNNIFh3uLiDTYxzt5YToLfCHevB7AUtmniWUJBrHNODS595z
H3EZKnxx2VCZE10Vhl2Oj8EqiaH+qRNWr6Wf1ytufPGrRebaqo0yrYGJ8MWLrrsv2GiZg5p/vJoM
RXuDjZsShf8TwF2FXlhwqamvZvKcGuAca5Y1nl5wLp5lKYuahWmynm8XR+QITiI4LsOk1RL98E1t
GIkW2C30GMxxHWJTBc5CKtQaEh47wC4rs8gUWwyK2XLRZrtqhG0SxX+5TBQsKpDW+TaGAO4C0BON
muNylLfiQyh+xn5TsAg4DwmW9p7h98Hj5dt+T73zApUM3JbXvX5xqYC8yWp+XOU0nO6/bsLPCgeR
L4Bq0Xkqpro1p61ewSr6pt6h2DUVjI6RYHJMEZvUUDsimrq9wIeT/WWo49Kzet+tpLApJ5kmESMV
Mn0V4MSux/NTB75EDGgGw3Ftp9418hEL1R3SK0y4BK1zvrK4iWiwLoNMstlx78enD6WATLVJle5h
BV3r6MyWg1y2K4ZI2fcRl2im7OWQwMJXFMGoW4HjfuqHF/Kb1GQAhwGGWm72he8BXUB9PZ7OLSwa
iWjmo/BGF+N4UZ2/JSx2HDFnaLu79UXa8guIxkh6Ur9tbJKmk37DiAV0hZF0TX7Nz2uqr6Y5Mp7c
R7qEF1H7/Hv3thSZTdhFqKJLHErg1A3jhQlr88nDMUVSu7GPUtOTBvG+Z8sVTpjjwCMRiHe8dKTc
UseAeL21scOyu+sCla7LON4bP2dxhqfVnuFph60NnJXBOJ5EK9ci8jaBK+xC3CWax/+AtcBC0b1x
UqS1t1RTUQ27iq1KJnORqwFcQFIoiGCmeOg+kNEof7hTOXu+OEMGDALKY00Zm9AMpPOgN1hKxbhH
H1X6AycFaEfdOh/Q/7WSxjVNrdybYn/3rjcHe6m3PAX9dT6RPODWjfjRDr84vFEJ6Y1YtT+JT+ZF
3LA2YpVAgEgvxka2N9mp59mvEXMsYo1MW6HpyefIYOZT/AJcpaG7KOuReDxL/A2bLzKuij1uwpsX
oxksXr55W1C4T3xmNat4Got3C3rX7isljMSP9rZxAOgyk0OhLFSrZTXHWuYn1rmVfSYGq7A7ptvh
5YlNIvEfkY06crHwvziOEfHDJUox1JWcuNFTIDjpQFItusKu4TcvQZRAc/erpRlPQqBAnLRHQDKC
44DJrLPP7RfHa5zK3l6GBxgzfGdTT7i+Obwf/ctpXRsVTuBESwZk+XjhNZQ79WGZK8A7ID6WHn3n
N/hgmA3nnXq5aS/k3md7uEWpg6CFFbI0zkjuJzgm/XoCLCAIVbN7J6jXPFJs9W5tV6q5SPMIM2gp
EauGZxgRsFYEn8uYz5nWEFOO9VuZymq3oIVKqQB6WzH5nq5PH0CNRUYReMpmY51RDG3QLqCAeN3w
i1luQtG1QCeE4Hp0Epg0w6ETsYj57bmi/mW7hdhbUvC/k/6FIHMD56hktbHwVcVt4h0dLDhPbJnk
8dllIjeIV3DPVs60lI2iiBWZ/b472NHRGsY2BL7KK0X+Hh/pm4HAPC8d9BvVCz6mb/6RtLnoK5KH
VhsHFbfoji6fLeahmk66VTO8l1lk+OFxSLgOq24tg4ujYL5UvkSsmRfI1oXLB+KLcVyiyHmxh9Bd
zOxMByaSfiG9o7fqN40zxD7uJVhWgAbsV9/bPu85T+A+lcBEE4B+mFZ7vbev0CGRA+cKzEAgC/bA
88rVpseWjuysWIy6Jig98uaSls8QaqjKFGbxStXLDcEw2EcVALLN3mWqQosFXB+5FT9CekL1c5ye
VrmBg6olijdERSzIJu4dobtdZt8R+kCOjOtqu0RXKEnIAgyVaufwRk8z4kCTqXvHGVwltLvfeNjQ
C3+vJ6rJ05XtVDEOxV697fyhdfw1sX7Gc52oVLGdtglQ4Be2XLWEiBvJR++wlz6uqcUiKCejnXuQ
42e7a6BAFuar5n8hqQwyd70wFCAvVyQBuenyPweuJds+0dw7mV4jnalZ2GCY6apB8SNRGb8mtU/C
TRZ1Q7u0LV5DL6VSrrbZ6tkl54gLD4qi3kI8ZQQcPQk9gsCK2PFZCaMv4Iqi8LqR3BfALKn6M1yz
0krdlVeoPHxOxTfsLpx+jyZURC4Zx514XRCRCZhS9kHiDYILpjFpPktTqpfDMWnjBL3MBxn0JPEU
OfuAP93bzHq6sUJn4baGbcpz3IPrqhkkXuGeYOftzTZIxcKafJ/MJ1TSmvJ4ovjen0dOQFHuvP9T
sDIxwTySHgGevn7Fg2MN3TYOLULEk/EtZ0H9T9BWiubCZojGt7TUgUGHi1RwA19r7pgFN9DQP5li
YGwvhXcJNwgflwrOG/7zgEEEI/+9k9Hg0EU+TTn6ad5+2CIGzLgc9QA/2BdqBgpmWSdcW0QEn8EA
5qrcTeYfc01TF/Wa5nj0R2t6PHav6kr27jz7WBJNSTCzfllkSRa37yrNJhyhN6oBsZHpvrEmYt9I
woFRlJPm9jzBOqH9NcAssnWN9AqucWw62xZphwRKCEUmnRXrLC6PzmAihVjhQiZvqhtR6BiAcnN4
V3UKnj7IYqNRRz5vfbevxzT5thblsgwBC6zD4cNlKFiJ6RC63AeHgDKSgVoLo8C4VBNRE1nvy1Jf
YIzsQTj58vRWy2h9ijLUI7EpX6Mr0wmAGDdIytVU4q5NzkbFQ9+EqAmEi08JEobl7dxEuT3lhS2Z
iTgFqHLDVJp4q4MMgJ2Gv10DNLSmybBejgbl/5F5XYZw7fLyZq8RO+RF1WwZDvastTBtxZ496JXd
IRFwX+kGlvaY6TtKgcAipVCcY5sKX5IZ+4e2LA4VP1BvyNjA77mq538KcxBNPJTiVIgXUrm0NBuE
S0ALUErgFNF6kYgZCb5LWQVG2EhalZEze5RbsG3S1HF1kshf2lMVuX8MyAcU6gaDiSv6X1VRuQM+
UrUm/IcqQEE8bC0qjhNI+/+YHIaTKXh/MQT7lA0ICYMVdp25l6zQKPbGOsHFFHpek24dVhsRLRer
RGsVavUCWKTfHnquUKttNggDDcFOeV+IdTyq3UK7tEGXdMpxZmNiDmJqbLdaxDd3ICVfu/oy7gRQ
7L4XG4YsTWV0D511VXTBi9g9DYvr/LHdeJemKm1Acmr5OXnoX5rSYfYembTahBwe/2WtRlduV7fz
+DC5U2XgaS6V0T9Zx7UPUkMVkWQ6NFHQtCsn9sW0xdFSZu7fVvho0d4pKE9ELTgfpJvNOJwtXUdh
Ti0INVNGA7/hlz3y0DCkDxjYFbLX57K0Rm0duHS152F8UflnLzcmTp1JJg+8YAV/VsGLxofBoAV8
/9IsxfmncCmgo3XwKFCwQGqG3AeJ5REAyt2P/OFgKXKud6IAkvLSkcqjC5fCY6vFgEjav8E5gJpI
2U2OzbwVVjnh/pqj3OrfROgQmC0iZp56srB0obP2pExVnJDuHg1HSM+Svv3pcLfBTz/J2MEughaR
94cHEU36UnKYI03qmEiJ2UQTUawNLfnoIFyGdJsGwaV6JzluMM625WxyqVnuGCp9Vp5sfHHpP0IJ
nJZSEdv0SxjuzWXrYDP+b4qm2ddpLTuBUFUfqXNAFosT1SXnWKQCSKrtG7L0aumYaogOv6vmLRAC
Ec/1twgbgPxrstfb1dQ+NZPYJs0SRayfT3ePKE8QVpcCsYNAyzmnXTcgXF/aojmaqlO5JBNaQHR/
0qW4HUremNHPqJBodidY2L82gfI4jBcJ8BQbvqbzFoPDPcmVUdTxWtMEM0s77kS+BxQzNPY46pD0
vbUW1Yl85D66c8Z1ZJ1DEDiWRWdaC04okmsgCh99ctkShXMhOGIVoELiJPJGvU1tyIXLicqrBFWc
xxKSHgbYZ728HgEh5+AAmdIGbEbSQ8x89Km2VZazaB59vDrLLaaQCx3bmB0OiWABI9vGb/Vib4Eb
/x0Mix+43gYjSHMm43/9yB2IG8YLy0jsic9F4SoY5llNMEuPtftYDuYW7p1YVCnYgNR29Xp3Poup
S+wRg84i9aVXtQ7SHhE12MgXZ9mVo5FzctjrTtqHz+5gMIlET76YEgIk1OKmXc9KB3hgnV8Kg+no
SO+3futeNQ+U5GBUfjEfQGGOqL7PaN9MWUaOAVqI1qZiWiD9RFBrcU4goPsUf0wP6Z17IzHWFsdw
Vl9t5H1bmT0vwp5FbVKilFmz+WCVewcrFHWqd7TKaM+qkKFChecmGK93wuJNQfjEe0jDURiwERez
SkDrFJHp6xRlVah7M+y0uOq2ZgD40WIx+3fKXMjsmt5nLLoq4Cdss0vpF7xgZkVcZkbpRLTbW0rL
5Mudn41vDnlP/iPTaIVl15/rf7da7TcHECetnPMnYRXF2Esd734oTctMeJ6s6N1yYBGif0QNzwHp
UCvBiSy2eLrdz+2Du3RrvtZj0OmVRtxqu2KT1QUxjnitJZrRQeooBz6pM64Hio0EcM5UUCxakJ4R
Tyyq7nicMtEOe5YCm/71S8XeX8LT/7jSQ7h8VfMi42SSFa05sW82xBcyqAFCKAECHlwvefMhVU9O
ZJEE/jjLdo77xYC2cRatpMSuGAgu5LKdFYv1aMR50+xergXqrcvvfiULRaB8/OgHkx8ZA9cTeVEl
O4OPu6vReyFq8vbT4x6gHoDNGDwm0934FvP3+Ste8+InnIRLVU8Zv1xrQ50FKAACYIN1uUNSgCqj
tldLRLGB2x4wX39BmDZQeoJDwYqu3wFWEEfNqM9vXkLYVgz32oEdz5l29Lk4sAswhsyNOm/7vYnD
dF5a7vQGKXJYrupKbfJ+3rgSkm22czHSFLu/3t0m7IBx82O0msnedRYf6Kj1Poms074tMuTqK2j4
3WGZUj9R15ud7+FFCG1tgDVMK7qAupWFJrs2n1FcojXkDX70v0p94XH7gi9CWm+hjF+vDhUa2YcL
lUgoJ25FcdV5FYkM5LodqgQpn55E4H9GRa0s6QBu+ROmSZbAdTkAUhKffB8szJY4CWoYLfw6qdiL
9PwEvgOuEqO33QzwVtts4/nwEa9wAEjoa1xyPcRWBxw+a8PPlwQFgGf32gYp0PAzP4pCv1HOwpTS
CUQq+zIg4BsNWei0sf5jj+xztTNwdGfzDwhAn02C6C4mj/uFMT6cOHmBah6r27du7EL5ot5zXzOy
EqZs3/+ljiO2PXS4dKrN5wZMOUxSA0ibdAbkUo259UtPx+HH0dyz30wY+CYgFe0tJnt1MCfyJdp7
EmNA9iHjrKXvVM5oK+mW+MVzckPxxE+TglIZAlueZfmt9d000s50UtTWhpU73hjctyfIV57MQpgH
3X17CcuJH6CXkftuugWyImqanLsvXjeuz0cZpQu4SYA+3Oh4IXyBV4BUp1ScMWYH0th3L5MzsYxc
Zg8+cvuuVQAmFsmBb1Ti4ltLPdPpzPHNYEPWq5tIfh16F8vfWWJI0J/kuXzAGRjfOkaC08TJyRxA
3VUSKaihCw7PPwN/zo1hJdoDlKf6sY6payjVeZtN1plvKgpHbH/VcX2FIGSRG2yU2OPwdStUE55F
Ml2tOUzrA3HjQfmdAi5y8jhFXuil2QRgqgdasX7DE6joRHBRzQmxyPY3G4YA+oRMb23pqn6UyOfb
35V8CxdDQu1PCjOQwuQSZJVjX3o0v5ocHhsCq2zpJRpcSPFDt6hxD7/VvIi0DFTkqj3a8/1YR+CP
PhDbpsy5MtgLh7YOie5ApiIvNE9KRPecmwI71eM81nasI130JRcsBIU1x3hDWfN//hkuVaIbuUJN
2qLp3xTbR4+m18xMbub3wI0uBc2NGodv19iXu8IOJxjFUM1S5kNqSy1UWgCDnckwcptu5yv9SP/p
xyZe+wkKlWieyYVtvX3js6SGB7/bJ1lNoftH7igojw7I9n45K1EsVZMH7UCZ5N51w8IQUqg32mvt
9m0tAZju/WJvAL8bsTCSpQwsPv20t0dTFWIJlSrFrR2ZZcQ1i0Sgl8hQylL/IKuNHWJZ3XqVWnc0
h/6AEz/3IWCMzwBKc/QqZo1QIksEXC9LF4BbC6UtwIGgkd57DSXxFs3JWne8kjdVU9cfXjnEbnA6
EBzV8FRa5Uv2aLOxSAsHhahgR5ukUGlhtFbbNN4wuJLU+I4cSNHR7DZ3obo1Dd4VLBs5LddwrQOz
GDEu7ErqVjKChHbyDxB/1fBSlZIs++IR3hP4i+LOgT8FgEG0nhWgQh+Nx8VU9yh9zxnsDGzEN0ul
dHX0avKadD5+N6KMOotoGjeMKMYR/+a3RhhgtzhhJ4uZi5vCosOHRU0e4z4/RbxMkcJXgdFJL51D
vCAXnD/mC6xBWVCWC2k0GV/N7txTLyzb/MfWcDt00CifCLMKSMzOMPglNrrwKbxiH2APhymI/w7W
h7JdMYpkTJuRhER945dYchAgMRGr8ePyDnN+FqXnU+Aj+wCrA+KV3CVpmR43PAwLnEgGWLWc8cT4
cha/AWhY22wkBpvSHChEwWIm5d0cAAneTRTNiVVbjo424F/mNxObmkGxoQfitjAu36dVAPy2yc/b
xs83QyjA4Tefiex0RjcP+qsTVUQE23VH0pq40xgvO70oQQHwVCz4BGimClEYLfaBZwJhIJqkkKaV
ZLi6ilzMsR/eNUQPK/7BT8eipqexkfWYMBdfWm00/0leF4Biwly5mAKdqRrTsn2rZnvr3YpNwrNd
4GJmN8U1dmPYw6Ja9Ay5/CFl67VIdtDyLnZu+vaPoG0eBZkqgTJWm3IVvS3ghZH+W8OZ4w1TqMEL
rtty3auhboGXNVwSrPZxMXXDZkK3KZX5NCk6YGicDSAXz60h77us3aNVYYfGHneBJop/ndR7PEz+
Sr0fiY1rO9RJC6ChgzUae/nqrHu73+ecxyun6jn6hRgLGIF5QlCTHffewrkFUnrfKvto2AqG/5xp
ngzcYSec2VZVSQqEAmkoDTfrWRQZNOJrPAIT6eJie7hCTZOaKmzhPLfGX0elRjsQ8mTI0APcvVqj
aFq8O9tX1E4tehZr4RXc2zipJV7kv6u7O8llRYW8XUntQEe3x1yg/0J8T2hhAL1nQXHcqJrD+WJM
9BwUvpMK/71ErUKSYlUEcfxAhrrirHD8R9kr7yVs1aEM96eU/X2PhKG7xyh/UxljECa4k+AKNPHf
ejXYjULhfm/R4FIn/ikC3xanFUJpmtAJrinb1oi0pSdlVjIsL2+1VvM1XcqO/NfKWn/zZOd+l9Mj
OjoJ/rVKS/sftyYQatztArzkJnrrXLZGc45WeeRxbWtn6bwNiqdNIT/GT+ye+E2r4yh9G69CxRs+
8cCF/CdjU5/KOLmCAOFfyiL07/0gk4EkAM+gfrJZuK187iFunscDBDzwVWqsk/RgtuPn4I+btbhj
LFFm951h7CiHRZjsn6w1AHQ8M7/+HfOR9CcHftvBEPPQK+gelDxEL1j1nUq1AjIwstazSDtv32Aq
CEOUpqpoXaSFPUxugYD0kF+o8IPZZTS52EeYR8evzW9CjtmPIr+3XiL6nLA8AM8TvJ0xXYj6F3QQ
l70UEXnpm6lkFqfNYOsRRFDpgMKllraCFuqDZv3ifl0ghCBzAwhy+AzAUW3Ys/StF0+bH8wpaKaz
D9MDky7X4QTtrSzDDswjMI4OR/OSqdb1dL00Lhf191HysSY2aYpMqI1gxIt3Py/z+ngRQTiHKUA8
Xe3lY6xls6TLflYhqiGjD8PeETVBxwMUM0p4IgbuE4GN+2JFjt0Z7w8J7Rq95GbkudahQXeD7kHn
LgpJMswy4Ag0sLhfk+c10OeOWJ2uFJI38YoYYvn2/+mV3vJgKUZ0+bWKE+DcqHYSI12USGAJuuN1
APafHqYecaNQBFjfqk7BzOTtmhuGsIotNlHqSrlX13RoNIdgUh8xUDo+JxvU7K+WcrPOoRUq9Vfg
Tk//8uHVA+rBPS6IwLUDuzoUCTjzxmg6zbEeayZ4oI/kkTxxbnA7pwqlGNWv8IbKYf+nUQw+8BSb
O+rNEBg4lNqKDThYx+mdAqD9kMJVImWpzVyFNfloJSAFXxqRj/fhqeDpN+ihQwNzCjLZx6MAB+yF
5bELFnIOfTZicuxsQtkImL2B/LWLR5sZruih/hLdwHMGfrPZpAPkujzlty60R203drxh/wzIif6T
Ky4LFQx6iDbwNz/zjiajkF+vC8ux+ya7Cp5ZQUU7OWQVZpl3BVJEDbcFBwARXpMjK6qyM43lGQQe
70CNnjoz/nJJjtUlaRdbRwXC6h6kQDfCJ6auBwFhIjTCovUTO0xECCqEq2uAKSpT+vW76CKGb9w1
AbkWOzGvemfPTSK/l2i8JBSpdjl3c87ddm+ujrITE9at3eprF2KTS+6Q0Nzr7H1kBJSTNLrD8Xp8
pDU5qD0Igp+6bDG2sXpsubptsqjg3hZ0T4jAzQtisGoU2LSCOCcyxRrBdLzq22mNxCPotAhO+O9+
SB+QTCcZ3vmEX0yed+vs52eXjbaWSgPQAOnV1radr53UWZ8kOH6l5rHsjFE3x6KXTT8c5bF/MfAA
NkaMfTuX90V/CdmFoxIDbpKWlJvAWahqYFflMpGIL5OL97GnESqi+6DRvYUm3ik2nY9g1F3V54Zf
iV147mEuPEB4L5EnolSLcxQy/ojRheNh/Dhny1MVE9fHZZmoNoLp94o+QaFJZ689o9UEtXqVwV8D
c17zD0W8yjJmD0XTo6b4XKVM3xMWBhhEU67L41vqXFY8mmpb0lW8K6cKHfJ7PJau37ElAhT3+qQA
R4quy9/WU5ee/mU41QOQP+leg+MXiwEgQRmaOndGvmPSb9sxh+6gxT0gBYGmGaF8TgAMEpxzCGQG
yeDG8VBqqC+zlJynp4v7BkfDa8OOoAM42Bb/9iJRRME5c3FKG+DGolUJ8Dpb0/ellmwWevdulK5p
X5j2PdBRy9Ce76+YbBbNeT72LRc09K8q0JZend6Wou2em1KIyMyQu7LkbToAPw9du2VXAjm2y5uT
7+mqEMRAwVPhcOx2L5Ioc0vLTBchr3HjSHfOtt6wOrBxZsNneNc7ZYNSVQ+yYm0zovU5bEAQY2Fr
saxfZFNHd8PUwrI/hqOOse699krgOC7NNdtlBzpasTqdSXb+IDebWe5vFRrwiKRb48IntPNnZ1rR
Da+48NyWsF2JgI3Zm5Z1oVQIqLS1fvmbmECxxF+TeDweUqbhwYGT3++2juzaryFQIPmDGKHjGkTc
ndrFX5QLS7soZmxKteGkAu8JrV0rsaK4oBYyodAjQ/95Y7edkUrSD5GJFhugjDGVYfImRV2o2UfK
4gMugKSGaT3IvwP8jq4Tfj3c9q33R2UrbeuFlCI0EvM5nWz/NOeds9DItUiUj90APeUxkfRQqTCe
jTnSOk025I5mB8rX5fnYc81w3u2SEXFUokmEEmL9vzi8UuOrBUtWfRqrfixUWajVXjL8ycB3OOhc
YWc82H9bbv706b24pSvU6Wpa62w14rUM+WgnOOwbEaIuQRwDZLMFaA4AcTHxOgVdMGcTlzKHb9TG
iq9xkTgFFmpU0v2N+kZqKsR2xYre7YVET6mc2ZLIKqobbExDhMWTva6Pl5sZGk2wSRNpbsjyErDu
7RJFRrt+X+fHIr3OFYSvNyMWqBXZySBG94k029PnMJaYj79bDqePjKDmoH4nr6vq4+BymKOoyPKM
3JXe669cmrM7d5wSBrj5xKq52YrV+ZhNjIsHCG7SxeTdze75y9LMrzaU/4LGDxjPnPl2ERTNwGEY
jqg8b6RsnnKebKQzT1JS5qNRqsg2+qy0OrYm7SHbkuagLY/YJXMowcFb/c8Tea+VH2MjZddn3XeC
sZU/ChvXslt6wdmbxrDx/uNfuEbpu9R5hMMWiXZdMPSeIfFSiXre8MFOQaIE5EGUw+Rc6DMdITlb
8fk87GuwOHMRAOftd4DO942Axern3lMWRDf7XxKdPl+idVOQQnbhH6ZPoQo0dfg/jLTssm7aa++t
errUlOH9dWEWO8jmjRBNNzdNCYWj6QJNbhTcYfJl8nxxTuu32RitduM3Ofj1m4xkR4w4NMjxNy0x
NRajfLtuT7VA1utwGV8o58W4aC1S7PTI7CSSUHx5xJnU5krWISOVt2A8eI5Fv9CuHWbGbg1YV8ZE
X6EV5Jq3wi2xTooBfaOYAPcFedQSqOy4cdFZzyaY+6/wM3QbOlmeV7FOGfeE/+v7be3eQ8T6LkbQ
rGY437X6AqICAANKryYlpLvfobJCtZG9DMteUi4PvGTXMwxqZOQoeVFB8M1ZTNiuespPyEHcIahA
wimcaKVg7jDp8deqpqHSASZCQ4fKN4m2NvuxZk730cF90h8s0TI/2315rHU+EqCkUG8a7TkExOqt
BaZMVdI6yQU3VileDB8RLz64o/NZuWhPljFvM1FN1ZNHU12U9vTvShaK5nMR+ImdxUb0e8KN/kdx
u2Og2kzu5f8GNtpztpnsPVeH1t4bqQ2PZuXb9lSGYTC8ke2wBxmivVivNuncSM8F8m68LqpPM7Ql
3xcSM/gCWcKq8DMlBqzpMGoeUfkp1e605aTlpjsmdJPIaLwO0lrCJ8EYtrSkutabU2cG54sfaRUo
nnWFvcFtLCIdvw5C1bqxHII2Hvt3DfZGVP+Oc7aMx53Pj620F7Qyoo4yJ9085iGPe6Rkp7kCL5Po
n5UhTmJPADvpTO6Dii6aKxiULTKISmRfWB4nvg+3UX4JvrNcWF6k1uCISd9IBF/lZZJ5AFUuA2m+
YoZj9PRh5GeSe+ipxJA9/SS3XoHhVnuAZv96BCVZ5JIhdu0kEqai76umJYL2b6jNWPbUCptJdmSd
H3I6i7J0CWbSLVssmtPD97TAyBjF7f/TyBzyRGt0POscq8P7KUOG8r717P8srZzS+WsQVYFfnRu3
Mnd3tDs18jxdxBKaVySsOxzaFczgfV23IWNxfs8tw9aFjy/eKD50b0j7UCwZO9bkKgZAnHNRgwKu
2c2HnWtzcrE+3Ma2Nb2Cghe1GFuriG4NDa2uOG0KPIvjowIjrPaG41K1p5n27kyk9jwvC/enLVBD
LxSORP4LhaDLU+N8hQeNkbu9PaOR9B0pXxw1Z5ouL69NyOtHGobtldi6vUfHdrv/nS6P00mo+qpU
1gND74EsFHPBB7HLvB5KKnWEBmgYnYkn/TSyExgstjTubAvkyS5IUn8euwsuRdqyJEWAGxiKdTGI
pIs31P9sD8EU3gK3JRMOWqHx21/Eu0Kwfww6MfsRu6lRbJCVvPICOhi4xImR6vFt0RrHsmS7+CVZ
jkex7RgAOvgB+gyBPPDhXFOKtPM805BNPfJwHkZ01QbIVOMXy5V9C/gXcuplME7ZhnYFvGhVM5Nm
bD3r0mJUwPDs2F0TT39L1/mJaSvFVYbTpiBR/WJW/Dji4EGIhlm+ZLsPy5jwcZIgT/739UT/5MW4
+XMNmJIeVAnYh6Ta6dLxTNfTGogJbbDqST33zyd6qVd0m4T4ogU28bQXtyHheYC3YMx/CnkdBJGR
P6Rp2tQgFyqBVdoeGcYvfUYQelX2+v+ZiywAmuoaSSZXaAmCEu2rvkL780D3JkSyNC2YHkOQ5HUw
ZBskwc5TjdBvWuMVqlBuRucckP+dJggkOdjUYh41/8cuz6lQETK1vAgugXtP4nR18SEO9BQJlxzD
3e9lYtn5NSQKwx3FlYEIqCvJsHbagAJWMqPMZohcNW2ABvTltalNHvssZ3H1X5qdUKX6y5ksY87n
NzPwOPAUzEfGq98Q3+/fK6t3obuo6UMWdCT2BsKa+WA0hweeOdxsrRoTABiavlojBPpfsr8bSkHM
rFjJ6cVXJYiAReGnaAnEprq6CUqa6Z1pTgOUSVvwRTuxLx984oPygHKDw7bdyvRtbgeew4a9C8P1
P6eUSN8wOjmZtLasUyJKPkE7QmvWArycURqa7ImwJ8fZUxG1m51qqeRwUJ4UVVFPTG/Nx5Fx3+rV
xInqXLPRDFQDsGDgc1K7yZHYy2GP9ru0a5C0VCcDl4BNZEReRvSC17Y37aouVJSJ/4UrOKIgltLq
ChWRsvWH99ayFg0QBUrzXA8LZ2d6fseirCdVfF1BErWxnZfVk38EX7VEvRM+KxKxr5wIsrGE+kuI
zy4ldgDGyrrRZ9MeupufBkPssgwiRUn0e72J6A8a7ajxDehJ8/dugd6oV+3J+/G1MpK7+kt5HaAF
blxdQCtEmIFqMhQP6urLTDrJLjVTqlJ6ZaBXFNAZkYutg9PAMNGN0iZn5NlvPI/yH4d+PDcpOKNn
Y3bsjdUgu6sa/NSXDi5WRpU3y/BNN6UaODFDMIZmixIX4UpLIp7SO066iazEDQvz4mfEYQa+2LOi
m3kZ6yBgm4ktUBVQ9Y+EoxOyqCaW5VkNYZUCAr+C0gDtXFGYpP9lKKJ76DN6vCoiv30x39ugIMcI
ILQpHydjcsAHhmVy5IWvwGEdXrIyhtDlkNRP+OKhYM23IwVodpzSFvmbmYwb12peABFGDk5nsLn6
ZBeGRYZT4WHEOTyuJtk9gHmj/6qwyrpgNlsGKIeiOOZn33Y0tGMZTbkHoke/vyLaUoRhxF8+IpRo
qHOYQtowclE5b1QKxdIaY6Haks55WDC5pXsPlmrFCXvFoaUT6G3fCCryMy5NfNHUKROZyZqvCR05
a3O9p1++F1YmwlhR9747mUP6gfNJ/NupuJCdSah1AlAFAwEVPWeTQKMxIQ+A8GPL0IbYsDWIBaEh
z/csB8KBXVPBQd9zs7Sv7Zjs5YDE2rdkpJvoP1fJI8f4lEorncLeMWaUwivvkoHbuvS/NaESJNBg
4m7tA9K5HeweX+BCIo8uxzvhLRP6cguXBTcMbjdJJ07M/DEZ2nen2Hlg8n+ZTJhSo56pi6s2QJIh
7J5V3eX7naPhBz9xktefvVtFSeGNC/jDmsrMuwO0UOi1maS9Wr3HfW2wgZtzzkwVZJN24/h4VcCt
MFd2/Ks5lDC/5kpXZzBsevYcQUtmZLkCHSa6nz+hyJVrW0pnCjNvov65MgxW4IhGCP4QGZU0T+KQ
0IO0O6lCaRt0EXXgRkH3yCajqytWladKaM3F2shM7LX+467FfWZghp1MCKTpMwQ6C0l6jdVQir5I
G3SCvZDa5shrI9Qj8j1qcrvE67h7vJeaMPvL0ehZefBnkL7Dzw+YeQpfSJw5Ri3wQJlHjAGhCLQX
R0LLnqYzfZq5WD5bOZnYZYn0O280aFGhCQlHwTCelbX3fhmCWa3hcXzcuR/8D39qrof1ir6S0GdT
szZqm3V6CbcBwxqEHJg/Uvs4JGQJgXU3WB+46B51p4eXejAhVJCwKcTg5L1zHD+6MuIMPBAMY5xX
e17S/JjRdPfLqF4ZvCWDy2scZIu7m3zkrHjp9oCAIGOP5pnXiGJxkCYGRFQUS2iLBV4vdZkmfmp5
7tEvIXDBuN1j3LzWSTC5nbrx1rWwQacLp8ojsTGk+jZU4MnuJ5CMKY93zoAtJVdpg8871f17nU0m
fHPIPA9cOoPySFFetIPplddG6FpkL9BGRNuy6+tm1s24xe9XvJf8iwtxfGmnY6qCQDAuexcB8OVf
WMypLvIn4F+Ndekm1b9Qe+pU18BX5ZKrA4kv0rWJYG10ox/slo46HTv2RKuX1WgKZ2mWaF79nh0g
sMYonufyTtBQXnBu/qbsUOdfR8Tc1VsQ+l7zb+yHjFAj5XwqITnloz/p1pizS5BSuuMoJrfMkQBk
I88yKLY0BD4x+6arck+5CbokneS7IrWy+8kg9D5JSRguFhZhd8/Mbgdv+lsENi28DWgeLLmUP12P
eugdZJE33qqnee5Cpc19NEr5jHLX3bor8lT9y50bsmvzLZVSsP+O/8tOShRM+26h3Q9xGlukUXo4
+ae/wSl3wuS17omVKc1iLKiUrZ7ff0ZHVkwLWQpo2aJHl8zn/Cr/ftPj6sMtURQrQjTxJ/i9O2Nr
r4yAhyjML/ZPkwVIzLhiDtQCppAuOhWmZYcgvRbj1SmdoiUVTjmSjhs+I04J0rd+/bPPFFw85zGN
aErH16UF3KIYGAmNNj4GgD7v9sNpc1jQnpdxS8uq1wlEwN71oSfqml4M4LQVN2ejmnrLnamHZ6ed
tmj5MN4iQkAxdH6y4C6SX0ntRoq7TsRypf7rOcZwILkn5i+SXXvseSTMnuhVTOqgVQwxEMRyRFpU
iRw7/+rEkF1CA/PMH4a7R1E+cvOkltxKnmpMliDENvfd0kZgQ9FeOhjOZXan9OPmOZ97SYX7Fl75
rqNhow0iV/gwGrtOSnmCOvs1iCAVFKXy/VfCyd+Mdb2M9EE96r6/vz5UdqUW3B+ZMS24HeJQCYjS
oWJYPfUTiL19Rh1ljr4q84udGy8bseoq5HR/FQnUHjvTRdH4MxvFYVn96MBGQYwTBsKMUpzb7Qlt
7KGs4JY8Gv8lsqjRUzAMwJ2LfB+bEgRDBupxBFIM5zWuZPDDaN6jRVMgbKPdOF4aSN+a4ZmcH2J2
d9/O3Yb7oHbYYdPxqYgzXgcl5gUeUSNbITrRjlM5CtABy9UQ41uaszrEBV7Jd03tV6eFdS0rivW9
QkhrYqa+mBB4Gq2Gab84gJMGlDHbA3JNwsIvdpfIT97IEd3guo3lee6GMw/cjuHIpRYfFqZELQYT
cZC2kcxMPUx45Dhzkg94Vag5i7Qc5UFZSiRlkaNlsfzM/USXsR1Ahnl6X0n8mUv0c3BqmLQ/Xftb
HwRirLZBvCU8YvnhPkD3FTA9eqye5M+Af9/GhO8SxzkdWMd0ov1j0pGJ+M03PFJQevYhg80ag6EL
3Ds5pb7JX7hrj07SI57Irc5XsckKa0HXCyXp5uMmYu7725mZjEo3LgdJmENuinvBAEvCdqYBtWgW
QjSxWKIcoZaH6199lqIxvoxuj4R/VecyxHpfFr9CVJfPBwsovUNOSfH+KUK+UD+V9CLuHYpS84F1
D8J92rOEcByQsQjDG8Q8RC13hchzIbB4TpNRS7iKMRje+K4REenC2duoVXik9oBGXpmEg8YNXJ1Y
Cfoa83jVzzc0MD0rKCsMi0P81Ayi24aPGhsAZRm6xQDzTtFwgrtkLpo9RU/LozN0M2fZCS5JPE8h
UCKl/2Gi/EYh3KCJ6N/hFzQo3wbU3DPAVovteS2fgQiVFr0s7hwZFgHsjEpQLOs9ZPgF0gMAVpyJ
J3iZP3PZ0iqePqPErzpNQJhOdQqqY2An9njOWOZRxw50wmQ/63D6tmCsV5HrU6QMv3hrlmhPYQpa
r0zHtjJI9aNUZeW1fqglB/iALjRim01SVC0cdf/T9aQTITughcCvthjcvTEcPfYlSmHXr0uORURN
7BKA7gkoybcFDg2Mt/dUPuyq7S51RKEl25puqXRE75zORjJo9le2POq5ra+3cuvNHSDlMZBSvOrD
Pwi1o8LcJ6kgm5/NEk7iXYCIKqFqWenK86eu3ljT63kjx5bwghcnnpfJwLdVNHyt9YUBYdaxhw9y
xzCUD2d3kiKayb5fGYixIcq9Ki9+TkZFC8yQ6pprYXWAt0GEouHC2T7Fk7IB2MglXTiA8pVBS72O
ITMZjdOo9bhHmiZ2a8Tqhp5yMrDh9OZ6cF/l5fnPy9ou5qPqSpnndpWSuAY9weQ8gGDhVjG3RaKh
WvswVn8T+n4zjwUKUZGlZ+XM7WawaLKaM/O4pK9AHk9DubNp4L6gaCDrXYCUptPPSoCby5vvOn8o
dyz3FBOvFXefU6FJoKdfgHX0NgsACiASFqH2OfVcTqLew01CrwOcvverTR2Sm6AqbXG2E5fk7Trt
aI2yTZpcrHVssE0+N+4i9wtCejLWuENML4iDs2DZ9sGUYK0vCxH5Y3Sa6IamjrhJSsiVfxXcSnbq
so3xIq2m3/AAa4jSeFQvwElyCyRtjqbFi7EnfLC2TSLQttXgJor4MfFkpIR/sWD/GHpDJ2+WzFwn
WGZVFU+je5TrgSLhM7vFDbczIEwjUdwtQ9nBu+UmzkhOoEV2RDYHbrMiAXYF1MsEEAYJOU89N0Fh
lC8RC+uxTLQkdW54Y4FeDCzaB0gLNWuzVgOQRNdSbcxtNzGe9yuHp9MizSMALmCw1KDZot1/c7bz
H+MJL7jtJ4EThPPzkthusiGdG1vbnsdUIsHhCqPu6J1t9K1vDUQXiobW/o46Ap/FW7NCJaYj+ohJ
mA4RyzcRNSDVeA0eIyZTYrBGQEBI1pPWFYh+iBZo6GKcwgHmCHKpRyM3dPEsuHRX6ep2J2GQ4ja8
uMaAoh1XwhQM0+hKcmYRgCYiGxGIjEUsvypbOb3rE32hWY2ePDu+XHvifcIpfTnbNhVhsoBScaQz
Vu241cfMHNPFNoWTJEL4Z2sicogUL6JlSFJ+W4q09VcOy5yKHaSu/xnIuOEP2tH/osDxqtWFL2MI
cIjzlUyZLMT4p4FiYCsCzscEJe87La1rD1TidiDrx8tHjddjCQpyj5+cEHjQV3GRlZ2PXEswDsMv
SvIl94PSyJ7jHPSVARsYxgTNggq3IWjXf2/T6+igGC8i7GNB3OweB/Z3vM+at+SrujTg0UmR8FlJ
xWagNk1GVk1B56+LlYxXR60dstXH70F1PWLdKXUTAGPdHqp/UN3XmclKN30JY+H6PyxeWgLmzDd/
rjow0u6SBGUXTLdWFYDg254SJnAxn3l8Bm1Wz0i9KwT3YBd//klETEhaxInKzOJn7lp82TgDY0UZ
S6g+1WgfFva/jadIvrnKkk0/742yjGqsVSitng31HEU6WXncxPeVFOzss+6tuOVsf0PepBacegRW
Cwd2s4gVvCczLuP2sekxSfd50HijcLB2jcanciPTAvQpJVgNHVtal2Q32vnMTgE1rbhdC0/q61yV
tpRKQFPG7SUYpmDC3P2sBmdoH85ZKb4TGB4ZKPWOS78bThaQGWbzwkSZAkE/YA4Sn7huzihzYeyF
K7Cih4ujsw7Hr1vw6pDzF17ckX5FDqYuU7W33+fH0I7Xaq3tE4I79ibRm33aM9bfKkkc/b4TQ+uJ
wqUwIAK93lsjAwQF3I0rj4dkolEleTX0/6DHmpiCEkpupLo5a6GqtKxrBO99QwxXVXpwtui/3zhL
tiqs2qRi7OCs3X3uZz8jWupTHGcB7/yqcMJdrI/+5p7TQbPqBn1qJd+Oh5lYFffxTgkX7cgSxrqs
m12VgoAsxZxhJvHRl3A5VnINcjsUObx2kHw1yFpiRQNeB7+TC0cKqyjnpwVhVNPgi7Yh9h83Pxbs
8oqQx9lxl3wadaRJnu5ej4ek5jSUgVegz8UY6HM4fIbo8jk5LQPTQUkCBnKWYLEGQwMYUxOaclM8
HSecRuy9a/ePm1DMcLIoXXnORc+ZP4LEnJ1DSUpYoqtLJ5Yf18aG+LY64ncdEL2WFjBmP8XtGhIK
ZlN0etprgWbXJbAv3M/o/AgkRgttqM0uGOvAqHffhf4hJO1B+HcVXmuLJJus2wTFhO9LAkhqUMJo
xzp32s1ZIlnpqiVvq8jMoeKUo06drPRZ9Yj3IRjG/3MNBWLgMAI4YPYQDgeO+IBj/biczUCb6NHd
WaKdvc8mgAodByyPw2TyFczk6tNWp4LB6dX1Wec9pDUZtzIKVxIxhGappubPE8sD8USKRCXRS51s
4kP+fAYgbSzoRAPa5Zt7ChcC32EwLmuj7Es9gnT88ox415CCxkQfcCKM/aUYK+mPvWKc9J8+inuM
XIwvP7dCYuJlTCeIEmsbeGt+d4f2nAhP7/g/gANgh/lhGtnqvXF9K65/0LfUvdlrkXGAlGEtHXzU
yqBUIvEIjCXJ+IJztTq9b7qWdf4UFtNRvnvDGcG+QHH6aEp43gpD8SJDAm9FJFTKc4TqZjBhiPOy
y4eGKhOQleRr0NGfc0KQNRrGQ718mqq+sPwsms2qA9SVdC65shgzeh6vFiQSeGE0nvFqknlZIPQg
mekQ358xarmtwXs6imnLMpEoyIkwqbGwmOWQ1XRNPcu5Ba3YPFclZGLyc5VBA0TeYhZptjHtdKwc
igxRCFl725C/QpBkBUHIPTMay4TWzOMZBITxEczqC/emUnpRwpXFI3vmdzdAWSBMPm5kJLURLBm3
W9RlzPG/EOlNv8WeqzRXHwEwj7PjHvmLej2USr+/rtrWJCfBkTWFnQLY07sLbM+T7zMnIER1++D2
uzjbQzZZMmIfyv6djiZcMSPGduY6QUPJw1XogimiYHrsg+Sj5/7qTi+pczUn2/SJofgfoKQsumIA
5xQ00yuAAo+KQqtj0vCPoz6M/Z7YzWD75aaTcVphDZ5Jzd+6tIbaCA2EBk77k5/cRXMBVkpeS6gS
XgoFEcIRKBjLvuCAhXtv7mzb6gyCoeFJaIQkvNoOzscDeW5CC0/Xp5QYjB6ZRc4kxfGxeboKzFTS
fV/o0y7576eTGk2nyCscVlMw88XQmjE723ncvUlac7+zKxg7/duHjlizLIKQAHHzrp2DTFK3kp5E
08jC51LfMoiwnFFox4FwAlFiotjsO8JB9CrAQOkUr7wUqxczBBjcJ2d8FUR9vrk6JoPF2Bk108cy
Se1FFTyKpcJmzVcNccbNaRBxjEHRtEw4aNaaKtI4QqXDfAwGv6O81mrQv9gpdzD31/cwKXfN7jZF
Np2PWwsjkTnOBjEtPy7EUnuZuTTx8OxNw8R9TCmfARYVIbcorGffkLLiFbcT4bhyAwA8RX6K5N6u
TjoXYTYwNhtjb/8VyKXPQXrIXkdZ6eCrx/GTQK+TToF18dwpzXW+Vyn3Fd3sXL0Gju4KQ+w6e/pF
zYRvmlDKYqsdmpEPVfsG2h7nHMWq+OWYu87WbrUhw5AVpQ9BAGCVuBPRopmSksaK6ZQgRnHku71H
JsgrQ6c+KvKCD0bBHLGC5eOqBdOl236eyU+xB4xRz4gaKEhXHJLuwc9sHqBGJuVGPRdLvZea3oJ9
yoIhTaJpmMzLUnIFmmQS3JFuUTYa06suXo6n47lsa4hiDRmzzpx6lHkYFiceeCH1FQ5Dc+7yG+7e
CCaJOXkvm7MoNlewuTHXiVrrRoS0ToZ5UD4nExXgNkOf1wL9E+6T6NOzXoTLtPta12LA6c4f/5Y9
AsJhSVJtOe/l14JVBIFUevrg0EhZscYm0dr6d3xh+we31W+9OHZKi76Jx/cQTMykEmw5WLsGtNBU
5zIFHbpM88s6BOrYWZHwn3ILqEsWn0sQXMAUBu9d3BxVyEOZjfJ3JKdd5Rn3IENVEMyjocVRX17u
E35WBFLS/WnMyK5gXUHKs53Il1RngXF5gkOpuqrgqZ/yiVbCKnSeyI/PYrxxjlkDJ8tmidjmuHcl
y2Jwi29O9C0MvY8zOH8p/MW8L5+tY87Nh2M5eUVUYy3xps7KoWXjwo/6aCaY5FRUZCSnmyk9sOus
CCH/+J8xPPX9dAUmWc0pyptcZB4wY+UieBFwvlC4wI1yloCa54LNGgtF13te+4N609QF0RlOn9Sr
i6vmZ2b0SKCy4JcqzO4CjVWnXUItZR4oOItpIfoRHcqTPssUhUNf5ks6ObaiLE/0E5VXhNv664/+
UFdVA0ZJyAcedqYlmull3Ldf7yESWOsrqdj+ZEUzkYCJ7rHsdoJ3Ge3XgdQH0gpiJ51DTYphD1lz
aSrlepq0K8jMSnH5ju7H9Ls4WRCChx8pxhQB5HysJ1ZHNR3ablVMlzH4bT8HmGVSwNQrBX8E00LG
DSF3p5flekJTY9keYOtY6AhdU9PVW70M1UXEDc4EzghKkalavMRN0uKUhmJxSmL6Tf3aH8r5KlYx
eiZinaiBCmzuhbi3u1EZHLaRBnGyh1AIk3+S28f58Ro1DzKj39fUiqRM5c2scRYsSWeoQK7/3cIT
4xXc7w2yqZWtZ8mpXLDrwzAGVYhXq2koyzsmgJMhoDps1x4Hc6hXRvOqLtdlFShjawTstj2qYXHJ
TcjOHJicgr4YnEyCv7H1GTk92criZo3dPbxmVwTl1kelER1BdXIpznqC6ypAkG6lS+SsOaSxGN5X
pPvbtGlmBT2lPMymqU1zHYikqq0dKfW9R/YZA7kyNBiw4gp0bTxOnRnDTdAqi5/BbwMAzDOvCXgQ
eBox/JsrhkOTGQTXfSGVDww2d8bvViGmuATbgsQtbiS9Ja0CQZT7/bwqXi8ZNypZeubfRGtnoAzv
lOomTr+yamLMn6VMw8decknzwfTz493IHPoia4pHjh294U7rC6X/SBKZdMYo7J5v4g+SMRbMUu7c
KyE5o2nacPvsvp1uddEneg/VXheZYBVO/f0+EwzJrED4n4zaQzv++drKdre6yeNzP/KSy2InIr+W
njkcFdkRNs0kVlhYwBI1WkLK20YcWZDvARYsGg1yME6i8KXMdy3Kn2vlb8QhNS8FUx2Oz7CdQm9T
vOvIKu3zVl0IpZXhdaKS0XLu5a+9HRulCjkyjWqqLi6eHMGhRUV5XwwD0XXRbKCLo/ShjByuWNzK
ErWqHScX9Y1wmDgqGKaTRqFco4VuHlg+EexfNhrzPJRbp57V+rwpR2btFTeDdnSe3v1J04Yd4EZJ
aj3rWhj9lYP6YYjXjFB4xmQmAz8QGT7gWmZVzkpfkvGliUyJr+NpxjakYXipmwNsyUtgLq3dHX8C
guDW3cvD7lb7AYouUiieFYcqxJZ61PbI+93T1Gy1xhvkMZ900Cz/Y+gKuBLPiSbCX0nxDEbDMh1Y
1zfDbN9kCMCoL66gqu9ZOGQsfr25H0C0nSCfRUGetx9S0aWJNgDt+ULqr3m00/WcmWf72eEwwxkf
8DY+czJ0dNm8dByvrqz0ehG1Hj3HQz06iZM79o87qhH4u/nwUxmKOAbDHDGeVsRrM/Jt19dRN+31
pvkU9uMkposUSqJqvL2Jl4EXCgXckKjb1awgrIXy0lz9Jh8nHNET0VdISTsuQuKSubDGOfbVwB3g
6bOMf+2ICMwuTfVVNtO8N9aA3qGQY3h9e68JAz0IO6ltMgJbYBGcFH/GkSW39B6YPefc3DCTOzFz
8w0MGo9WYpI+oi1aA5QRs1Xwsrq8NNoQQMQb2Wf2MwqpqN7dJjdnTiJ7gLCTPwEHjnXdVac21Xhv
KMk9lDOoBAzWuOejaeJ2T/nhAMzPYRtfVAknpE04Qx0z8056oG0AnzzPSiT22kutRuQ+gJ69KJb3
dcA6IiB2lzSw4BcLBzKrctTKOkeyHK5Q6KLnSpvtXWy4txN6M4O/V511KLNGuwhK+p2slKfC9LfP
0EnvS9Todw8IkfV8sV3ty4xxo5nKMpihknosNZfqN+Ct4LNM2G+Whzlqobr9vS/CT23S306kNwyv
IcxbIUZK0EEBW2AJY40bPKZQIOtqgB3o/2zs3IDEAzVk9P/1E4vu3c4utoqS8x/6GbGXvaN+S4Du
0ZOXwr6IJ//IVUlEHvV5jfcuv+HjHkYYe+lijv0qnL+H4KtGWO9jcasfNpDwaJrC3bCif1hurBul
9+XvFLdzbPhrR0uORwjchGMJXdOMma1/hiXvnjqrRvNSYggf6d7cL4X9tiV5C+YCE0/Sz59yUAMy
cBmhG99+vSliN5xibdWjKa3RBLSmFP8KyRtkzf8j0KzlnhLuFiToDGmTqRU0hxM/o06sNoSLvKYQ
xyRONybbhgFFtqTty6XcDvfqeSS7IdtbSxL+qXvy0iT/V9TqWuTkxKO1zpvpIYZTklvqemk4HoSP
iiEpsyjh6z5jJZjIDBMXgU+XcklztnNUmyB9/+k2AdH3VaUM3akvY/dWhV8rUa2sQPegbVCgViLe
VEuh7HB5X56elhsiAsinO4zh0uXmrvdH8kc2WhiDNXGsw8+qj6+tV8UWMsZSOqlmUTKtLPNwdie2
uuV/SxU92VGvraoBzKGsngQrkwIhdOs9bU0SzmFg9X6O1WK9rQims0zCAxCMQlVLOkf8+1VePNEt
XN3JOGADxpKpYw7hlJAg6J97KnUMy/t6+WKh0o45/2ld9kpfiRQ1aNXSD+WugYrFgDIKoVJemGcA
1m2iw+tysQbMMKNKqRJLhTwAFCUWnjwA4KMAGEYUKNdUZmZ7BVsUWOZkPgpwDrYODO1HzAh03ZXX
46fFSrfgfnRmic+ZxKDDmzyyq/j8bJZiIs4OSbzeFD2pyO38sYywb9/VPgf4J7ldidKx8Y8PJ7eF
CbLoFy+UVU/YLgnj1WL5fJalm2PMbFmXEElKuIiYwBzNpyRmRwj5RzuFNFPZpKjNJ4P4NM5q97sm
wHHQndtinF2dSuIiqPBByMVSU8fjhluISE5vwN6/PybSrp+7txP5TJk8CNDzIhM63twq93GFzW7y
JCzNOBxVlzlaUnnQz4OEFwuUAp8EYcj/0HXLjegPALvWHtJXC36ceX16f39zSsiDDV1V2DbTBrfw
aypbhXHURuIXV6tC89gDL+bA/0NE4YIQti9an+6TGDlsWi0bQr3C0lRQmutsXFSBfKXwRoYxkX1g
l0L2YNOuVdRLSjdDPLJ7vDP5d0to8YGdsNltI6jzkwxIwWgi6XC3PfJmjvwj54YFH1ug/YOKd7q0
T+RaSCPpnSApsy0T2D0uyWtgar3RKF/52Hl1DZC+BBj3KDX9XvhPl+XXpFy1WJzmmN1I2Z7idVdx
88yYwJU7j5C5tSrJxLwIJcG4H3b35OFwfqHWG5WZMHBzDHeaPU2sM7YpKOi2y4jNOcal1S1JXF0S
mUXD7ayqp/tBqE0LmcFqaiTdkVfS4SHe2HSbfsQ9Gr9ifkU0Q9k8VBLJg+3rh5/xtlho4LKNkOSY
BjlsJU3h4FEIz8zqAlwSppzvUG0gDqRpthpvGkKGBUQDJ9yhjdWJGnolN27mNejkCx0optSBORH5
FqmXNDYC6u+BqYEe3IfHoeGzOzMRT9jbyy2q6uxlJp/WuSK2QyOzY2hkrK52FwugJluqYFeH0Ue2
o7RClngCYyxWVWCrOuzPL8zfS22FwbWJt3fHWRURYTxLDxAmDknvQoq73E6z3AZtbmN5PyHyhi78
PoLobT39cG9E54O1dMRtr3/87xyaomGAKOnXR8hEwEq3JxPezVCtj0fWaTGvkCYNwKFKEBXgbc7E
IYq6Oce9hsIn/vysSJDxiga/VlrzSDdn9hDa8qChCPc838zuN3vIRfvVKj3JwkbMYcQWdZXFNVWA
lZu5w2cP46M31yDLGLFJFkpewrW7+wjBvUn0mQl07eC5rgB80avWdr8PqlTZg4wW8oejVWCpI9CE
j+E9VV05liZzgTJtmADU8h4+tCNQtmKMSRPhxIOwCy3uPDmnOth0OSMIuF54w1gOSsk71GXGzX58
+pgqyrhbXk1o/AK7OwndPT4IKoHPxlspQJfv79YOLE8l14O1w+tKiULxOmQwzVapdkKEYN1WkVWq
ytFASVIY1ctaxPDPSmUThYMZDHOB7nnOqzl+TJ70Y+HOxEPPEyuOSoFM9IvPscq7Xn/fIu2fjsW9
tZqmDakeeLz9xnMTfdGJMfTj0Jx1GAHL5wXB75OEyO9kZIiWGnxSF95vX8pGEMvrHPEZJZ5SEEsn
JKwqKEfPUQhU4GyyES7W6UUqkfvKlCojukQPe/KwQe8x6sqxanOq3VPJNIPqdXXuNVd7VmJJznPW
K7EKkmYF7gYcvnEUi2rJ+GYbhxkF8kILl28NN0LZfugt618usHrwelaJ2Uu6NNePS9MIwmtUxSXk
g6uUhjSSgd44TMsp6UWezBpt6rjey8Mb3o3f97qprxHHxl3yPCvA83ubTJwPfHCGU4M0boTl05lh
t5evqD7gV0E3YEF8F5f8VXnU702kATXjaDnF1KzviF8NFnmrbofJUsglvdtVLhgxLNx0/1cFjYY0
7ykMCvhcZG0FroaMXPvvpW+ck9UAd9s+m5LIVZY+OB2mBjrm0S0Ld4sQQ1W0CCoRqubNBihOex3Z
heSWWdlDPPh1Bpo+fT7iT01+A+r9Ngnp+Qs5CtqJaGp0on7d1+m6ibC9Qk1NNwa20EVtJk+oSZFU
pMmcaFYV2yYf6jpTwbL3MWw5Sc5yhT2aeSLxQtj/XMXg7h66PYJHy+noM/pQHi8QT4q9DhINQNMI
3Vd0P+m8flVzqKrHUOSKu6qIcgK0+iCQPrQykwYHtEoy9fTVxqlVgdtf14UovUgDxvPm6GH6BDik
iKnOKww1EQUtZ6a1lBFvNgc0gCllapfKSMBKs4cB1yQnwx5GhJ/4nh6rSQBGofl7KjW6r9/oWDon
8ZLS5IW77ozMvHer5d8nJ6gvA1Wj3bfVRu3FiD3aFuqNw5E5f3KcsOe8SUGfjMqdJMfaSanUFole
AEkof54jeXxVu4saPPsV0BCbHNoNOCmlUBFuyQ21f5Kzf4lyFvldNackvoMyFvnXV6IIl/vZaP8y
hHXO4o40MRu+Jhp53DxYe9kqpy1Ks2qulOMRzeokSaNbKzy+ro0n7XgkeYBk7iyreVmkqgxnoZaK
150KlBTtEB8p/0n72OsLAhH83hEze9c6/XH0mdlOc7BNYPSC2Hkaq9VIQSoSxUZskRZQvsQN3zNM
RU3Kwh2fNWFL85ex3uVhpzRrcAqoCU7qqbeKt1E9eqlCDCEc1qrj7R/qM0kot1Cvns9Kzxam0T85
JTpECBQAjbGUwnJO4pHm+hCdXwGZlo4qpyWOnMd4PEygEpF9Mq8RACVSup5IyL1zNWkhzx/LZ4lm
ruOV/zVec6qUAZHH6o7jtDTulz8+t5zpFj9jFwIAtBHSca29oolf/khrNuhaQuKXAvUPysE6/5/T
IRNllMQVeaOSR9ItPscud5Y74Kj8ZHEP+fz/wfrtinnkUo+SsIUlBPnCvycGC39NRMOFENJL5Pxh
LUGFLSmVettUDgDUXjYyWfd3sKH3/iMq5dgzprT7q4f9zQipKT1yxwDtLRKCPGs/d5GNDjyHjGCb
Ic1vHT7cz21SceO1ioaeTbBhiqVaI+XUyQc30EeSFzim3HRGisX4jlCYRXNZo0fEarewYhm9jNYQ
tqcf10M5y9t540LI3yHdWcsw793QdqXOlVUKAI76ppEoZi14qeMxa7/pQiWfn2wFEM2di3qm0rJq
u4IUc68SSBNEZTIH+rij4BoLb2dhJjQReuYQVyml+bzMv8OJNyGHKRtD5uIZauxyGcUhZBCC5g1J
SvT0iYhHL0hd8sdWlkp9YznKIGUE6X8uouE4VxObDnwpGbr2Fkg+H0y4IMI02Jj380vQMxYIPI2x
dpqp1RE6+z+086yO4bJWmW/uHdWAJUWmn5ZbnBi9p13hrlT1w8mxYcfcuvwHqiwGRnVUWUw40g1z
/lTJsoYkBE6VyAW57lAtyAtiyWZ7qfef37A2aG7+6v3FiuhS4eYAMOEqj4JUUyAWfaJhvV4NsLog
UrTpJB/EnR3MdwkL2tWQqHsTuuKjKyJgrdHtyW/ZAbakub0ab/EQ4fqWLJKUrLxSBEmeB+wF9eNC
Tx4GpQQOZZ/BsYvBhfhJZJQKXG1E7cMvEQLrYdW9ZJ9caZWnHVu4aainvAIHt2wNT6+r0TNXQuTg
rCmls3MKF98dYXzqu8uGZ1dyWe8xHWC6t0DYnhWu7JBE7q7+5bbKdg/pLE5ciYQhyc35QwhfmO0A
okbjknOm8bXzaX79QUhxJaHWu1d+Rs+E+I2/JjulT6XJcDJFmhYuVwNyf8031vm+dOisI4WN8jrj
cKBmm6bjK2dOBnvF0onr8FU+lQIcDeT9yGgjRWOl6iXkMGmXm52E3X1qZztrvAm4bRViFHz1HDqN
giqdSzIoQfFwViJRtM+bNThovDH7d0adSAcnNRASabFgM6Fe4rUFKorNBewNZUT/UjM4/toNqDQB
gBBWRdUHGMcvHSuxdSm447rxC0kr0N894pwaV66P6CJlzz9fzmK/R39hL42iPvE75MswtD/+sJEL
3M0vEW6jMhAEOdX4Sfz6RszJjWoZJh6JUqCzl2Jxu6iMS7UD8TH9c4VzZZHdN8s91qL6FpQ96xEs
gAKky1jw7dU7KyUk6uetxaxe4JeCcpTWgwyfMwyjT5jKzNSF7SuxcCaDH04xkBL+5ePQ1PIrwGQ7
BaPgA8vovDHnaTC2UiiIQySmEA7tjx0Z+ExQwCzlst2ulShX4L6/x+2JQaqmE7VwcKNqqwjRwkdy
Z1ewvD7XFrAd61WeiQZn/Iz9Z9RfwxqyNHP5DZzPuih8O/HNTwOhnkYRVtTDLz84ovUBTxezn/h9
A35U9SulVnICIPrfwaylfSa2yhpITeSQadRaYy4DwtZif9pLtEws8YEUac54o8RFGl+ql3qmp0UM
HKC/oR7uf4weN7Q874Nn0dClfyl4AsjeNRPhOrLTWrXQeOu7Z4IeKAmfOVL+tTNkCWno1hYacPot
JhTCimNjIjmVhybYstnDUrdfD1L+mXBKacndRPm8ZeUHF4RA8qyi86zks5F6GBVudce3o6qqiS9K
lSPSdtqGGkWwZBrfG+9PFuJg8k5cpwrhsBaOT2NcNgaWjlFPbOWpI3RS6Sgf6QmU1cXL+aYNSllv
5ewH0q7nJtMKm9Me1HzjCxyu8zJVNGF4j260+wo1Xm3T/1RLdW5zdBwphkudbTvFC1iCXeOtogJl
9yxriMli+PphijfIS+5kCcYSSZ96LjYOWKO3wfBxg7xcxblKLNsXMdBBs5XlT2e/T8BNOdlsFePz
IqE2+R14/Z/uqug+9hG4TXpPe/a9qIFK9QfN/scnt5BIawH6Su4qe20PR5CCFuaAmD8J6FgpxpSP
59C5X6IH2PiAnHGyFoaugoh1G53Bi2j0J8Ow+fGbDKv2WFu+C8DZnPHu+GZKS9rB401fszYdO33s
12VMq2R5S9vDtJJtRGLHKr9WjQNkWvqOYlka5PdW7LNvqJPza6T+g7J2Pt6iuirTawK5adJHsZyE
hjf3TOdPNjshHzYHHAOdoj3gV0mOEPxys+3tAwjf73qg5EVELgRBJ8aOK0BUWfqA247mUZ6Aa2Em
oZpdQ/GxXK6U4y8Q3rFvxRsRBJH42EGMJdA48nW0xEm8gaIIJkTUEnaEV4sy/C2VpFQorPApfZWS
qmaEd1O/wKZ8HN2hUKSYuY9FcruTpsU/SYIbO/kmhYxs1etqAQagTCSWvlrIz7xS9/ikbIDIgd/r
Mo0HWZw91X6YX2FQ8w3GXewR+4UgxT2KPKbeOCFYXl2A4kKHmRpFhSNWFdBDMbAp4+h6SQxxI1XX
li6WNHJsgFZJy35/UlDUq0GZOYYZdCEUalwIrEX6B/O73Wr9S2g1fcLTmlxwkCREisMEcKO73w1f
5xIAirt9xMWX4k14wEEUMwcEUcvIIAxXlcoaeCm1eKhxgvPeiLEZzjV3s3Ht8puzxmzY+Xpq3apq
/xbrvFb92dCQF2WysvgyH97Pq0rTejpgXmwP3VAcf3YOlSp+i/88EHPalNojHppZLIBUVlW8gLU/
CYOKVu/kIW8tg5T86t3NmYeqec6UstpEApSn2FPztJMg6XSrXxHNEsi3jDCLZXVjDYX/55OeMXVK
yiqJ41J9MB1/DnfCjrWxg3G37/AwSmD9OQQrtpFHvHsFiaI+UNbavzscV9Jzm7zamDY0JlTfS/Ja
DxWo3MTcMEzFap0vf8zyYpIb5xC/NTtp4NJ7XOgGwrsFq+U+n2Gpa58CkSQGl6/VdF5eJaGRyGs8
xHigy3WR1tI8Go7ofukjXzw5MmgkpmI5ShimwSqwgcWopcLVTov8e/9NYrjL1Ye5LwYL6twaeKNx
Cq0WLTh09w11FyN8KPnNSkr6sJPkzVWYnQYlqe5rSsSHa1cMHABuQo6GI3xx3u3u7Ga3+chdeZa5
SY6rpnnrW5YnQ2MFi+DEI2xvJS67LDO12D25lNNoC28z+XE6BEmAWOcFsezAb+fovfW0Dg6pOr4W
4jjJ4AdeB25r5wdM0dQnIK/zlkybA4qSazjMGCSHXKGla+Z3OHDjtYZ/2LuVByL1kUdoP7EmbcF9
Cya058u+lCn3iGwLlsI/fiAOb1wLj3WWlJM0YR0OuZwDqTgTvVlfzjpnkjlDzICcLv9LTt9WnNNI
kSCzXgNc2TKqT0fwXGBal3kTsmnGSC2msgGmTSu9QAC3Q2+owdzdQxTMBxXNoz651Y5pWAfE0zL1
ijVlVxVsKxl1f1h8toy4LDW6VTdElg/kcO5Ye3pwiP8WOCfXyVlPUzLDKKUMJk7hP814DThl6Qh+
37+58DKFxN1I2Dkfxqqeulb2njQ4plb4WgkC3w3T1lcS3pidBq8KgN++53MoglYOuHfWbFmwBCqO
mUSWeAvm7xID/6m/h6bKHzbcl7LoqkcRIRFOBCfeQTjZ6Jv1eYIJiLynsDZn/sughTIeGixu4h30
BhjymJdbpP1AA0+PRhzkP0qGKk7w+sG4EKFvqXKCDju15Xh3DC5FvkGqwhG4f6VpjEs0KSKjR+Rf
BOIGo8QKJjmonOLl3TeOy3vYVOh2juEocP2RQyBq8H9hlGy2JnQD8aDOLEXMlg1xhWQVMVmXYbsY
OxOEoCxgyuERmzQzaT8DrRGU44QvcbluurlATtsoUqFifMn1vO9OBx7tnPwxI+UIlPoos+BN4YCv
0+fs8IPcXMOmWDrZILBAbErXP+p40QrPDd9RM/8bAEzwx2k5XvJlMcZJsXBrBdA+GQcjDcTjivTb
Cd6ggfcHCWuWlapSKGis3NagNCgJtm9cRO6GqXnjM4/WFUx/9QDuc67t6oi7N7pB5+/oqbRHwLoy
RjJUbcT0OB5Wvh2lWINlvF20RW21xYQ3gPW5V0/OZEu0xWqaa6+5Ou8lvUG+YSsqWhv1fqi2xxeB
wukke7NQqPjnS9kXD4zXqj5kSlaWM3kM3a1jrlpKv5/MSX4RCI0sUk3N5XQ9Eh6pkvJEpVTFYY2I
ohmo3Zzl0/qp4Xw0Lq6KNMcV3uKuhfFkLQu+fE3G4nMSSGlDBzQwpOhbhIt3lBImdlVWtR/NMRJA
20MEFKYjc+bO12Reipz1TnVfi5qHH0qtESiSGBYrvEV5+TT1OThHE0yWXxBx5JwFn/6UCk1VobEg
Z6mnNkH6GzsdH1T0D5PNtyPntHOuaUEooDavk3eVedpPogu7+GWp8b869gEP0kwk5KL6ykI/5Z+w
iuR+qfEwt4k17CGumdE8AkHLq33B3jz01w/Fn8nl6dePyUQ1wOgi67i6DbRzmdyCMFr9rHYeud1e
633N9oVamUB6ZkFlIW+GLfF2RCa2J1DrGHsM5mHKFbY7mzl9JxRuz0DOkva+0J0nh0/GDoA3Gej8
CLEZcOSeTEounUw42qkkeSdQwGf8OS3NgRjQhl1UcnE/dxjKwt+uECgqjhLtWlX7bgpkcbNyZ1uL
WcFjM7iCFuwxcz1vlT2NOUUASIpoxRj4hb9FTbr17Ogwz5gR627WtWDbuDp5V2GiL9fLTVcNoLUY
KFWzaAwkSNh0sU16JhNWiiAeZnyC0cjJldowL+LQ9co2qJci+w/E2AGYbF6TWWjT1dhM9NY1LWDR
cEZRDkPOl0+5/XLuruwBjRiMuU6FBYs4eVc1YKCwiN79N/ZnFkJURsrN0Of1AE7SSG2iuLsffXTI
o00xxfmYbmaudCFgFfON5wrBdiNbhsdXITxgnS0MCkFxwMr4bU1fsRwJ/nGtbqR+v0te7PzwZy3E
BP15R/kNTdPAoGVEGJunH9JeSdRg1hWXdsfhBhCN6UBHjPxiiih+/KkdGvI8uddzun+THjXOSm6F
mkd8f6u/aW5TRuoFEVLVZjYznuUpBoYWbcXulqStvnXssXd3OGJ3L3wKFUJHLQMOdC6Wo9oU5Uwi
IEbXE0WMKkeHlF9n9UkWS4tPv0aLpB9VO/ZMsxZJN47iIy5cU8zzfmkEUNA0i305uKzmhoTEn1Uq
emU2ooPOGma/vTv2Ex6w4a1idhoTMU25uwmxyG3oPuG9NkmltIjTQZPpgmly/1Vt7epPYlxccEe7
WQsANDh/kgVrUMdtn3jkMABMtvETxLJzBGVtg7/z8k08ZQs4vF9tWojRkB9N7sOaNWl266SKcE7m
fkKJZ1eNT1+9Ebv4i8z6Vpp6Jk1zqx1HBoSp4wtVt6pMX+omKhCbjTrHxQqInOjhsMHrTcETxfxe
cWc1jNHTnsRUMyruSkpOxuRgri7cqE6E+u3LOuZQltPOtks7dc+pwsMX5kwLkCYGQhLMXAKFLJvT
IhBnJhYyISBGwciNHLrWBa+f7hWYIZpD78qOCp3LS4/ybUNt5mJl+UEsPbsEQK9ceMbFEkX+6zyY
/MLvRPohsE7wLsmVHhevMN3xrAfWgHQW+MXnXD+Sy55bQD3H7tgD/yvHauMmYeDB1g+3RX5Q4Y8+
3wTrtwcpm5qUjGVZDpgyqeEOZs31UZw0wEqSfxQwQibGpcPDUJ6AWTk3/BM1G+5z/o7AIUGfhl91
yV7/7bDKdQn9AFc1VqG5UOqvGFDHYKrFZSUsv3848kuT6qEfk+tHeqZBXIC06hL1AK7gGlmk61VV
TaIbZSOm4bxlEUAAWW+iHB3YyS5/BpOsqXKglfhdmS7MnyRU3Ize3L6ZKrQnEevIb9vTJcknKDVI
i0kRT9xuUrkxR9YgypfR7DRa41hWwC2X1Ahz2IIVmp5OEzmoQrNbVizehxk8k0VzwxtI8L8TOoe0
4qrUIzxwyeH0ZSce7WA/U5xDnmiwmCrIFAV3LmRhuP0BMndBpVTbAP51DVg6V39DTaO4px6uZSHW
odSjhlEePZ7Q1coBZghBJOIwlE/x+26dIEFrIAb80D0pZD2aiNYGcgMXp5alHbNsLqFpWwuI56gm
ONaVOuvbpz47UG2hG8uVHyEqQDjXrm3vSHVGo3UHYbFWjOFqoeodEJc/X1Gjr9iQRvGxnzLrFLzF
DEjUGY10d8Rq060zPORuLlBOebmEfmudsPa10RZGEtIMtTUCoy0J7dUsBXJZvbUaYBRLTRfs604j
P0Vr4dZzruGhilL17K80m9Cx62yOmG6gIE2/DNoKjYUr5Uzv4gXw2H+lOb0jjRTUOZVjwkOVX20m
aB68IDReCRs30US8JO1U1lWq8BUCJQTJijWzrAQ8CwLYZwFiBVFErcdHM7lcLOLAe4wkTGImPEn+
PtypEBX4kTOwd3gqMUendSIbpHec5rRertKcgIR67QrLYO8R5+zXKTh3+ql85eJX2/zKB33QFbEs
6bRQ3hthrXa+BWSoqunu8tB4+FBJS/El71fUxvAUTSjv1i5YNJShVkPXeucSVqKM+0r0fy/hjuUM
tdNIdUUgIuCC/LFvZAZ8+kx0fEQfUDYoNAC6gCKVbN0hbFjKQcLteoIXCb7eT5tJvC5MlwQQ+bBb
WJoVwEWcmkkWz6lb27HN3Z/JfK+gM8cDfGfGQFbb7q80E3pEydNMS6W5Gr9XM3P+GAgBCCuHCRGh
xXErkoPXGyEjpxLx8d1P7l82jlTIVGYJl+BTjo32Ob5aEc9qKrYr9H4Jnc8slOAZnL5rbm0kY657
bv5Y9nDu0upCl/hMWlbk/w+SMxFP6lZniQKnFO+nFy3H57rhKOZLlmexhz+/Rt4DifY9FUk3xXVs
uwd95JivrLq555czuEvWJUxuCKEypXDIPstOEX4sPRZ2P2B1HYwP0N0n9vvcVub/1klsKgaRDtnH
mm9zZ5kkFK8ypUZ5PMGWKpEpgZaHLhMLyrAhRRJKFmNGd07IQrdnDI+xvSYcyIbLiKH2XZkhkNuD
AnPlGWGZMV+VAscWfO8h/6zCTDz/61ndjEhSJvhRCsNSSJi73Jwyh27H6stGQkajG1jhmQPqF+dO
3MpIu9rpF5+Tz7ngHoWU00rdgyso8nRgCKfZINBx88PPeUBvXGpnG+1yDIOM/HeLpNX6N1eUyXaj
rtaO+5pFYz+glF3GJCj9USmI7i4lsoz/v/DOtbEVi0x0HKw2ajOKWxzyGgtA98j8zh9kfvPlbi1z
qx1mdA6uxu7x5RwEz/VC9P4jac1AwrfvKBSrmgijhjs2/6Xy6NMgY7JeNHXsfbIo5Hczk/ntEaWK
ONoSEf4nOhlZk3z6/qYiBUSFp7hS4W/J4JCmZ5WthuVIpLTC2uwN8tiN+rv86CnF6E3ErEo7Aa76
pBCO84nBEs2XRmZc284diCSPqQVA/DOnc2sOAGlW3h3juzsuykD2YdGC9CLQi0d8rX0C98cd3Ny7
iQ/qnVhA0ioLlksQxuN4fPvpp0qUzREJfFQDmYlenKaaC+pWw8fhBrKKlgc5F1mcbROVqg2lhrC7
qnvIMI5uiRcWV/rlalAECgVhzgF92We4QjG3QJU+hRXCN6J1M6J+GbOYn2/j6u0MWn4NY8oqvxtq
PjNZ8zjRtpGJ0NRGGVIJCvMN6dZ503mtenD/YPtPZ3FVyTv1BnfEpACanDyunUQEM/zbeBQeV/7K
AonzMwSDDhAijewcZDfWeIwvKHeGygQehge+GUcYM7CjT9wWZ3Jh7jbuvw9Bxzb1XPDZo6SOWtqb
0VdLXpv1CTS0BJ2WqHnJ7bV51UYV3aGkOG39tEVQgpZBo7npprhTSBFX3L7xuSwQVJdgfzhEp7WE
dO6f74nNfEvxT/+Q1BEprWJhg4SY+QmEHRi6fQprIgudslF6EHPA2f9bCWaSDTNWa0Wkk+R/M7zI
TZcs76QZpgiN4bGGDuniPuFnuw+UKbMIv8RtG0TMYKJ4c0lxFJVpL/obAttZxKu+TX0FoWPKs9Hk
UuFBjVJTmzStvzNlz2RWlfqtsQX+bsBSvpJAbEAtgDD0p4izMeTULe9fgCgX+hTqYWcpFVPe6GPY
QcOYh/+NncgW1nFEcsC6RG57m6D7VcAnoxK/EpsbRy0DCkSPmC+VuHmpH6C37JSAVqYKn0ImyLar
q8p49o5IjHHN0LzhmOwJSUHmJNnNHn1XLrTbCtObfmaTpV2EK5wOkuagEINNpfs/lVZRNAU1puGA
DONnljSA4tU/cXcfk89yJHlaLI2DWd1zUtFcSg3me07P6SkNZFlUaWzTPJj66LsslKhhfLyUKTL+
TxyrOgqZBX78+PhfsHuxddGsR1PvxSBgCoCXMeW0Kk/vC+sgtkfWdSg0oDXBQ/s6yv61vCG58xm9
uv3n/sOGJw1Zx0wv3JSr1ZI6XKWJj81gdtHEZfKexNT+LNkZT4ax30Wb32so/7+p35Y7V0XM2id7
Qxe9G8WoEJos0JwM6wrz4bxBQx/V3W6IX56g0SJcqBJIE/BCoqCkzz6/3Wefp0a/64LXA7vJBmcp
LObvrV6KG8KDv9h5BoDjWP6HnY42DpDGHB/JzrS0F5gWpfofrPF2p8mAO6Ge4dn3YvpTdhEP8Ikn
5qzWORV2wlYGrjp+GH5lV77kbJOBh75s5otj0p8hgwEL+Kkf1ODaeGA1Meq9CsChHaTr75hVO4nh
tW+nefotrMBhHi4b0DgSuFggzeb6UtT8hQyA71QTsW6rp1bKoTgsE1YhK6VvWWlX4vaCcjCoOO8R
87EB6sjJRpgS2bj6xqxvHzLtg/+IyhAYtbGdhkxe+7MBws3gwnRAnFco4X1hvqA6lZQGEOJJc3Ux
ns7P1pDvWBYBLw2rxn14M2ob0Alrt9HpxC2e4d3O8d2XczUaUF08LQKgIlXgQOwHHeABT5+bWZVR
Hu0xznntL0GhLyFP1NDljrL8PVzh+L5bc2cJKnTpgnXSGK5vRHruCRd9DtZviNFow7VA/l5ukkxS
ZFBxnBc4miRwaxmO0DEf3phqTjNJbkI5Zvtm85rWYbi/P4lUfQpNr9+6yVyBPvIxrA6IgauQMvzt
aRAd3O1vp2smsI5leZNLe6KD2Qn101I5EiDU+uV3bmOYUb+VVK0sz/sERHxuHoME4YHfyJBOqCE4
U9NGSG7HdiMyPvPuotRbHtzhy2T3X6XJcdwRgKt7X1YeOR26GMPGZyKkM0ScrYMpCbeTStBq5pYb
nVulCxdtN2UXiqqeszfvPJh91dZ8TSvRirEM2wkLjHexNNsn7I3X6nH40aeb7vcIsAgWpZKhqsdq
zQro2deEunMxzDTnb4r+EDRhi/TBvFsP9C+868kPUGrjdA6QGlYintfUh/h9iHS4UssVVX0VA66j
05/oDSuQVGNbB9MzW/pyLBW+blHdAaw5or6Jldyq3bKUlT7qZFaKZx9N/sXEtvXiaWJaUByn6LhB
kUB4syRUURafNV33E+Yk8ChdqFOEmEZGMlcXWp1izg0JhLaqwKeSDedhNs+d1v6CkjuEtzmWIk8f
zaXS1S/mblDUdmv0iWjjoMdgNzZvp6uCnsTBj40X94Nahsto/8Qlw8p44uZxQvha0LtLmQCYpqEG
8mj9oMjDZ+uTwU5HojIayzezTX5+5fAohGOZb1f4J3AEZaIAApqvY/QP9OT3hn/7mytlvF76SMI5
7riKPCZcuoggzt1vtJz2JdNoSuvxawEI2Dl89aHBk94nuO+cKyH2LNE0EkVWjW2i56pP1t5Kzq17
G1WpBA8YplpQyDp6rHCnsYtRPOZVbWort7iHwrRtetbU7RsPch+YwSr3ItbG1LWHaUhTWcBHqz5s
r1yAFnXNRUx/WUIkM0Nd7jl5oM6uanBNPIUVAPN+H8i3GmcGpVVr4KGasVKKiftXG9wXDh3YhAg4
RjZNnchHyUQ2iZ18pgM/vxZJRlta50Npwtu13cSdsZ62l+FupvikYX0UD2Asgp6ZluYQ5maSVJ1N
Fwz2G/y5lxvVLCziR5LsFpqhChSD9hbbmpV7zYYdApPF+LXwq/w6EL4A9boF7XE9il3ViCm5HqIf
M2fOUCDD20s6EX51kJ+GiQv5zpjvXUpC/Oc+QzoiBDlMGsxO/XbXE66K+Khz5xIrL7uubnGyVULM
AcZ92TvgZ49U0b0dh281kAuTMxLIcVYl6vLZ+fLUd5HRWcIjirzroF67vHbt6pLl+XA0DqsEMOBZ
efGj9cJ7KGm2Zw4SnaWBHBCsb7oHO4KcgraWVvsZkBZ2z0ljPcH1vbLIOeLXVNDk5SifNJjk2Ia2
Hc2D4babVdtOmiL8uu4AG7cSxRr0HMTgP2Gal0EN+ZXJxMpVnb2SDQ/xsEC/0ZF4FVd2fKXYIJ8y
gVptOYF26ErNDiB5LfBJTZT/ZDLZM99hlXaOrlEPiWjwmNwPMmJE/wYadu3U1XBFIfjwy012CIpp
ps69RZr214m53yuAVs8Ma8uHYrMDmsme/+vLBW6uacGO8PZt4/tVtZnRFaL49b9BTW8O/p40abjX
aJyvPOSZ/15AAppbjN9fqCPYs2mjDmK0mqGzl83oju7CJq5wlicxKifs+1jH9M/sTu8uu8eBDiMz
lQGQMzXEm085eYxOpDj2kPYtFn3/XVVqznIonwdZXYsC4vgX4GY4lW8yo66o5w6gJz/WeqjscqrF
evgUg9crbqUMcUrwXX+Fvluaci5tnobMVAln5JoIeGbxNKo2O8opXxmuBbo6gS1bqNaVvEwFkw9v
1w4qj4JnOjPQ68nGad/JN3IIPOc4kjSWkeVeCwXS0M0lRjTIRpynDha2cSGEv9mCS6K6WgItJlN2
EzV/7PW4ET2EhZ+AT59S6JkVLxutaWfX2Mywqs/T1KUHLI4d+FGlSfHJ0q8BmMjJA/X+M4Sq+RIb
GZuGJeg3UluAlIQh7KCp6fgJD0uOkTjfRLDxLd0ohp4Oi9OQUZfcnBdnoa1RtwoP8OGJCrRBLeOP
N9PpGXhWGQrBPmrdnGi6RZhu23yt0iNmsp1hf9K9/jXYQ3fNgczi+D6gfIqP4tjcMebDDw0NJo6Y
1LwtCDicz6/pmI+ZaIHjm17ToRZb6pPvgI0IosKH5Mg/cpkSY0oN0TMSmtICAMtMYRToWS89/HPI
6bjSby+EFr2SdMBCHQmUHs8yMY9//u5LaeJ8oBTYTlu4tkQUE+REg4gNd4WxpPY+uCUEbvEoyCTB
uJZaAepaMT/+VDxIkivsZhvs8lxIUuJH38Ba8TTICFhIjpwVltdqZyAJ1CqWKq3YZa4aWqd1u+Go
M95hk79+eJeo0E+6Li2wFM4dmw6FN/0TT7ELILsljASSjyfW8VF22oJLfLntV4p4CMubhfqWJNyX
8zlZnj0vdrh6nqZLgS0IDhxZP2K2lYQ+PUMr3PgJrXyAAE5R/rfXMHbYuN3igvynloEzxJNTAX3j
+diUtyehQVtwKYqPnQj27sk54JvoAaEJqMVLBPN7prFvWdjcYqb4FfKaSTkDAmwpBGW+NIS77OqP
XjYi4TkZQew3SfjB9Lp+8ynkEYj343+8TZ/N1ciwRga26Q9mlnNsF5hc3c0gAhlb0vgjCPCBDmAz
vNbHU+Ita1m73lxJe0G0C2WkD3Lg6J0s9Z8G0KAsy8wKVd0wfzR/myD11tBsZuKN7NuSKrKkxwkB
LHJuGFmVAwUpzGm0eZHb1Y1XQbw/JU3hizhkAHCBN+2coH90yAV6mqvDjZUDTGk27x58yVboU2sN
EGYbm0sSm4sPHDHGW1QfREdAVCrYwL3Awxvw7VpjY1UCmwU698joNA3gUgSQ9AsULVDeYm9JE10o
lsh6Ll/5W4WJGuSLDN044PIOD2rPZsCEmSWkPqtwQsUHWq8zlvOL3sgRQ1GaE+DA3xT0YispLAq4
dGA7wjmq84lq5FxvoJOAnXS8+p35+BE6fKqfWGEWnagnnPUlgfCJiqFCfaL2yHJ2IyC9vym9bIIs
xpQRS/RgxYYTCc4N8foPMHNPgpuLjF7XL5ccN+l4To/7zi3bqsLhVll7REhjfot/fxVTEy8e7/zw
tSVTNn0KP3d+5Bw4s7VApe0LF2hAAC+UykAfMA34t/ean3q3a4F9bX0NdStqEl1h5lWuhdQPxpew
QO764K+GRw59NlsVJcxyMv5lNtNo/EgHHsmH7W5mLIlztaKuLG8VaWQQrQduUcFWI8ekJ6rpw9wu
JlFmE5/Iyb8OAq/N8G1eP03abDfHdVcLAmGeiaoNqcogh0fa+8E7tM88JA49bbkGFJhyEamNKdgg
a5om8I1F6cqQRJdHWKLtm+eaGe4Dac56PU8di8LtIrFrfV4e58J90nA6v0jh8HRcSm3zqZpPD2/P
wULgwEYPX6xZLOyXEISY2maxOwMOo5u6nW+xSrtgzIWEVEdsmVlx1SF8oDraIg0viwbShDhvRmWR
gdlqmnOb6uIIGNUBaH9s/SoRqUq1NsxRpTOhPYnC9UarK+0bxqzpRYrQGyBOYqMH8g4h8g+VGaJd
f3rWFPU/I8qqwP8S2loZ23E9gAkNnKrX5egP6fZB2meLY8UD69Wl4PwcImA5/OvyjEueO0QrnAXQ
dstrwtD1OskJMZLtXo7mfoD5ToKU8r1e6Rb8X3boUUSgbpqMQK64CpaI6dpCjPvNHpBHzq7ah9xc
zTxqToLdSay0KEn0DUu7BSgUon0e/pUI3J+ZQuus89waSFGHzCf4+hUnwRCEbi/uObCJB085idcc
2jLBwGP9qQv2g47uYgZRJIUpjvWb1NPQ+vZjlsWfAqLNpFChPAiake6w5yn+n0GYGn+6y5Ln3sng
pBjREOgtl2xj/ltj1LSZopuIHK8YisgfLJScWsSOE5GzPQ50+JbIgKWskQ4tjWM1Wy/W4mJSWitb
ZwqQUN1/Kol62wf096x1oBzqD+aKAD4ZB0CBw/U4RQf6eNJ65zi5p8qmCqlXBpG6FdmoXJzBwAK/
GOc9DdWB9sce6OGCOotnJrQ1HrFR1OFNUsbmEDKsFsB7oGEJ87Uxex5tf/kKqOxzH9/ZfDmK57UX
5TKmsxoU1VQxPzpcRxtDl5VblcMB8rrw/OuEW4tln/sd/VDdjRc6/qHnG3scIyYBATvSmQZRiCTP
deGkhyId6YJ9CgDPHHPsHcwqfaWy2bOPSJO9da+DKukTzL2P9Rfz9GnNfZvcdoUcg2oh+Ome6ZaC
qusG6h1sTtjdvOFkQE83RQe4AZvSlWXFToRvmZVYD/2G2bin5HNbi8jW04DryVeSPXxt6UCpLdMD
RVanRMys96B5QkUyAshNkL0hNBtqilnwG/08xhI/kEfE7Ja36Xy05SRgb4Ae7ExVKIDAuFIi8vuC
aFFt8lrNaSs7zYuKro10pmsQxr6hen8eWO9/hYEJjlRWCV8PvhvFFxBFN+vbgEP65pdYMQnMXFAi
tRjQRMsFX7flYkCmpiSqeOBxuAkXS8opxUMH/TbK+XhRuJXIW4DTpWBBGkJC6doetxgfG4Lhxyy7
XHas2Y33zCm/1AfNri2gYl5jDRvkvM2NSu9/T8HWaW8nb/6c3SyFaFEFYBrJsV7cH4yXtj49LtNK
UnTo/dBoqY45F7AOiDFs4259g2IkkhOecQpvvS0rEVZ/NIvwHeWCAIY6bYgTLdQdjYnuTWyvvMxR
bOuT3R6msBTD24PAKRB3rI2HnbD/6rBH4MH9cTIU9cWYzDSzlnDkHBWwQVwogDnus6Jy383/kPKF
bDnhSIH4uPuMSCGaSTMO4JKayogxbfJ/xrcr85pRmGjgNuNTGEiE3FVrOy2abztgw6jE1qXp/AlV
DzBrOoRHqGPW9dlxUtXBqOWYXFkVslfDmaKNk6pHXZxnMXtW30oStkrKwGEpWG+OgfbvmGQ91Ouy
gr4/mri6Dk2bczQbL0ohNk3uFqKNZfLmGh0Ude+JbWOX/OamRQpsZvJ/yMvyrHyk4Cvq92+etPf/
H37O+M0oSwUhTpNYMbG4DQBPNuKTQYjpBvfhsAn0aa1VbqGMNNWDLrtXauGEJpynzgngks/rOQAB
AqAegR9z6urbTv/VB3WV38avu3v+eTTYDVjVJqBEGDnGeHr0Sqi/D57vive1Rzw1DaU2aqyY4YL2
g0d3cbdZI4vdQIXexaEqXYAC2104KQymRUxXwsXSIx6D3yFwaAmNHS2uXkASkboO7P4xqfDoKfKM
hwrwU0LjP/cHxwlGQyEKV/DlMhZqWQI1IPbOvTmdpaPg2FD9fN7eUDGuKx2ELstiRt93M7sLvm7r
qwDoNpZIDQOiERZAiFXSaU0yam8fovwLdf7cXOM6j6LMlVT9Src+PEZ/udkesEJQbEGSnrHDrlVi
lv14j6l3WGtKtseUZLV/1kloi4TJSTftjVU8uBbzc+mYHaHNEsvMiy8j4I2ALhgUqrC9iZ7ojWdL
69x0HCQGrjqgEJwf39FTra2opsUB5NP644VImONaL7JvV80fqTVVgjhQPA51zbjWg1YIQxnAg+Re
Yld//cYeaHgo61pcJrhJ/oxzRVbje5yaj1LhZFZC5LmODE1NmsMT1gDfiIW0zHNG0gLw/m7DKZBS
RYDcv/khTCR9MqUxCwPfW/PEqa/DSMkTkbrxHpLHzT/XSoBIBsle254rC0KNKCLGMbGKQ3LoCoLh
ly1JDj8Y3+W0B9UtB+XeH/QFpeWTdzcvqWC1YzwoLqyyz+7FL+BBvkuS3PVj0Z7768Niosumyt/o
mx96nzwvtF8rPywYU0vHI9c1BpHU3rj/9skz4/f0350D48Wqaei0N9L13moFxtbOs/CgTellty/4
nO9TkpSRXam8pvzfDVkIQNALO/mtzN7w5wr19a9mP6ROTRrw5Wf5thA9Hmher4AG9cqaW3wrHuL+
u46ZcIoKA7ZLxwFcjn42oecH9q/TG+V6gRFuxm9TTVXGI86DwCCJDNUmebaPSArYEwkZKvvWNV5r
sK5LfCXmB0BdQa/Hl1+odilS0ENw2T0EodWshUF+i6Env1kIhXg7Cpc3ORfNqWlF2qmXN1EOZMry
DC3ZuNJEVHxIGz+Ja9D+tvt5PlH6qiIFRHEtL8wP897h5EPFJWP9OWHdMtJadpSP8BL04TGP7fve
VeR4MiuuroHSNhl8dxIfUvtnf6rqnbI4qjy4cXk9nU255YCvEnw3MCukOY8sVPQCS1I2d8mjyTHP
eSbktJBz7xirOT2QPfJksjxr+hJgw4mQdKdf89PCvUMd/3ZSBSrbPYJzXpgrr/I39cAGlZkR/oz6
ZBt/C5+Loe+ikzlE5gPzSV/KOZFPn0koNiPhGoil0zNuBassxlJ/mDRUROHclBHcayqQcBiGry2g
f29II4g6V8/xlX0B4iCFM80WnOF7IJEc9J3QuCO254rKoLptxVb/2uO4v6grt7I1VYgo8LZuc2Li
Dwe4sKPBU+gRAI5sizuPpSqP9IK2Ke50kmegRaNeAZUNlPXi7weORjs59dxyZ+/S7xFjXfE/Yjt1
aBftbvxyGaAuDu+Mn+SrnOQrFqqQhNEr818je+NdpcFQ3wYDvGhbOkssgefEC2OhYIy9Xtc6f54o
eekBbKgvFo5L4miJcdyq3TCy3lBIentztD/okS6369gww9fWm+L1eRwaxaPvlpromUMdAKqdBd2d
7sE02pv+KtkE2fwJXwgyBilqvx6DnNdmrYIn6FkB5EMp9UpQyMFjQu1QL1E1Mj2OaCJEPH0eAX3h
s+bXDBQqroCVVpPb+yCu99J9+79A1+DEoKjt0GPhXHJTZcfHQEX/aZBvmKtrEv/CJq3Pl4mWwnYA
cFxF3f3Em1u/4bkSwNOxRfR3zaeB/6s1+cdNKM4TGpqtYA6v+3yJtRYJ10dVEjASbhXWmXh5BLD1
nV+pVs2n7GwLOtVlKwmhXF9Hkh6kT99LX5ldadkbIgvVCvMJJGMspLElhEBZPCjVZ6nrlHiCqIgi
vqWtzetv/lE4TFiZaf+OAvJmu+0NvqY9eW5NxNTF/jsuzvXqqy46nq+Mq21sUdITq9KyeSAapIkm
ITEJzYcqoHvlLQGVo3HTx/GZ24h0P5QlIr4MFUCpJq+alVht9oJ3UIkP37XMlxPMsv/zQmWF+kBJ
ND+b3I5wdAWlDxJhWsbCmDcUtaqnuzc1r0CABY/Bsa7mQel/66IAIX2dlg9YLw1nYR9/QuvgxapP
ceiy6nZLI5OtdUkHA6CQzN7qfKkG2gz/l2uscvEJeq3d4Boipnt6C/PC5DUC9DlEee1WsrxCQYzF
Z93n5caTX062XCdDdPKppuPY3NZlj7InTWyq7TfG95KqZjo6CeYDm0P3oTmP1rbQphAaDKwlPJeZ
zvdC+eDcwb6YhPF3brjteL+Pq6HUabiSoB04J5MbCnKpnGYKtOP1goTCRCaRjXtTVJ3Hr3qLc1mS
ttUdFNoeMnwKSKNuwu3uQI+/EHisxwq1ZkBvlkw8AVh22tb2lM21APvEHxD1m/5cpzmO62Ly4ad/
G7lq/chLri9If05FUGq8W/7M3PE6Lnfmp0A+dPhCWqlLkQmZr8CcJc7t8eVMBGI25ilLpebATyD1
rR9H2SHCQ3vovVrwmjVwrIwhgRdiU2Ws82cM+ojf+YP8CgKcbBkV8MEVs/hsWg3bNQugMNRgXYNz
rB0PT9vAHIpIp5NAEwCI2gaOuHap78MwOokYI9Tq/a7nJOivoICadSlrk0KMnyn55KJ/0WZJhnNE
ORX/I8W87OYva7Zy/ZImnebVtErqYYMh6ZLMtnqn/pCKWh37TXn2mjdj14e+cxjve8y9erMqSMDM
n6zf2hG9j3jF9bQKC4w5TAa/t/Kdh813LKSPlkeW1K9JB3Wc5OnVqo2/VvL08au1JljUBP1S0ykb
UMrTaHcB7NMEbccEt7C5nUiWnrDjOJiy4MWQsZiEUZV/L8/FEZ4Fy0UwKDLQisW08ioT6IXjrozw
ntscyUzcFE7LBLOiGRXbDbFrzBj8r9lLlE6a7nfQODenf/xBkYIVgtfHeKr+2QmE9VfYjW88s2hb
bY+9L9qgt25KHlxpHtgKsQLLFd87vmR9lCXZKH3JAlniiMySBczJX9J0R/pZ8IyZBBW0G+DoTmAe
WDvo3y7jb7jJWz1BnHQUeWKeCfMwVL/SrcGnM9mU638nCqSzMrMJWPiWlfVF9scm5mffJ76vodk7
H30bhfxu7ZK/RDCylhWzlNqEt2hNJWAsjwkaNRIZC2wA+O66axhRwkaNUrcE33k9HY/A09JjfXg7
KZgAkmqmuO5njt/kVjyzwBuJjpf3D3bNKVrBu4j74sA9izubGydTeOwSFiz52IkluWvUF+GUOUr1
U9JkJmMFP1GyxucxbeaUC5iggWBIvCC52M8MMYBtAHE5azOZLHnVxALnpiS+3RgEB5l745FvlXwb
A+2/BEf7wkcRqApI+1V0TmEWOTE1TCxz2jQ1auHGlR6ct434FY7nobZBLd4nmuwf6d1VMC9gOwPT
TkUrYQaREP4TEVOVzYdkQjRgWUZ9fFLA4DTsr0cRHDH5etwyXYREE/z34SXrSLCGYrKwF545uVBK
iNe4pfqJIoJLPtf1FFWCGpLZtrNbkdVdmgTza0z3K806ucxBQot0my/to3YHb9hCyzr8V09JprjB
0rkO4u8TBT24rZQBgIXno2OooAFmcp/ieUBRGG+r0f2yTHBeMSGH7PUwAOo1ISXJTyW8JAaq1Z8q
Gv9OEfOraGwQFLmCNG+Jvek8ktm31h4M4lLsX9dkQGPNay3IrCXrpqN0RwHThJ0jsjESWhmSTM3A
GeTmUO4QZYg8ReBbbuPriak5ckCr9h5dKTu6h3C5FN7K3p2LApnxeZe6ZQMIZLnRqoN6SOufwYIH
PAgzuvwJfDH3BPjftS9fYwu+bhtxnYeWD+w9QeP2U+EAR7MatbvLmaQn+H7dZuAQgW4VSfLZmgLp
c8LFt2CJSoBPuUs3Hi1p7CnVhc5Q6db6xmWlNTGhMFomqE4UVh8aSkhvCwZNKI2vvB/c/iWoxWi3
B9qfsZVzDAnuS/nxoEvh1iGG4mptpcerQ3EzLZ3sPVrKhbtum2pjur2PfWInyGq/FG/Sb1qBgQHp
DQUBRuelfEiV6AYNfJBCe6+jqoTrNJBXh+Dy6jqTRTo44jmHhJMKY3dYLpiMa7u5J8rwzZC2jXMG
yCnK2uwFZZu525gus375461TACzKb27ckL1xUPDg85dGb7FlDF1lQc9j/nOAEm/6wJ2J1VSleair
NYqED9JgovurYIKl6VE4xzuiu/9xScMYbl+0swIRJmIWKncDyAiUf1S8+aNnfqJbSIjHkT0Gtnww
aG29rRbRKqNWYc8/kimg9LYfgWnz7dklMwVCdM+gRLymE8FX4/XSfZsT99+ydery67QhYW81b6yy
8KUYBW+yLoy7/tOzpTV3aPTy3XuWW08vvxKO471HCy1Xoii+8Au/FgvtwJxOrvbkTe5ygPdfrLGt
blzvzCEc1bD1EEphWbaiVPDB+zaEL2L/Q1NGZSh4BUSFMh3ciH/4akwld8MiCXoVlOqYTF2iIRVN
OMhVH8JYNNrGupzejinIAO0zUMc04GyW9hGLTTOfWg3R4z01TvAykblwcWB0zUosLkkjebmiN3QC
sTPUzL5DrC8PxXvp6+sJC8XlPgJUkP4ynjy/jK5x94qWb6tBqv+AywAvgds/LJy62f068pbVtDP8
BaEZvYyMZqR0InfODMaFJQTkCM508Q1kklJq+v/MDcQ+KHoQdfbLB6GP95eLaWvBT33UATtFjvgQ
jF/DKFsrN2eymK78h5NsvZjjn2biwWYiktxru9p9qgrTLixTiz4eEUJLftmp3WKGf586rfw8o99r
YehIx0ZKwAa6OuROPeXh6v+Sc/JfAKswPhOnDbI5o5fY5nU+yGVm/LCC1pPCGQoVWOSAZqZnhkJe
E3aouP4VNjXgpvU5qQFDBLc8wSP6to9NI6H3LMVI+VE4tkW3ebWC6Zsgi2fkbulFb/j/4nJzV0qE
/6pPdWYBi8nm9fCqJdvfw9qRKPRA7bfpN1uEaOWXO+nP5ZPRZfNR7w3jbpJPJ5SEYQpjYcxJazPY
cyJeXzntGZnpl5JBpKeQ4Dfh6skAd+5b+iC16t+MixSVCWXYkjDXegz4Gwjzy9G3P6/Picc1xN7Y
khOLNUtBsY8hXoJrhBcwPqrulWdhkdsmCUK8JwVj/UYoyBQv1RRfT6b5p5GDR51ckrGhAZaka1lh
fptXmlDNiXMlkBXH/TSOjmfUzYDGvkGuJL7scLlboNLAX+ix5SgSvZNPjJ70TWFIGlszPo1PytFM
T+RpDbwDvL6nKby3K8PHS3eB7NAKc/wT6GC1jGULif2QxiG79Zpo82lPzrQd0hAkcFO7R92mURzA
YxQRb6RbryCPLKMZ2NhDDF9ZGoVymWss/yeW+5U5DY3bKLyjiEI9qbaCl6eZzhy0fVoCyyMtnin/
yjOfYizm0EI96czNInMKDVPtYZ3r6e18nsFURXpF2F3YMX5qsDNSD/kGaZ3Pt6PirxdCvMrZAS5+
HrZ3a+mIPFDpYIenQ7cJDhrFx4t/NbUPbhmd5zB+pzdjmOexpZkwch6yB+BNc0bYP8J9XnUzp8Wd
ZjESLZB2XBfXeqKS5GAydIs5PfyCAgQ91Ndd8zGW8IMQsJXNxZA1/sWh8mlIFaa8CEVc3cEdlXcP
K5+CW7JHy/DXNRJC+UY/nSFPhRAQxzB4l8gzVnP/2OhdjVKuJCo3W6ZMX7TJuaGgV4X8PPPp1LsJ
qelleKIWmQRQpK4OeQ3uvgfuz/OKJ9jLlIP3EIoxVBCfnegERY190W05y84NrcYYD0igFJnMfQ3c
o+uw+rPxdy8FFdN+caLrW6KJNqskHaxQ2MDK58evUI0PoCs4sIBAha3/8T2pNJan3wwyPa9T2dus
2ZtKiK8EJxIyeGQwqffHgO9HYSxAs8DHuK/aCXS5glcz2LyGcTfR/weSvfgvBTyd3RdiC4hLuToy
9fd+Qg9zKLUyGqwlD4QXp5T2v1Y660/npUrJAWJ9KgtRM5wLoTxfUrLxiS6toegDuZdreV5x9LkJ
T+ZD+bASNbuJcpqe/LLAInVILEizqqohSSz8pOEe1ULATqj+gnf7AoRPeEdlyjgyr0vneNnACSnz
CTW793vxi+LT7BG31KkM3X3+z1t6P7y919K4u5WGOX2QrwWx9XKyino9WXdySKK6DPs6lQhtWeG7
3kgWH+fgiw45B0hQIyoubNaum3jnSo2+lDW6fZLKCJ0K7YdSwopFZXZKWJD4o7T7KMq0GYQLkr+j
odqmixvFvM+lwu1pRQy9/JN/OwCxfVrBs/WoYqkID2iw+4DghXo9caHRxU4pECzV9FlBfZL9PsT8
NFX8hFgvrT939BRID/XmEgZCDhTsiJ7dySWqT/uV1TvWn67BbenNFt6HPmSotOIyDvyq6mEYG3fG
5sfGWucN9G3VEhUi+8pvyYGzs/77xcm7sxRqbvkXbvKehHDbsBVlghpNFgE9jso6zBHRhUsPdcLD
u8j9/Jhiy5IMdOfQ10YNBgzbJmCifEDOrTr/M2/miGysc5iS/yR4tQwsqBsrHcgwJFsgoFO14iOz
gtq+WK4hwWxwbw7bnqicuhGbuN+TXQ850KP8+jJmg7V6VZvhtA0w2N/q2rJVfR7dLLGZpQCSIjcb
VDj2ey2lc+pnyuBNMNpxgryRg2/5Qd9rCjtYq0dwG8sG+ry46LvTSXMdFz1CXQVhBRu4mrB1CCdu
4AY9+TWS4Isl2nG5JkFd8e2BUT3ZMETzZaaIptNHpdNk8w3npubFyL/j+EHX1D43OzJPLfBZ+HZe
iOxCEt50WicDZvjIRnS3Uo7CMSP1WfmzqmbrA2sL70CjW8x4wXJ7jPmON+Rwonf9tAxSA5EfxuKJ
DnFolY38rKs7EcoSJP1NS3b40jO6Bzg3vEbCl9W+XUtcZq54d+YHDdUgEm5TQd9SvVs8G6Mfk3vi
xM4jAt+scMldgcNZ6qwVx002vJqUlrb0AkM8hGwTKik2Trj3GCaGe+myoRqtWy193w3fP1Gc5rIL
qSIeHzK7n0Sv8vo2joIiU17+QUj2HqrCSKKQItxrx4xCdgtmjEj2/c7pVDs2YnXEscFvW/VvJNJO
hVcpngpGYD+35O8ieRg4eVyCCMc1sZr7WlOsCgIRX0JmFI/ZzXtcIo2PKlQ7WRH+z7XHyUTl8ZgU
frqphSQb3xGeq6fj3TLGmskzyCWy482exA9qL0S2rYy00aOl+QGDSbbjKrikCbBsIWRnViwC+uy7
MCZPGW+JQ7GiRnlV1M0BqmJ3C9bXFqlPyA0AOCJ1+OHm25/yxKUaFHjp/ikMh8cyYCD8WTUc8om9
Agea/xK6nXO5bkV+6VKeECC0+qe5UTm+LIG0qM6hfTOlVzjoAp8jmpBSuzmXdudi7YozJWyw6L6f
KkS6VmneajgsrNmGcXeXzTgUa4LhXlK+s5Vy77aOL0kKTpdTrcbBbl9Izcie5Aj6g7EIaYAuu5/Y
hM+kyw5K83CeCQkHxzaaGJGO/j1GOwxNwUe1vUOvA5w7Sm5eXjnfjmAdx/zBZWfqg6LOWkXnVrrd
mbWj+REtOrGXuWAP8aYWs40lMAyJ3P66ofWoNn85dqfM8HRCHS29iiX+iEcQaWmsTHeW5Z43mz8d
2QLRGPdn/T0vnJJbxMOejMrCOvzbVHvo03TYpAnjgZ4fq3Sy6kmd6cTkmkkaNGvqw8x8+7oX33yS
4dS+3g/EET62VoEzEji078Kfw79+B+pvvd2z3Jh+m73iWms28WDITUiA2VzVL8mgt7bQVzOMNqIY
yIuqUXGO2t/ay/nwtErPnlnRiUn2gal/JM9Meq+E5M8TbmQC/Ngpgw2yK2IeqowAY1BxN02rAknm
sNmyX4EbX+WqLAAkPifR6E5p3jHU0LKdiHn9da1Zh4m11i89qFPL8JBH4Tmv6VzyJnsHOCBQlYlE
GmoiUsE4B3VgRpaUTO2DKzcpxwODXvqqJyM7mZ9lZ+/yDFVWwqlLFT4GtsoNl2bVbZ4fNqIP23Jb
3BT+lE8AN2Rj+GYrgyD0nPyEnlBOK/bmKCS69Vg7Rl3/6gajE6Cz4jJ0t6TJcrsUGyqgsKSEFBze
g4JQm+ZYD7iRKY/2MMiYpdjkOselEgBBGFxbTI2R7mHPNxOa+2qbRll0MiU/wuy7fg8F+V8lQXxl
sQ52HOWtSloHKQeslhB/OvdySmD/XuFQnmsPbXCsev3MH7RIiSl5xa3NLUu9I7S1YzqTQKmzkE8B
/BsNk78liS+6rXjsieqyXFRGJM4424ob/we7hR9dF1RbiGaLQ6h3YQ6MegZgavPNqfcJW2DiIhYg
7S4olEip1GpRHB2blElxgTweWqVzeDagYsxZDNtAzobv2roEKOAl1OTd8FiiRIJTolPbVWt5+KHX
1tlmlpjoNO5H0+S1bjsRkLbCVMjqfkTvoSkGai8Zrr6RXX91y73CvGnzBy3QK7hoPW5UZgCKcYtP
YPSwB2sk8EzqRnOKfijOX9LlmyZ3Y9GYeTMAS/vuS2Vea33tZyus2tsHeGsxU2tvULumBfBUaaD4
mWdn+t13wKZzzQxTNoSs0jEFtKUqPdlBGW1FglwnhT0OrfNqufd3Whc011hpy4+3SCPCPhlj4UnE
5CIERiozRhkG/2KGyO6MLCFYPnSEkedmQtErFU1OLUmmn1zerte0g5Sny/GHEYSgp+SxZoClYCUV
31tZ9kETUfknPXfe89VuYE441Z7rFi00pk7FsnXIGXH5kdE4Oot3RoX/6irPhcxKjl21aBxgjWop
Wxs4r6m/ZWyqmROe1vHeDjacPJ9KcspqjDsfhwa5q3XsVnxTbm0sp9J/QM57OiD7odxfwdCbCCXE
rG5JXwcywQCp5VeYX8MyXdRfYSDF9RIBEuPwZqm/gwcK7VZn8X6QAtvUVHGg4HGoBNdfm9IQ7CAV
uQfAN/eRb41Ijs0umzkLThsX1/h0eOJFDWVpXwoxSoxT31HL5uk4N+3GGbyN4/LqXuxyM05YX7eo
qwuQNsE2nYtUHdOV3vZ1M2gr092uS7mM833mwR7iXhYCCcsGZnG9TgCWdcxrrnNgpVb/BB/16YwT
SHFmzYIM7Lmz4swvFUK5Uy7F9fhe04YZdb3A1aY0nXKws6PauCfB84A26wmsVdjDDdqsjzISqHFT
3HM7cJ8lq+hkisvRId0Oip4VWFT1iGAq1pfdEb8ekdEjahoehIq8m52oNSu28gw+9NxQZ50kQ5Ju
5BXxND55XSCDqMTCYJUD0+U9bpKP0SwdZavxs79CRSzftgj6MRQCjPykkMFGswzntdLHczT3HqQE
f7U8XFDSQpQuN4lCayRQoFiyjjZ8un7q5i2rK6wLX/E5fP7kMCbq/34rbgXMx1i2i5WzNz+Szbh4
FZT56oWw04QUtvP2+2bI4sZg6/Aj5e5VXdfq1xjvo6Said08lB7iv/XGRahboktD/RRPWJD5nEWv
G4HQbjaGYgMyhUuSNsyt6vokZN6tcyH0pbDGirtHvz9MBYlwk8vYslcdv4BaAtTVXpWGsUqiiIj2
Dl3bbKlMtzcWAxikSpYnTc07KAfOmdFaCs9oveSSjdMMUJ0tskxSS25dprz19nRs4jSzyjx5JizL
DCIBYZ65AfTIXPqTYH3SOGW91AHAfReDWIC32AU7bcECiGxWeoKAWCjqkRnwXMIzs0SmPcqbsCGx
7qIwuew45XHAiRp5GU1CByerTN+FZREtdEkcSNEErCw5rtnMAOXR+6A78NVWdTGJ4xNTHfV/hL9Q
7Wnr7PHC5cXrr+8LztLlzK+iH97/NiFWqHoW55jAJrXA0PqRkZlR1wpIxphztCVWbxWGqw595UOg
z6BI1qYEk7JyIWgfqby1D9Am1fEYp2fatTa7A2Iqv1c07ZV0nkcQ1IwAgvyA23wQN3GHO7reIARO
ttQUUK0DzarPqdgsLLbQrcOlYnvz59x9bfGkPYiEb1xRoUvJ9pIPy4D2LGzwL6EBZf/gywyGth5s
r32s36zi+RdoUeG7KFMC/HyWC90u1CQl3C5lNFgEgJmvpP/MxzVCh+8x+THZV9gfjkV30MRdEyvK
qA/A3jcMDEDFlUtGDdq/TtYHc59h5YZa0JM2B1lWyjLUx1vUVsjplPKV/uFEmMdnXn+qCiyzMCwb
996AAJNCRj8nCfT9ldKVqG93a+PIZ5ax0X6YoDl75ETe3jxhvaUiBOSP87PV+ojS/QQX5vAg5icq
lpTjPcMmoCFNK0Op1fFY6T+lMUZUQUCknupKn34L0/clL0tYVDbyOBw/HSkjPS/Fw3BD3eSVHJC3
pK7oLf697/fZPLqxxp0JyrLznOfNk8n3vM+AHM4KD9ouD138tqOzkOuI1OmwoaxrCbsi77kzoU5J
JuJmVmkurRcPybijsiP5Wm7knSHZeY+D4JZ+p7Ky9AJThKBKlWPiOURzQ55L9NxhPxr7yDcNqxtC
1hp7szXlAuDqds0YKmu111yXJ9ZgAeiV2K83zzhFKycQ21unOK68fodkwRDVGHDiuV2NiM03GOUE
3the/+shq1flNzZ9MWNzqEkm9x7Do7OLUh6DeT23TS5A8T6K66N0rU2nB9Mq8DdF6o4RaYTKMkvS
X6Z5TmkhmRAfj2DEtBQorNeiZcVNO4Rh3oi6wsdei6elUYvkI4quUAnGKwW7nAOpUOK7jdKhs3gn
LMf8zpVvQl5XYNr5lqrcGV/rnj9rKU9ONZtSrWh5wZPz3kjIY02rR7W9u1UDQY5Sd6x+F2bg8BGZ
yB+Pc1ZFT7tCWtrSRzOVZchUQWK1wA1MymLl7TFbABl1Pbq0TWDGt1cZldkVWT1OLJoKcubJrvRI
0/YylN8znQ7RpomvOWebHnCggAgyTlp1UCmibML++Q3U6iDrcDFz6X4fgb92jSVR1JQNlTQVnzg7
Fv3Oeq3LF16MuhcePbDA0SiPG6xzRPNHbVrV3yQa15g/yhSxcMObkVBraEnbDJek04YlsE++9h/O
dWJR85mSUBBtS9SWI1OOlITx/m365qzpi69Z2klCVMM4sGFJ6LiqlB5i3VXX/g9o1RAuXKtcSVaT
VdU5KOdPhFlIX0V3e8XLc/Ep5Aad8P++jicywAuU1xqdMWfO3mosEEldpbclRK/uBbBikvbiR0sR
GdrZWYst9CMcGCKVs0lTQ5fR/Gw9y2dvIIQK5fXbgtAbLGNTCOJToIxrYej559mnH9xSccNAahzU
Ytui4Ab43nLV4IGx24Bj7I+2t42oPNjp1zMj2wxTSGCW39tZwvLzIrLaTdvsleye40rHEPVmWKlD
Qsqvr5lWAbdJxF56kN8KzVB5dBfFMP64rkn0SdgOoCEae0PzqpSuZkHSdi8+lynadal9i6UsA/Tj
AQZzDfTQVtQwNIF4ugEhMSOX2gL2HiW01ca9IVbtbFLz+Q4UhAzsDyCrC8r9GtLD9Var+dl+rMfb
tt0uwYoUkJky2peqJntKzrfqJeHo8u5JwxZ0/AkZy6oNrKbmJNMRPWf15W8lWY17t7at1NlefRpH
TRfVd/j47bSl3z+NpBqeEhIpHfbIGWgFKLKZW6cENPkAC0GNiKPUbsYqmxxYxXq3wY7QvF6jx+Ri
gpF0cc1g4DYTkc9he6l+1SYvyTDyx2DtQtM5Rr19vM3AIqnehw1sCm4P8KoF6ddsY1Aeh78ysBnE
AkOchny1Is0MydKtlWD3ldNipIFWmDRmLI/xNi/GVft0pYttPhAB6tJbA7907SofMGTUJTriv/pj
K6hK+FYeO0tRY8ScGskvRM0xTD1wvn9/WR8kw4Y0w/fx2NtI8uUOuT96INJRO2ztJqsiZHE1UMzC
BCLj8gejtLMi2P8Snt9dTVAmKDf3KqHAfhN62Zrd+y+nXi5VZ2/i8N9N03oHcNQA7NcftLj5UaTE
jvBnZxwEbj29haYtN8kO7/h6LDEniV3mVrfR58prSq3TPSbedfn+96ev8PA27ORgShzwZDd5vAgt
sJ6yZv1mjgbK5pZhNotW4qWcQ1JfjH5frI76KUDEhk34uF2g7xpqt3RClMVY1qR76KYCPUEIO7pE
4EJE3iKIXpwkKvGkbwByXafSMQvcwe5vpeuCpSnT00/aKEY6FHxq39qNkSluBbuZ9U0p3StealmI
SNyhYgKVQKXoO35sLYHuLbs7XWC9go4UF99EzvMiqiYJyXKpfCuct3BZWGP+MfPeAJHqkLtrKoio
kBr6Nyt3XFa27ltJrPOcio7JLoGR1Q9TceqI++WFmLnbE34Ui5jDSSlNNTyh7GmCDcbsD2faQRvW
uSfk8MlB7RK3D+diOtX4OaWZ8e5q+nu6S5zyh3oyk/PL0iN3BGs/b79XJ65RGRep286DcshUG4Hd
Ipvyy5BkFgWZqpxpJB8FbgflWvB4eh1j6IeOBiI6ws0Ys5uvy1O67drI5Vamuiy3Y1rMSsskcgu9
p3ovSLFujvddwwRf5Bk6GQVWEXTB4Wiuj509zl5IgyphUVHvCmMezO6bP2Z8so031JhKIvFb/uLD
rfmN0V0vK4+X43Fj5qs9QsFXhxMwxQ/N10jJsxnrThAaLcT4v8Bx3qWc4j4oxh8wpMKgTwHKBjYp
TP5pXO12rb7/2v+KO2IP0hshkUWQ3/e3x8VEa7zqqsG7wl7KAiqaERLgnloDev0oitgarMQZHqLs
zM9/90dTZ/d6/w+U4T5OWDBoMvIgPawVx8jTBi86zlZ2Y2HO4U5aDrx4EqvtVMczlDy4y8f7EzgW
XdPQaA3g6NYI8jXCRCPI/eqPGdk8QaPGt9xWBdbG2UgJG2+waG5m1zDg8Iosx5dWMIu4e/B330lO
AhOeJOSDgvfT3UTxSLStd6rzzpV1U8d/JxRNrV5sIWPy+F6T6BdszY77X6mPvVXEvC0EbaeSE8VA
xLgkPvcJ+g4xuqbI/wg5M11J/j7Y2wC9YLnfqOJXG7GFevYoZ/ZVIW6YDoJQeu2PBeVmGE+T2b5f
zPcKS1ovn7vI8IM9/xmHIudO8vJ2u8p6uSY0d+ZzqKXkAtqERzOKpFZJyqadUE4wRQGaicAtoN1v
GqP6wDvdMq7//e3afX232HJgb67yEvFMuDqb9BXxzc0Xs6q5hxtEDMKhfiXx297G3qKO0oNt3qDw
aPxoO5+AiGaKde/ATgCOPZ5Az7yF85YMmAq4xrBflPzBIS3lk99e8/DD/HAu3fFm5IkpQIjL2+KV
DlNwdRmBw70rycDtxalNs3MXvMJquxj6/pMQeiouxMTkafK5w+ol3sMNeafnUoXuQFtpHSnFbG2/
1YcNgoR0nwDd0fi9qesySeuahNxiIZ4igwp4x4CBVV03D+xmDilJULpo1KYc0BYV89SpSa8G+5bv
r7SqH9gZIejWi9sx51/fv/Jrx3e3udVoNbEJEUSZG4H17P7xvBxS7vyorLG9i0nGmflS5PvllrBt
Ygxq+dTV7yLCUIF/UPvNhAaJ2cwO0a0dm+9Lc4uoxLuV4TYH8WR4hyVC1BnguXuEX6Ui6jgshaK1
JafLkBpTZ/j+0BFOKkBlzbGt45rGn6N0FthCoJ8HjkFkZKGg0QR91lCe134ZZn8RQoPmsybzTRmU
x/T35tI0WPMHhSv/pvJG0hAsPSoNSoX08bjm7beW+yVDAxbGcXYC7A9hwEAXjYhviRE8rY+sAkZe
FBIngyYrJgewjOsB+XwkrQP+vhsiRco5JS/+dX1QVgwxWZ39Bzd1vlma0cpJ+r4ShAdUGr9xgp+t
PZfel3XH+sKJrEWBJIEr9qmlxpmnfsWk+AWzu/allNVA9Av7wbw3fAZTpveR+cTZ7NKEHTiV+vQP
vpqwv//0RWN381lC7MFGOv12AXYAjqayMjRoTWw3r/sOr42DJA+yBCPH4818Ss5mHPrUvQRGRY0C
jE+Ewyo4kTalVx41UNNLEbPt3TRJpLENkmJsjE4Wzm7YsV6AUDjkiMGTAsxr0SoeWX27v88GVQvC
C2jAXFi/uwyUDToKUBs0jThLb4Xm6U/L5Bj//uLsfbBZuNDZf54OSMKHJewK+EHYXARBelM08N8u
fwfhNnP6x1fYUw9OVcb1I9YvmvtA6vXhoDLXgZ0ceM0qcrmxlwwWUvDamxbBgL7VuSODEnGMtVvg
tsjpdv9e8+EXXb/FJ0Cnrurg/Zdhac8eyTFcrNAsyK2a/pnxY9mL3f7D1INBYcp9oRBXv+uWRli1
Nsfjds0dEE9PLGmrGj5ERrCddiYWym0uSwCyHSdZCDXtn70xuZugPV5HVjSesozEofdlwBaora9G
ueFhzNLXbRr4YFwzPBOoNcksy4fBukYqW/du7pHBRn6jIE0pc9a7OrWLwsq4bczGZ7JfzVJC0/IR
dur0SbIhk5Szg2/Qb6X/fiF5Gf2H8ba+DX4Nh356jPNQNJm95t5LAlO6kMKK5swGdnfbiSnPQM0+
7nKNCozZMgqJ0vsPzN2GxB9nPLQA5LDREEn9/OcnZCs7Ejl1n9nwTZG2QY5eCq2KfmPSfegCz3OK
J9aaSWqUiu5EZhH+yJtH4m4XW62mkTtr6n9Uz4wD54VJ/j/QzrS+SBsY7WQSr4d9qL31u/qYI8qX
qTHhIgcPR1PvfIlZwuEZSoR6L8nvgTeBBthyoYpGN+/2r4HF2EN2+yyL3jIbXMWS77Y+CbxI5ioa
uWCHhM1nwtmDYGSDUckKNEwVmEpoyN9/2BS+D+5euH/DV7hwbsN8mhmmRY8PGvdMYMea545ft5Sb
Tux4l+SoPiHyNwGdMbLM3d/x9aL4FZgPVQh0qNKP3rI8gUXqDSha9OtGsev7vP9+kBwCTmLb/trl
yQgTDUk5IH00aiWOiyH2ggC37avscLvyNV4oBfSAd/IQsNBm8h6UqU2Rc+oy7MQrmyxbBP9xjd8o
/L+7JChU2Mtz5UrOqRfZHkODr4lde6lnElEMFEaeTKsd19APbK60BCc3JltU7Xg0g7MuDmfu8J/t
Fv4zpYYBmArB8m3zOee1BV+wBKIDxR/WX625eW0CxvDKaCPhZ/y7zWF93q0HXna9tkBCBxs4iMD6
2rgKSFSsICAkWP37jBxyfipvFg7yDESTZh34AZRA2pZGcOiGsNUqLl+amEEkVJDOd4SYoxcaiYFd
9kBzxh0KP/7GU4XJ6WI9kybtGidiUxtLZTRD3lZ/q4D92UoFlw0IKTV73mMuMCu83OQtWj5NBDLl
a6W3fLXlerWTriJ38I1gPSxvx9ZdokpSRhpJXCl7J9xfouff0hCOEqyqGSEI3yHzJcJI7XNEB/Oe
isrSDrG3y5rKSvJbmQNrdZHnFFeyG6K/m9Qh2Y+QfBFWUZkv7GNXkqQcexmIrLvnLFMNwSKNgpd7
peLlHREOXXdmqaxprpxhlDwTPZ9YSAhpGyYu3cRQaGijaBea41OFmc48Ofx1ZSSdlTqGsixBcp/T
o5Fm7kSSWVyVuYkhvQhBRtpa5pxG27UFaDcvzrEEVW30/pFJ0jKnn0jdFPtU8FGB/KKg5z4hPBNT
Plmf6KyFaB9QmLFdhxUPdcQdAyKzh2VN9zfBLKb1YtkqrftelBJo4bKjscSatepoF2ANoNLGrzPv
+MAkaVo82xylJlRAMu3bDTIFEFimoLSxVRHtk1wa+lbFBPla7cdgXOq6+HHgp4LH042cbdlO4i5T
bAlgfmJzwfM8b9W20g343lvvL01mnP2WlUEb7jObKIysQwBbZnNMQUNze/q6dEy/71pTFhP3YfpE
mBd04lmag16StodzLFiELxBlcRfj6bLpYaqgqzAI4rs8KtyQqypiJEGIc5RtraUeUYSecpHAiItO
aTFjjZzzkD31atPTvyDc0cXSDDQsPRbwY3sxG4cGHPARG1BEyCdU04teFzofXv5RW+K0T1bPH6XZ
QeyegJ/RtThXM2QhOJBPUAqSiJpio8viEhscNXai4biuxm/Ykzf/lXnsvQvNTNLT5L9y+MCsWRzV
3gArGjlsSOMdBHiBV1/GHStzfI95nyEdcYglwC4O9hM15lLsgoFcRJQax08BFmH1lANx97KBAONa
r/cpziONG+iYG91IgBbLUWX2uTb7lFAso4lL57uBIsgMWhUbH7Q7TCvjdrFskpzwBS1qP1GFVII4
I7o07xlUyR5L1dPkS5tBDcH3/o7IAqMBh6Ms6R0OWMoFTuwoTWDWNHUgkZiTkiIXFFmeFOOOrfON
TMfxOBqh3FCTyoJR82QyfkfQ9+KJ0sS0E5UXsFgS6mVFfDm9I4L2JnGHXP5pnmXdswzEuAil89Tr
rnRpmaPhoFblclGQ2Tf+abrEkuQ+ef01mx1KTS0G+mk7J6YBzxL426lvkR1WOtu/R7B2pWmW5gIa
gNn8yPBxotkNe0VsqiLhVJufwztnoGxCXPbNmo6Cw7Z2lZIDpWkCqnnVAeBNSt0DmvTYJfwWaRWH
1M/uP4Z+GpK7T/jHeiz7ct50cw4xBcH9jA6fWD0aP/vlWp8BRNUXos2gsATf9kmGCHPEKED9BdUN
Xj8pesymmV5BEakL2RmKQpnb9UuoBsHP/9wCQrQZqr7iTdEbBZySkraG4TEh96av9TcNDYocCb/a
rN7zq+kDYvCq4ur0NAAef+DsAwHHcyHVqblCCuefhjn9aqLOkkwug1k4UR7onSG0ahHXBgrQGMFI
kny1iWHL6urO9OuuDR+8hJViR2/LJPHfV7Zcw0LcNoWQa8290/8lwEdRebVZjSoPALzZKkCLGCyh
Z8uvAsz0tnVR3O6sKfLxLF9DRCKvosferke8GWmgcS6j9IFyXyekCQ3n3MUqH7sz+O4J5PmpBwSq
UFQitlOsgOPFmDP5ljVRcQ7N0GLx2C6/mO2v5w6uBrwMFeS4OySPqrq4W3W50KXPcSYRIjL/F/hc
djxC/nYmQCerXg7tGFXAQ9B9an//rgss2o84oZUMGaKI/YqD3RYNACHYVVxJGdOmvMhLHak2rnqa
+BH3dLqOPWl3nj3D4+XJD2AmZvviI1yePQCSGyd/SAzZilGFHapId9qWJ9srbzddDO40JuXbPRLG
klAd05ytVp/3/71ilYlxLXkUIAAN4zjIiEy3XvO6eBKMjV6WJlf5owTTMkS6qvuIzbvxkYoI+VxD
VhEfGR1/BGl0Ptwzh6ky8wh3/uIGH4yf2C3ByyKZtmayC5yDfN2y2vTwVh2ya+7SfMQPTIU5HvZ+
CbEiWPATBqkCQdtKegLGLprRfB7nOx0bJP3G31DFHGqq7ThQ1iGqnS4k/GGrPckwabKbuOOCH9fd
4/LcKl4jXQMcNMoxp+eX+aKGFB77zUblGHfzhlG8wS616MVd0itra1RjDdLp9Lixo7GDqcijCPF6
0aCsL/9UhPj/mkA4Ek/5eyYGudZnGArEfHlPttXoe92fAUc8SUT0c5rrnPaxz/Ye5QvmfdQxLvnD
Lvnm+QCGSK9oOZlIDBLeNTBwTqptCOEdkyK7/xXrfe8JHzRTW/QjeL+hVv9GrybJYLkmiAJoTA58
uUhrMpmggV3r5WY6fbQvq6WzVcppgEK4S5RzySU6+n62Ipjx0CJM/pHZwK5FPkYOifHfN+0fL+Bn
naEGhSEUqG50kqwMIYN0oN7W8llpM4WZSnNR7R960rC80OSTn8BdCdhbfFC67FREiATB/C+Y5inw
q+Imr0KgYzqE44oQ3q0Y/lkeCnRSXwKlBaWAQLe77QigJtBH8hNIdI3aCj+Qsm7yzvfG4JaP5hRW
enNfIOhQqAu1pMjiJfiBvObqMPGj3Zdswo2gWxxF+5V8kl+SKaW+ZpU9D3kJocfQnQmIS1RGibgu
hENtpKKrsBSG2d8qSDDf3H14YBJjlrY7oiyiIzc4iAKIRUg6ytsWGrb1n48rKxNeB7t3WuNr96cy
MX9Y+PiBBfyUG/+El8tRGk49Zn8J1hY48gL4KABhdGmUrMIUxepfplrf60u6mi1jW2SRXAzllcCf
+UM1EHxbiO6HW05VzniiKYWpVsVKU9LXrTGg15RO/CjNJ2bZcC+v+l05FdS7GSLg2pzL6HRlir5d
Gur7BIuqmlXA6S/eG7mjr2fiCIiw3/avC54u0e818a2RRpeCuy6W/dPpuGy6xP4GRgStzzIVGT6l
fv1vhbY7XVdTDEeG9h5FybOKHwGt5fIsIDS6ozjq3rj5OnJvhInsBqNXvvxiu4vxoS34snA72oyl
0+8oXhlBup0sjFaru1bXxPv64xBt0F+q/vOiWdRNJpYRkqCsjTrUGNL0eezbf+Wi8p17awkcqGPu
JU7CC7l7VUHHxDINrWb0JbN/tln/NOW2rGifkm9SdSecVd90n3MA4G7caVTIyNSFa3F6WdPmOhXv
8N/YzOAiw8islp/wsMguGEus13Jfz0AvBu9m1LohD/8IVSr8/0Ll69ayvRh0zsHsUV0bJPm8viR7
fuuT7/SDyh6C4yiP54IBrFWE5KjEoiHjZakxt3KN7OTbLV780ZBKwrGbQaOtR4oJlGu0431MwS2N
w2+JV9pdMn7bUUucLQU3GzzfLu5CuFgkdDIg+0F4UQYYvaQr8KrFz4zWJ+K34jxyu2f8w/J35MIF
9pyVsjNmquM+Fnt6rW67mB7zXCgVnVmAz6IXbdqmm7tNAtGw+mq8VJfsVh2mm/IPvhQwmXrie4Qv
/ehWPYuZcDJWPNN+b3Q+4OgVfFE9fDY/SEAIwYj9eJnmodbMdpa2GjzHpZFBqOwaoPuYEvi5+hc1
3tCUo0PEb4F+scOfJCpMDAhGkTsX61qHV9RArIsuTyx6PfcDFzUPJWCjjo5gsxw2mvVMUqq4syXJ
x2i38HdK98p3pRqg02wYCdfkjEF6uQznC67NdDLuwnCA1zPq1UTRKsy+ccPnhpvYQ9+zEaz7TNQV
X8YEbtAeAqe6wj5ulM8IIGJOhWG9LzoxzMUWKG/DSm+v/m1aS1tyhLXf8YYN/de++lWCqfOF/SuS
eaQmRza+Sgpc6XUGZZ0AmuYIquIL55T/IgFTuR3+WxhM/FPgbrULgf4RE+4242cL0KFIjceTQZUX
t5YAVvjusAboR6Jl3IFqKwjkB6LYshz9aKWefYIdCqYMRasQlEK0GyFzSCnNF1u+xKLo0rMxqpfN
hvwFxddNou+YDrCuVd+1/n8jbqm48bWc8eJmg7XwHrzMoqLLPqlEBchI85bp2RTFUs5XsZukp/yf
Luxurjm+JwdWyzsRu/xIrczyUdPrULPkNoehJAqavc1hjFS9nMW+jth9LGiSOVc9r7511RK8A5Np
CZBoHUPU5T7A4gt1idLtHWCJrZ+M0KFQr+ne3F43k8dLoPhAll3OKZz2ARzIs1mG0x0r1S3BPOTo
bh2SiVdIom20oLL4OWuajwOUji13mnSup/MmJSLIGme5M54HBYhkBxO9yc1rd1iisH6E8YEfpi2H
3TXzl567QVCGcyNEECC25ydik91iOZ/5H4nCuVmIDVBNVxg4SVHU8O4dPE7TQPcBiQkYUiyvFIDl
BcM1dJm6dfokjnUlfwlfsc/2VOAG39lbL1Gnrlhv9dYeJwmXneQZSDdY0ml88hg1FHbBQ7cpr1jW
JYkHkY3JV5wyKApGgi4uS6MGKBtzcCZJSap+KevAI50T6YJDgrO8ikoYeTx6QhsgqKYdQubTS1XW
uh17ONQ74mWhVkixcbd9zczI4p2u0nvkKUwqMrbuQ/iE0cRBoddClo2XGwveFIT1oswR3q8PhO/W
Tjy+HuQjniRw/nwlcJN5u937cTTI0VeavXw9Wy0lBhIUD5m0kw8H4dQecdskUCRkARDvrE870SUM
RIidUjdeJaCHiT5+IUZ1MVUli9hJjjL7eYCryNaaftkBBWP1y3QQ9JLTSJFSuYsNcSNzF4dmzb5i
oITxQR2nebOTIznkx+PSw15X52owUqUC61EsdcqbqJkJow0wqc5IF9BEqkU/AkUKs7vxYVlA82J4
tcCGGzk1D+DPeseyYRBwzsaBPHN7aBz7xTTozv/pTqT1JCVtt/kG5jfODsAjfyO2ut4iaUY6HcoB
vQClg6geReOGmCqnXTvIody69imlIljvgsMyehDzwJMQOYF/kV9Dl5f7uwRC1CHiLV87Nr0AYSMX
8Sg8bvcN6a1W6Ynpd/MMj6L7aUtddOK05tPaUG4L+pgY+874n1tXRHkAvCG/Ni3EKktLRvXMY9Xi
oLH6c5vy4bVEreG98KUmPCt5LRjtEu/+9MYEgbTmNtw77zgFD/LUClenKm4GctHGh2NWdl6k2Xyq
3P6ncif5FQ/5U727pYvBJCUxThkL2nEiiPprsoQpdTt7jaeAtSxTqo9X1/zbDQ0YhBN0bRY/59RR
XhwdE40K4yySQ5PjVpT0i1wQYrpuEKeszg6k89jG0yP3Jnx6pQAMp6uQrLCg8jvyS8hRt8aRmTo+
/lrI3e+B/FkmpZ0MpO5X+E4Jw8uy3Ckd1Aj3BviGv2a7oIGVZW++LSf1u6tp3jLUfSOqBaNjK420
UCl7iKlIqbsU07uEtxw5M1RelXe/MzPZ8aRwRFzI4klrzVJuVZDHVkjwhMCUYV6iWNSgJkcG3fRU
zCGbyvE9NEUpAon87iVucegvQ5qUt9CibrsepT53jfFdf6SeXeU0zrn+a9hcN2YhtN5Pd5e1Anmx
GtsW1a0bMfynaQaDS/DmYhIaqwbZ0IlIcQi71pSguhk0YmDqA5XCqS1x4udRaCurpH2LIluR8mV0
WP26IeK9PqoKSuAGZcfHMLHWJ+wHTCwNaeop+nAG7sY4vsNpsffBh67JrlH7JXJQEv+hxLZ5DdGq
S6JA7YUltDYeY8jgpLSgfXx1ekUSNMSinzvUHpZ3NlysCR3nMMqh+ZjBV/A2nLoh+QJpCXsLy5sg
oO+NUKMzj57iQFpkVVMnTkxnjuk2PkgKGUlaXbK8kMo0vTo2/6PP7fGmgap3it7mk78GBV2JgAKI
y6df3ZWn3awkbY+fMPZ8wkqJcYA5RnBfHy4IYi8bV7fhq5bDWC3Bwj6XblUK2psyfalJtT4pdCGP
hZyfUH1tfA6s1FE7UrR6wdrmZmCsUSSFQ7MvRHmQfM7v/G7oBA+KQ7k6OvMaIFqkBId+vJk/we5K
Jk9fOsM7I8Zn9RlYh4KlMWVSPo9u3Jh9WzIrGboAu8Az8Hx1lvxbtNKrmoj30UjLOGn1WWyfeOE+
53pHmcocBOUSjzkNMzwIt5au2aejFv98z3C16/uOIhl4CuZBr63tT3rJsSlgasyXzRxY1X+dFpm2
cOW01Iw2nIMkjjf258B18eb1/4nQkOlfeAjGHTJIwnIO8qb5gzQlkS/qhGAbtauBHZR/W730utzF
Vupqdpytd8RYgkqVHfIOiWpzUxUbbIYgyF2IrRZgOeY61NXo8PgmZqI5TJyx/JdjJ1IoCp+19Fq7
INOe1IzRqZUT+T8YfxTq4iuob5SUgg2qysbONa2SbCuxF+TQKzOFiCFzAri0hg3LNsH1ldLtpYPe
oCHlLNa0HhCfxzNiwl8RT0BgiQLBzqcwPUZYOBnhRJjIo6WLzK7L0KS5+oIguV0kTgsAtknFa3Lf
zLQJfvaxreBmRlxx9c9X8jQHi/nDm/MDGgzUQWwWC5ukKc/DTucmmvBJ6QMwXDIRDE4r6qardfmq
Gzb+UDkQWGhs43+55yTNFLbRh5cg76xhf+lisNziMhDYNThbfw/gAlSqGsZ6BvFAajoouZh9Q5PD
ERk4YXs9NRXMLWI/F6G8vkSkmANILUjd7j+xEHlTpTsUFbDJxJsm1f85At6FfGy9TkwDtm9tIMU1
IWgNz/s8/rz5fxMsYKS9yElEOLKIG9sSHUDQBkUlowlAeMJYspkZ6bPZ9ujayJI2FzOxdXUf+WZs
hoL7NfTwLZAYSMBJe+nlv0WaLiP5pMflQYjpFvJ8S6LSSAw7mpWldjEwTFNaKcF0iL31VeWwFliU
/fA9gHsAsbFm8Jg7w7emks73I4libFeGm4ucdKgy9XZ/q+E1ONqHS/NysOsIa94DINPd9d9liGUq
kJikdsL4l6/rOgB9GnYn9W14XMkA7p2q606BjmRgzmACTtwysrJGUFcXec6wkdBGt94y+1Kv1IxS
zmr8sVmpoAjDQ0M0Hw1Q5fsTRLcbz3aEzSA2U70LLtAXwW0xye37v1IXAZdisdqJvwg0ICUqy2X3
a1AjHafewu2//Ax70o0A7d7/nLtbmDDPzIKbVith0lVIaqjzmMm9TlDPtqaNWztNTzHsBfQmxxH2
jfJFmxWUG1Grj09uu7TqYRB0PvR+AW2z7vsxc7A3ZWcRR54sx1tB4kmoOCNMGAq1i0TlQEo21LMk
sWuHVtEbHzjDHyV2gOOGwFnsVBaSOAshokrSg4Il9X7SeGJib10/o23Wkd2H2eOMtpA3YD3pt9QX
9LRiB0/nardOLrpe0Pah61Way3q5aavQbrUrPto1Bb0m6ZW3JQNBLrMIBIl5FlDrzs2rx3trByqc
QrIu1EamQvxPHwIfK8VB5li/gs8n3u8SSy3IrQLrAcAzQ5cMEP8QZOCvj7iWyE4fp3r+d8esBOSo
7iFmJH12ayUp7BTsaOiluqoWbMur+ZxAFf+eroMc5yZPeVS7wjK/8Xqt6vVBKENiFfa8gGKDr7ia
QJsQdCMcLuxyXA5nMhCrvR2+igaxTavg4a6uTIgASocJEj/rL/DODvsHhN2JnmRWkDJDHOnjK8vJ
e30LZzo2cs6Rcsa/PKMe6Tex64pM/rUFPeYbFweWpOomLSrB4exf8IY8+8YSgGQtJLPf2wJksSxL
gMNMP7+5eQ21j44PUAVz6+9xiXZdYIkGeCaPwjlo0dA5HLDcehAyn0KiRw0vF4V5Ydis/m2SOtSX
aAlpckRWUzAF4iHQ13TJuNPnopYhmNYSbDjftOLzrJfREra3/MsWyPlljkkQATyq46Qvjev2klBt
Tv9dO+KSoCqjTy1uFLXt2BdI5LKhQI0kWsDzAvX75oPsfKZcSGM0Wxk0SZmGAxIP35Pp6herwxMN
b1AImWGXZkLUWC6AtQOfhBthd4Zsg2UsIAOWR4r57f0c05mvMKWu2XD9Swt56dvc0JKHccfDMTjj
N+GMJeHUwRFQujyFtQovHQtptigze0YIvCZMZvkieYn+ROPFr+SSN2t6/FkGZEoM6Vk6NNRDZjr+
EaGfvuq3Oxaxxndv6yZlH1qDJoPdORh/fokvv8UHJeUbJEdJkVTPAdvOJQZqMn8fK9V+Nmrkn3Pu
H9IMUz4XABG3rAwGLtbkoDrPjlRJunjwIKfJnPWNtmn9sx1p6Gm+V7eeSKJ0zxg6ksKekD/3siJ6
+PjXKxUwH2p7edsB96xktGyP0loYWQDRyKGRdygxeNzrSJVZFLDE0Yle6dqIKzsWRovlIGF/+D/R
Pt+ADCPx7LJ5WafkT0urz8BMoAxMCchsJnS3IOgOc1bXt7NjBts7Ioiiqcd+MAKKq2ab4bRabQO1
951KfmQfmyBFkuOq94fA1PwAvA7DZxEAuhAT33ch++SpZRYDjkh1IbKsYv9DwHV5GLn+4KGWHVR4
ofQQM2cmauVpJQXv442X2bgusH1va0sWpfgSj0y4nP88MZgLuE09gw38Vji/hHl6SJz5ohko0s6G
m/jrYXzdOK8P9BTLvu7dRSFdjkbF+P4nIAp0A8czMuuO0SAXvayQfqbEV/j+9iJsWRV//C3kxjKO
cyswYJUEzsNa75X7R2HjCohJeLyS9mQD0ww7XEKCr+hemr7kz/dzRG0R3+1u/PlGyrBPshDu1MEy
EuL1HYbdTlqqTJ3U3zJcwk/HdLkTKCb1Ixo/Hk7IexBwe2IPqwXewSNVVo2qNu/aQFv6AFzZV663
AmjEMzenTiXCO+FIH4iAvyIB8wFGO6O+1LDf6kOJ3dBsLl1JPExgJ+djEk0NBGHczd9b3s7afIJr
5Jv/jBVyB3YIsesZ1JbEZYwh8iqxL8tHwpRUnitAyHLHJQvc3rvX4M+sncT+fcXVlDRzFBu1lHD8
/pX+4xJN7CqLjiHWemZZb0aARN18F3xbiliSixC/zUmUC7mZ98YA7RJ6j7VtfoZkjtTwcdj1Fg1P
usYQxAWW7r5gnuMZ7yM/YJpeE2RWOJjknKxWyu2s9QR5BlLXhJWLbyqwe2zv7kmZSlgTrXCMHUHY
X1lvJTjZfhZwZvXkapUPwzxbovXfdURPFIfOODe6guNVAFDq6b484J7NnlsgqWCpDVZ+U+N4ER89
jvY280+owW1xb4afrt7OlnoGYc1EU7ce8TgJbjkNeoll2+wBX5IHZvRr/rPnV7hGzhHbSU4JgW79
phAjLZlmXyP0o5/lJgoUtqbVj1rSTAiPCPQSdA49z62POwAzXtNzQenj0ncUXflJ5IgLxslpHoLp
ZJrFwS8uv2DJNxTMtai+xGfHwiQjzDitaACv/qI6dfg/8w9M/u3NTCU/AhlsCj8Who8h8MBEVLh+
prcw8SV8Hjz236yCrBq/ctA75JlLEwSXzfXPhPp076OOKfSc6JYL3xKzf2A0nNw8+WhRI1rkdiR+
TVzR77+GR0U/BsWVGse8l+FpfuGtTDUxOfAEzpmoOc+MNnma6AVZUnKyv2gcmz7zwmpmTcVvEdiR
fr5WtT/ePzZK2n8Ul7HXkNidK9FWnkzvybN7o3k815YMEirk+yCYHyuXaDBOmRD56/QkYOqhgHdY
UMc/SAN+DZJCngAUFCb1kT1z1CGF/6/v++5j3kyfjiuSUbbAUXu3eLW76o7D+C02p6hr97Hbcv6o
2I6sTRwAbRzEqtUNvClbDoGq2svpANlkHWU8/DIm905d4nGWI5HvMugmVW9Aku+NMUOQaH5719KM
NTEmlarJAYSthFah68RGDpHi84HlHel/qD5zKvfpmdj74bgVp6l3kXypA3HsGOGFtrf/fiijdM8/
GVi5SthFhZY1JXELjBQqSBtwJ1vICAvpRQy2EZYRKIbfriGzK4H3d9HefIvm5nZ2h+8zBI/27AvH
72JihR/FZIqREJXg13Xvp1elAyWcKSnt8T93YTdkJgD/cpt8v7lANoBB9wOGCrXZsVhpMp05dzhx
eXBsaHZcFkP5H9Ox+IKFjWiHhExtxhAPjy606G+xULgCWx9pGzgdXtSRGy8sq+yJhfpEMw9PNCaS
jnMj8F5N8Q/IDEwae5AkqM/ziYtxDGBhHxMAsX63khLHLGh9xzmuBTldPozo0ns1nRRI9SbmmwzN
HC7bhAH1f3TND4upTsAbIAwXIeTdxmvIevmj3p0EkTx4upwo3T2wz6lNn4duWUcBjf5rlZbNh2yQ
stkI83hOzgr+cUUJgStbSp7SlxABA8xyVYHgsLqmYw3JFe1T2HudxpeytnWm+2J2S59VF3P42Lgy
1B4Veyys3cQGpObNwUrE+Q4b4ZNe5+SWSXLVlxZRRsdaETI4Ouux4Hc7XsE6J15tUh2418Bb/JOv
JJOapaEjqjDEnY31SmA6Tx4kj90c8VtrWWQuhtCNcdPKhcj9QxHmIZLxsmxfkcB56mju446qNM6i
OBNHuQPSRmya9tXzNxyKOBwiwZM/xrtNsI15v9SObwHcVYBUWdZsCRutUhx4dh1SBZeSWoZosIbW
0NLrno8Chmc/UAh1MX/vkZp/GTrC43PxB5WqLlPggRWpp7OC2Yn616eMWzb04bjM4GVK6x37REOq
Z67nL6Fd7H9maSXqnX/2VnMKqPEaWBi/QOF0NawOOAm6KhrvLEAr4Ub9ZZObQ2WhDT7wMcJSkkwf
zyHnUBqb/qF9twzTCQ06TWIzjKz6Msv8lw8oKD9RleCpOfNhnZ2lNqPMNF8FvA2X9ncRmFLwjTUq
mawIuRvaFx2gVgON9K+Wqf99Q3j3kfAMslT4rvP39v5VhnIiE4ubf7e9XxKXhanEUX0MqEDXSs6P
W6hYK+g4kMEBlPGnT8vYu1Z0e8+h9GpD26AQM5kBjB1rjIMfao6VdtlYUImLgXSlDhbn5yZFnA5l
W6xxwYSV41ncbed/Tw3sAc4SfoHhkX2egS8jiWzVtj2E7H5VeDKb343giK/BboTSid1mIMfr4xkN
keNm19GcPXOUlwsU4uJo8/fw4K6BZz9vGC2ZUbGu/kxu7bKbJxF0/KT8UATH5oHhGEoGm+uqiJDY
B+rpxU2hcEKZMav1Z0tTZ4q729jDepovKAuQRqDSyWdjd3P92zr0Mb4lR3leLUTCdNUqx7UM2rna
yDW8hyYegQYSEfg/cRXwegpGlHzPmPph+2FraOFtjIoxJqV4T+0zfgH4gb2dHM3FyI5K0K1pMjQZ
qEehWlhrfMctiKD/5LhUZzrOmjfkRizy9Y+Z//3/heKty2an1eJueqwBIC8n0arky6U7EoJn6Wiq
caIBQT9bmuv7VVkv5vmGpjdFtu8nrUrau79tnDcxAb4NNX6kVGWXyfe3YWCizjIBgoQRmv2+LGo6
FV9inX0ZIqq/FxQVWXa9LItnacDl1H435lljrmsgdo1DTg6uxquib/felzBwFFazGEYcRVwtGHHL
tV3OwRHXNqzfDFLvWRX8s5yWhTje9pCx/VKaClsQhtcxbOKBe7AQTuFvoSu/uF1lBxN3lGFKp3ne
sFa434NJ8fccX/f8IF0C1OQlMBjNdg281zz2NY+d32IpgBUssE3BoVb8R8zscuJ1TMgkclJI6+5k
PZH+FO0DwlRrg/XFh1IV1gzoAuXkTtdFyvAsXXXNGipjAPubTSJYF0RPk/0TqbrsxR4A+7+ygyGy
IdxpK4AEZ8FoO05SbQnAKrimaOSLuSKJq+eQWn0Q7nJLjSMJcWR0lItPw7hANc1Vv/ZgzvjS11oX
bvBrI7Ce899Gx8HyQPlVKu/Bvl8BASVVh0Ey4CUFhVzoha9cLmp9WKFRVkm3PSZpu9X5N/URLIHy
xTmCeTwV69iCzRq8atVxLKRH9GiVe1e71JuuDiWmeq8CAcnuC0OtuzAxPby3dc0zNmSujMqGh864
HgYoQFGRAv3Q2jQAd4mOfhw3fL2cl9Q9TUZ48ISxuF3YSZHsmY6VufWBiTpM84RCUD7t+E3wjZEF
+NHoUWwwQbLKjJFH/i+vvqpzSVCL0ehhYaCWkshhGVaTsMH+xzei1Jc3x8jXuzwqMcCwn0obpdgU
fbQnu2j4S46dGNr/56p9S73+a8BdO13tHapeFQEvCFTKeH3L4UT9mfBe9bcpix+G1R4P/2MhSkmV
OF2oGHB25Pspi58YFdSsRRk84d7sJujwCD3BMPFV6yPanyCH460MraNUbNFve94rSz52kXKjTP5T
nNcoLaX8lTkjF63eU7XrG8mK0m8ZzNgS+R2pRYpisTQbyOBFxcdhdqHehFxz9U6WETgMKgZprniq
gDAvNfklTOH6QfblvoAGhpTVSUofqdVI0yHv+YfNSYA3GG97aaT0nfX63Rn8odsx8XJLqdGI9b+C
do2WM/3b6y0a0CUh42/acNISwp88WBvqksJl9b9B2TRsvopWdurg5jZvI98lrrsV9wDIqeq3Jti4
5UyLK1M5SkD8xsA5XSM2TUeWYhUQbSsvJj5EiNModSuq8lRNCGvWuJE4t0HO4sjYiW3Sx6lBh2js
Y9DCBfqYzYG3AIur0KyUZBmjJd4rLXyA0VqUCF+/ockyQRdgkVQ2Twvk8w13AhCQFZScvEqsNrT0
Sq2TLJFgNh34I8otyzfMgihqW1z7WqxaUtzTMhvGGCzPCQ3cPVExk0vfTDQx0ok5JddEpVv6tV/w
qiJGNPm2o+CuqgzUOEwCJu1ZeZtIEVpR2KGPBVuPYP4s6aXgAG/Mqd+hN9+yTKgfEdmDqRze+BFo
Pz3oTVeQBOyaaBLKKBBeUMUm2vOe7IWffnGsKNkHfPl+ktt79I2p0SUkRPJG2FArutMryJYpSGmf
tcbsCkO0npn6VFl3MU7nOEf91ZPMCe3scL3u0R6I8iZ8T4jtU8MU6dDgpayHnXunCY+KiztsdBMb
AUh4868AzHbqFCedlAELCrD0mD95VysSWNYVoRjkekSayDHChLjoZ/3pXaUcs7OE9kygO06021ck
Yr+qzBoP3r1yKLyWv4Ry2LNzmpSQ1GxDvfTGeoG9tzapHJiN+LgS0pt5p507Dlozy1tq9qmUwyq2
QXR+VrgR0sEWk+ClBvkzbTsnLrZjzT828QtB22C5umglNZ4CkyZ9DdusJhj1oAFMRSWCt7rY+UHW
Cj9AXz9oDcEMjykK05pDFab2u5SGpU9N4TzHZ5lsryiLT+Srs3BGiuw/iHdtp/a32DsCPs1sWL9v
UFJL4+P5NbGe2dHiZg2i+plMgytQEb50kvnEe+jtcPJD7U2rU1/8KK7b4904IxeMaBSKTitNijIw
bpK8sFJCS7Ck0gCQU5t5vJK/fePuBPmxHNJuMhLfiGKqOhmvbWc6w6WtR/WgpN/wsHBNFiWq8ab5
H483rrvsZd6Goo0/fMBVcfAPKZu4JD1v7Br54V3IW5ueYFkTvDV3kFljN1ZckhTTvICmUBhf+8Jt
GHlLwfMVIu76bAs6AseINIcgy6NMN1b4RA9kfUd751smX19c+0frAeNhOZj7dejxWUbbdaQETwdT
+jOhd17wsjdH0kM6s6sOHyvajZprXAzQi6ujTDBEizylz113289EDCcMbCUvibqhNVtdsYNicWTO
qi8Nos40Js0nBLnQznQYK5UJ2oRD6eJiFDzoHukks6eHWtnvTGX/lUTeRK3Dv+8YV4pd+QOu8MHy
zN/ZIrkkVfHA8BUXuyVEcANkqsJrowoWW4b22PNEY+R9WgrwXHWyHLMfw3eaBge8yo6WsP34Lu/R
Hv7MFlntW3g5rTbap+C/FHEII2Wh1pMBhg2nDM1GnKtNIpT1Eq2zxF4qrCwS+gey/huI9nwd97/q
tuAowdZyEQQ8VznfEVy3QtR7MSSKqRCu7FKmYc0YyU/ncbJAfv7cqAZPWZ6jmeHIUZKWoB0b7zy3
qgV9oSrMrREc3gunPncBR60l94R2CWIatj6yFvKP4pjW0rdxCc5j7r8MCDl4vB5buK4sQiXu3715
JjLoH5k8nbAjfhTFDeHB1p0BQEHB8e6Fm2RaEsxE0t4CKLglLpQaTZmQIYu3MTqt6/CfQuTyboex
NgaSyVujlPICOs32OfXZELHcyEBAPI1pykE6lHECG91SArsJGbKrGXd+segBfgmrjSRZ5EWWosjF
PjaHavxyuQa6luC2oQI74x3vW6aJnqtlLkmog24Jru3GaJy61OZ7hqdpI7Gqrlp/nemjDjXaDQo/
Hnh8ewCFY/N8ht8KRhkm60XbjNm0UYzIkcoLh05nj2eno51GYERAeQCFhjlB1VONmXQz8E+i0vjQ
Hcj3MWv5OodKeWByMtEvB9h5WGkvggBAt8zJWVeFwb2bbBPmQGfwgpvrKUNjIM0z7e+l52DMJjX4
OaFgNpkT+SwZfuOucb+Qibd6lXBX9VHmxPLEIdpBl+RDRgkgjFB+EcJLS0oJpZ99KctO34auerjh
5VaCzE07hGO4lIkaESChuyz+nNt5j/fLDj2pBAOy5zzcQmqWuCWxyyyhtRQ2ZD4xEsRU1Lf4QIKm
+I/ABhlz9Dq9c8Tfo+JcmqAoMSjcW9afiWS03wyeBZGB4dNiNtuDB/IEtpzbPaQ5s5RvdedQ1t5O
YOFWrHkRbUhUf5LIb6Jg39JOqCcoJ0NEoXa86bmYtMfYPNWhhjgBhDXjS5g2FFGziu4lyBcyrnRy
vppD4NwBFyyTf8NEiBe+g7y8pNWtTS3i1qS62C57qB+qNkH51M3UB2c9WU5a2h876c4e5KfU+95H
8apQp5QTGuu6fRm/tTebTyXao5OZ/GTTif7DeZ2pxvJM+f44CFiAEL/k3ADhAFiuqbC1iMqwTPe7
+NVseLvmGPfl6Rxc5OUjbHDwxGOtW48U7w6z3Xf6M1MCH+h0Go7AB/0WHH48LP9CVQQycRxa9iFQ
V8ggyhFRUYJqrWhUS+R4HD6jLd3MYuJO/ojnEyOzLfSANwmgmuzulG/p3eRkVLLpCm2eH3no3qh3
J51F/TUTgpeKD9T2XULzBP9HNhcJk43pNszN2TSR3LPFEd8N/ZZ9Zaf1f4xAFbpWPWGG0Ti1LXja
Gx/zWuNMpagB92vooeU4r5khciFxtnqbH05pEHPFmS1HiYjnO/4tX1OmEGQmaA08NmCBQTUfyOFQ
xszAouMLSncpbw0cDEbSyEqxw2fJsk5KvYqW8WqmgXafTjwaF86x6FpwQWJ6WrPzK6/ckAZEx9E4
R+nU7DvLyEEvtnS0fjVUcduBcpeGYq+K1tNE84S4YDiOw9rFQcTo38j0423DDf182CHBZo06GMqN
DyQuGac+Eou8+gcVeL7g4CCaAq0tctdmr3fsJ/CiWQSX7Oup6F06u0GM/tN8l55AxMm7vL0KrUrX
aiQCwlz7QvktsQEuFqcJIh7xFuuh4iNwL6Lj+R6M7G9I5VwFkigjqWgkk0rDoJSaWRH416r6cVvW
+QmwG/3Jz6bBlf+6ZTYI4dmoEWX3HqAS6QDWMqKJ4pV4NYCIXavEohuw2dxsUXN3kRv3n4TR/TgA
o2jI+3R9p/k3ZNnYZou0IVoA9abRFAIus6u3PCNXYE9OJpaz6XZnawOFG9Ood0pVrlQt2hp4vKa6
ATC2YT6i90FPWsN1ebwsJAoSDUO7/jkjcxMpHVv2WhN8eQj+OJXAYYl0aF88Y9xww1Ko31VQzoys
y55VYBBdOAQrH6YRwsn0HxYoPyKTuMAsx6ljZv61BXgGmUYELN1EBr2ZogTTYrbi37OVwRNcz0F3
VZshqQgpHOWP29yDcJJm+Jd+b9iZDRYcdiDF3wqG90or3q2w1MLJUH8rO5AWqQaL0R9QVoiCMgXR
/SawP+5d0VhejILjI514U0w4gVAVge7Uxe+yIifPRc6g6aIPifv6TT2/AvHM2gs3PBMM+h6jX6Ze
cJXrwltlhWU4qGHFvb+cnhiKFZbF1s2ISRt0ggZ79CtSgJG4CcWkkLnUz66GFWhYBjbpAPSULCUA
5svmQmpJB5hk5U4y6kNmWDnQiaXsZfWzpsLB89Wk6MCq8whG2bJzTvs0up23XjZVqByrKfB2r4BV
5wzlP/EJlDgKaS/wYxEUTTGvro/B/dL2LLqMMBRJZ2s93kC++tKtP2Q+p0qScoRa6TQPEyuAhRo0
schkErjFnIXWR1L3Q9SWg9czmLZlKlob1C2GQRJkev6s/dTrwHQ8vhz8YUnsVsQcvvxTZPEyW8c1
n4btKUZBUfSHlnxC0X7q8iUsYEYFFxAfpPZyOrp4enJMFlYXwIe/QjWtGGXuBaZjqqrpuztV8uSL
06KscH+BWLE6orXUGeKCxaoPnkdzdfWOqeyVfzwX5bf44RVTBWkwLVGfSvJKaSSRjtU6qx36f/g1
dLKAcbqiogtS3wLD39eeoslZmhvdl8/4vPmeKwLbZdTTipzKRnrAPgejg2HOmTgngH3/RQOFpfEM
eNqJGCS6X8Jg5/2zVTNSrhjLSuVPbERjEV3X5p2pUKD0FI5ljKC0flXRu/l+xl/cZc/p0lANfCXg
zEJU+oFsvRdVi1A2uGX4F0PPGieyWMWD7sYO/5MOmI9miIu2qeaba1/g9j6gfUVX+58mLfn1Xqke
24bBM+/LAMhwh9akaPAqFgvFAsG1JJPvsIadLQEBhyRtUZecQp9pAOCibkwxijC22VneC2Pm93lZ
YEKbiR3SOYl0aCD5NE42Pa29HCl7CpN3xc/iqe7QQypIyW0GoXsBg+IGef4z0my1EFfBRobWB0GH
PoBALzqPF6k32wk2YbmYpDIa9U5UZUDMHDvtkTqgINSc52Rg6GirW9+9ehei2IXj4Ue3TtMAsLDl
0nysLJ2ONp1Wq3V4VTGAVpDj3M0Q/gegsSw43Xgvb88i5UnmSYYYs+vmTPh4doK9aHzdS+ou6ob+
JVd6HPp4/9WW8P7bDN2cVRIKV3zE84opvUdLfWjgsV0Seuykdhi3GnjZWvK8zdHO93Ka5TeV0mTA
NUvKqqnuMZhe87oMW0LtXp+kgAsgObE2zGVYY5Fz8F6LljUTsWUChkKAE3CW20KpjgkJm1HBwmxp
swn7S74LfEHzXEGmXXM6SpQ6ASwgyc0cuKygrMM0ovmeTc0tnTDLsUzLK/5aeD9uqILS8uL+R2zX
4HeUhgERtH6i6/fHeByT5cTcZqXVbR8zZoNfO2zfDFsgbtZaGWcMODg4X0lX46gtu1Og2NqiBZKe
48QoFHuDefoMKcH3+ZDssEjdLIzvohGEga7o/SHMRbASBSjll5SoO/04ragTe0ABVvSGak+U5Atn
q20a4Z6zli9zI4i0zev1mOWJFSsvXPJiKdRnCS1lqzmNNYCsv3gSq02UIXbnHlfFAsm3QmcILoRf
QBd39QNAXZM4YATiqWibQwJTMPkSpHrOF91oheqhaHSk8PUhZq4M86ZQlOh4wHhIMnZWA+E1P6JS
OB1b9A0nMnAIeYjwEwhfRrLHDmiRqr/ceTj252wL0lfGGHDYA7lpjyTikW9q7CTs/E8d9xvKiZj3
YhWERMzmcuzDlLxVQM8vJQzkko6ZyvYx0H+OXmmu8QnRq7Ebkx4EqreqmoTMfSSiJZ05FAy2P1+B
0yUv13/DLwZP0/8cCKX8zZ6yIRejAGTjOFClkCbdjGNRW/tZcpZ2QrAW1naWSoGHGwRhVXMXnfLY
JAph4jqGqpyZI8GvyhWmeWwHoRJZNRZZRLlQMiGQ/lu0GC7qIKffmP6ye6e4C3j+Q4VEEmd4P3j0
2+CSRDYZ2Pt7fJWBQGfIJmuCMZoh8v2RJQs28nSskGc76lY9+vkG4Wqcy8Qu07GgMscia2iNfSzS
2CKrIWxSK3lqjYB6z+oarcx685Qqfox/KuZTEppN2a5wVEG5cGSz1L0cYSzK7Famu2T1yAhzl2cr
fgV6XJuFl6bOhCC0971v6Z4V8XZGaxskRVw2XfNaYvUnQ7CxUiq4Gw3wQH1VDtxcFBf2HZ8d8+3/
dvw5MLDF1G7Iouee74LAukyzMfewBm5e9JdNuunShtmmdgoHMcoPgnSzvpIgxKneV2JNHiBqJdzc
rZeGR9Cin57vvTJIRry1o6PkO8zC6gX5iWU3lpoztsqsnFEZv9mu/bflYe0lEKAp8cgBfGbz6Bbs
icStk6xXoTOmNTgbt0dfPTOjNMTULYQc5uA6XQIAHr0cwPXu9N7pFftfKuBvZDVnmJBGW3wpC4X/
Kea03G4P+1f5njjHJ9kQW6iki5GbXUzth15+adYzx3tmgiAszfSkMR4Ruzq2LfZ5AFWj3TNTTQ2U
mQOjWxo+hb0CFgfUqdVRHtIfzGj3Al5GSQcVR6ln33aJCQZwMPNtoSRSNQ930es3Mf2hRBMC3GyC
JHtM7Ud9C8PwJ82QM9MDR1Y4F9ujogvaVYeQybzAFCk736H7ItmSTwKrZZ1nsNrAY7u6hKJapzfr
hjUpduL/C5YjEW173+iNp7NBMYBxlSOmx74okoFiqMSgVBJDNftlUkggH+wLx4wfN/L1lDwnScCq
z8JJDbkRT6iZiskZetHsBCzaDT0nEnONK2gjM5mHd3z+RbSl69ea2gROKCjy60R/P/w7XYTjrzWA
RyQj+qn9QcvHrbq3kQ0RGjaQanV3Fy9Gy+wbQJmJ4CibYERMORu17mjqeYl0ZMXIHSMrFrG0Pnz0
V06WHKOMGSZ34r4LJfeL9a32gMseRPcqu8f0Dw1oJ/zXkspsGC9aHijnG+Q+4kPdAtd7xFqHLfje
PJu3Tnj2yZEGXUGRiLqvE4GUdIz3xh+k2+13ukQivQHGd/1+Ms8UuRnBLLxp4aeE66AxB7YrI5t4
fZyFn/5KT8v5vo4yisxpycqHi5DCQnkYnne5RDsaKwDP6szG25wRfvS487aQuwGEy4w7Q+u+96UO
fQ36iGNn0/vRGNUWnm9qwsZBcn5yltAm5VVjjuL7aUerz0bd5AdhF1s+f+M4rb/kfM72r6tA1h5M
GYRWVERhEvBeumsOr8yD9QJSVHbrzngsUMudAMHlUmI95na3FHdKS7YcJkvrR3RdM9N+TAEsTN7i
/UkXqdR4Ga+w6HouGkneP24j+95owc/rrrZDu4YwKTA974d3rLwVrFTZSTX3EHfdwF/XIbb6Wg2Y
NtOsQ+VvC2aAP6J6pFNDlsuwdMj9mGpK0vZ41/dNnWv5wlVtLn1rLGlnKCOTo942CY5oYxulpnVJ
W+7Wn6jchNy/EN6MAn7DurrqnhYIkA9rm1+e4FFqPCGCFcQLe+wIZGZIIoqO5RT3xim0NCEzY1Zv
RXpHqr0gCVvaDBTnPwAwi8yTm2g7IMoHKOVIG65m7uIF9p0etWyKWcC06iLdyHeQd+P/fIOaeNU1
Q9BJUWz7uikZpBJ2oyRoo9a0CYSFsQi+RD19YPX//H9MtE3QoEgzCtbxgmldrgFzKbDjTLQDfdMd
Rxuv/AH1PKPcpyhsOJL2YtggOB0U4R0wgsP+S7wguBl8Aam0S2FFChPTrIOodiAmwz4ZZXEviutI
X73d424S57J8v9eaz43slOFJLRXEAw3Hv/SRwDUCt3jHxUy69kv8AZeVrtwI4nbjqGqOlZiT3Ap6
+wOK3iWXRajB/q8iGii/lqEndGl+kF4frLcInnekOPCkhRR7TrmiUSx2egnKT0eL7kIkw4mDMcp4
clS3JoQvC7Tu7p9GMadqy/kZDdyzHFqi/wjIc5RSm5/Tl58vdQeG3NCUovKAaqWAafELxx0HAuBo
IpSUYS3qR3vkQuUeWQQMhvNJkXM5pYPIdp1Hg5G31Lt3kSDC1raqIIiqEKL5mTvbq5/zPrwsrUv4
7C8BkmFzGEZHsfy37CowvGQiIGWbDIjNqxIHolTz9Ckp2UtGwyripm0SgwUEii47GPcFfI+k7/Oj
jsbVQF00z/IAbbno5IndPs0QtaIu9iKQygzs/jHlsIFEC1YQgXL+nTA/NKf/b1kTAu0CqHgbji15
LvFxdsaRrSZFKumSFSgoiXUSrUc3+N5MbIhOSPkQAIH3mC23ILaks0i4SbetQ/GHeDUvqHFrWY4d
9xjp+qvYGBJiRuDjgmSFbWUfT23H+JBtrxzeRtbL8vWPQADai3ha/9f6kuPqCw3SNG+qOHwAxGti
5/Uo47majVZVv4mV3/GgBCwjm59UA9hlh1OziyccYDfVs1UfkBHS3z7JXkbOnmgeN3k7K5qGvL87
1fA34x3HDTfoXPKwpgE69up6IN51fUqfqPgblQRPBQY134bkPylJQi5etDRhKz4GLrHodT8rDi2Z
WcCND+p1xy74E8Ewvnr3o7ednlLEYCbeAGWpQmYn+dL2s2bH2tvQ2y5kEPwDivE7gTgU7QNJeQUx
3fBP1XJhMPxe20xxSY/5ZqgqMdjVCXdRJ3J5S4xSPJ6zB4i6Wljq4J/2lRbEFmWQY02hvKzzxYiG
If2j3hz5Fez2yeeEVTNm8tgfmJzex+Nl8cIQzUVlLBvTzIqWUTIdjeG/dIZFKJBYjIAKL1L48i6C
LpxhBPVSB03W4wyZejVUJStuaYCUtxcuOpgqmXXVUNIaWHaGNo2i2ALqLWlNC0ha0ILhAetXPUDu
hyucat3fYpaUx0gitm0G4Hv8D/X8z84IrBQYTc8og/TEoGAH+4rDaFR76vylFRNKZLd3GuR6Bxpu
uw5U86JoDLrusK1QIM/9NKuoy2JThoeBFW1Jq+6kxBMAFH2ndE3rDbrRViSqQ1IePrRSWXJp+5Ya
mhDGj/bF7Gty2kpFaXLJm93jVFTdR8iOjuKDNsuWYOD1KyxU/CxMz9+Jx1h1cpuQ3PXiARq6/Iji
yyK+Nax7bEhdQl5yipqIgAcFRMJIl1sYnac0C7iDukFHkoGOahmwqn7pIqaiP7et7OBcBKHqxX79
RrgtWBvl3XwlHoM3PUdGUCpN6eS0N81KWOtAai5UkOygafGEwomvdS7dZNzDpdfA+wezQbydUUx+
Pcu/jqopRaKG5MLyaJQpeThl+lPBDP7D/RCfsMIjUzUsDf1R9VLshJdsTuB+t8ok/sMUZYWzbQ8p
PxlvikkUVO3jptzgOYxlrk2SlTHTzSwHXnKCY35wCnF4vS0YVUJ3Ql53NuYQaoPZuzvMpQZLM/2U
XCBo1VYzUePZEFbAL1NMej9D7ajOGFffMbkswQUKHlmFyRJ6FD5iECUcdg5m2rWyyKgpJgTjPK6n
HiLdlnBHFhMBk4g4UiGkxOT2kLDlrqlIaG5/Z5rLnq2uRrc/I1+8hE++BidPfYTiTWIQcu0/2jc5
1/HkLMkE5/15BqyHdHbpVqcGK/t1KKVFvgsNJUWf5pqhnWgYjQStiD9rHIHH7aRu68Dgzmu9Dlvy
d4hTzwe36eS+IqIzqgeMpzXEbxtJ0/g4VtvW687PyED2tpxYUm26LbsMeUKs8xbEj9MMmKXvamwo
wDEsnE3TnMcdm4a7HhpHJpBBg6AsSQXRRhSooxkyTpDC9fyw3PbobXpyhh31AmSFeEAAUqCVTNN6
PxzeLoV6qWt3hD8q7/7DaBAA4KTb+BHNjB2VLM0Zr89mhOEBgyxkPK1Pea7GzrU097OoDSoS94+x
++nZL04EA9agUttFrs7z9t2EojxTgSSWAVcz1y6u4QN0RRudfL10+tuNgGCDxjoiSlwogrOpW+75
vIg/hhp0SOk33hNe0VpIoL8t3bObpR+jdgSE5ZkVB7tSQhome8lGkkJ9T8ncf1KxdzlF/URu+0lr
48ewcWE6FGyExWyqyzq4yCdGOYCxkjiNtU1Rl38Jln9S9Y9EhLF+qddl7Xm5bAZkJOC2dG4zsowI
PYOwr/jzrUaUJPHtDc5c8GHM+ofF05vAEeZ4S2zxGD234RuBLxMlT3T5FFGsVQdkqqZjHz32JeO8
N3lcvcsJH1lI+VbkrrWUgHcHTydR0JyhicQpEYMxa1wpJkDtpIG3HMSUePpPi/+slcFykhx/x/rW
eQ5ExQcKieekL8nbtdF1rCz5HXTtigj1LJ3++jYE3EsVvnuZOTyfq5bsxsSuSByKEQateZDhYA2l
mpimQ8drEr2E4FHadGQp/3+T8Evnz2+hUx0jOI85yhiL5Uo0JLS84qCcntqW+UHQGebNN1XKLwx2
y3jC2sB9KMjVgRpINATm/IrPyF+g4yAZrMiCYHVc0TLwknmKY1v4G0odOfagcKEYnzF4EOmrbJO9
0jPTX3LjOe8sJnQ3i42zotbygqJfSJLbY9T0oAtkeovDp+qhHqbv7GsDQWsrXYV6LpGHZB0W9NIX
0eseSdENsqg+JbSburkvSBqMr4kbWu7i9mD27ejcGWa+jSVDwO9GZULBh7suz1OSb+WY2w3QYJF4
8nNYS6J2F4axtAqkzAxM1m8Z7lMf1vMNf4JXi2fdRbJ0awyNsEnxRF+cOAIQfNxuDDg8aFiO8m6j
hD4qtsYpUfQ4SQxLHoNXBIY3m/wg9ybiw590UCu40he/7V414aLHucjKoe8jQ6BEZngrA3iHETdj
GacmPS5DuLhT/sb5LIaBpAUT6Uweg22UXskx3AhaO6lt3Fvo9Hl8R0+LZC0hshKGBxi3GgmCangm
nacZI50ERuytK/eBVacE3LaatuiUF4P/M+UgNXTaiOjlnOkAq0B9AAjhxytkIF/JMtBRD0Z16jqr
l2GYve5aXAbOKr7/GpXBS1vhXeVZ5nUJpmJ8wEVqjPO2oRfyVwTltdICUP9VOxZXVxqVS8KchuO3
VyDAysQ/IMyahf5nA5s9mIJXe/t7r9tUTBvhtRszLQrBs8hGbKH4OM8P0kTaWKtmSWplHTxOns4H
UB+SrnbVlq5mG1tJfd7DVItlTipteyVKaSLiqxeCBcpBHC4RXM73TR1oiv0UVBSAT3/5d6ZlWw/b
uOCOqMDqR/ioreiAn48HeoTyLIL1KNZWKiwNMQooyI7050CtnQswblnwDgEZuOnNki0Ush7gOK3X
yW6F+qv+2OyjDAze3N8+TB/IlDgaLCKoKaEenLTK4ZeBBu7jEJ5RO6NAvnQPEYfREMJML0zFm158
dd/Hmzju9aIwShkCE2hAy/L7rgE2p6n/2czGrylvfSOZYfztJ+/Tf5S8ez6VdbRl9Cpfc1vERdH/
2om2XTP0qD07hNejSZyLfI7tRb9B06czIVxBMb6iVDuD56ACm9QSU/g1ofEz3h6zrdTOTOTpCjqF
YdOnJy8DzDiH7TNIyfNfxVliYGW47Rt+qgH5nFf9R6PjcVqNE0oHo/MYcGyuJUy+2Ms1F1xYZNCt
qe2zrzbHH9eeqLPe/jR6FqLRUWXtj/iz8j/ecWETyTyVh7a6JB/e9CoDXzGikMyKewUslqfY3lHY
Ps61GFb/bIEm1AlES5IcnmVzX1IddMwZV/sKW4iCfrAvrCzryhbObWr9xU5XJ49LepRv6bw3g6p7
cPfoIQDjt4chJVihzvEFYIrmtZk4dCIbXKPolRNGGN9kJ1i2SUhx+XvbD3gA9Tc+Xi/6I08pQWti
Bi38yCVPMYr9aIA6kvejitk1DRgxfn7H7OAQYW0F6/MihmmPmVgsYaHk8bGLpmBCSIngSfeGXi7j
ARjyCA0RDAeYBDRo9MADRi6XP8gsgQYtiGd17acQnGJAkAqBaVWdY5DjU6tMnRnQyexxIfCX455m
PAxSVfJeyiwmPX+O1H3mWIyOIqzXQqmSV2t7aUm34Ss6/sWn7xaGSmEsh/cly8LFYZm6jkeuCP+n
tfADcM6+Jyhv/wJmE6CQbN0nZ6z5Hh3RkOGS8fn4uQHbioyyVYBuXlN1+GR6ZTW9lbge4kVGZwUQ
NuGUCnF5j0dcFXErvBa5V+6cZU3kJ+mYofA1BLl+6Yi0IVKewZPOv61JsSjCJ8i/K48l8xoN6szx
HnZyIMPzvWMw8A6eaCe+QGBjvXo0ZDFSGeXM61ztOxIszaIQM+C65D73j6oVC7RJS1AfyC1DY3J3
5KSjXiH245NBLatkFyFkluZUCbbl40iu+5u2OgglwG4N1eWAacIMpXYXn6GuBWPDx584H772xO8C
Ifo0R1g8YwJRDmeop/SW7P/bVYzNRfbJUS4bTO/4O0O7mizgYxmdlbgZyFIRw7c2JU6pAzdwgvTg
nD8jJWFCUIWYg7/rF+rfbaXvpQM+2L52SJohvbO8DuZmaveykM1t+oEwe9IZ7bw9n87kGYqU2nVQ
iQu8S3wjeoB3nmTWYo2dET2b9zOE3e6HhYLSMLgSH336aaBTpzD2+JbZMbfHlp9lTwXoQqOmgNnJ
irKoX9238tILbtWx/NEEL1Fj0WxLmSG+1UPham5N8D3anw0TpvM+Olxah9TFSLg94ajPS2gwP0E9
8YCTEX/Fqxsbm4PNzLkepZAUODAVm+mLZXjvYNyjptiPuc5HkMJkYUb9kOvJNGQCVFYaUlLBxN3H
uqNvW/8xyPJRSy53svwQgvSNf4Rc2VQaWf26TjcuOh+wNdadJbK6sCfYUwpbGOfkldQ0bPEZCZD9
jGNqxnGjSNo4QNYVoikrwn73GC1287Whw+WXEdiRIe95YTZFO2SmcecKRAzGtC1ThhBfvouohh17
pfMKJzFoZfc8mdhUHx1h666WTNLUnu/p+G7DFbqjP8EfO4CRi63LPSNefVMrzxby7evEG5DztIjm
TsSo0RPaNv2vvc21i8mukN5kh0dKtxFhsBQKZkyNhzG0en1XXJB7IvNa5J0/DDL2Q1JKfp3mwd8N
58jQgnsdTTFXFp1zSrPBA35H11tVfXC6wiD3GqsuCKz6+yJiVOiWVhiqRDFY2kfzNQDFMD1SMh3Y
HIkrPUxQ1kwtwGbKkAT9rRkwNBOz162mHK1xUL7uJ7FvTTHGuUSu7h2aQypZaHrfWm6VqM+YXbfZ
20G5ahbHzT6brUa5kFL2LINHkrdHeYeUvH07NSIZO4H/Xe+Kdhl5lAu4/ePyj+h5MM+O44ohlJiH
4WWOxWDKurJhLJ5UmVg+uzIkJsGE9XNfftRnQtn6+b5B1zB48DmCI+iM9TgZhFRX6RK9ijAMKVxX
DJT63X8vjuSxXq2tXR14EcjaWA7xG96PKoiIViF6TXpRSoEp2OMdv3elHxt9+ZhPpqIOEDt/kgDq
7qSQnlcmn1GR9TiV2eiUsF9gXTghq2ta5v4WhD70es8q6NP52DPKjU3kX0KUFSvyhLISBJ5R87UB
ft+JMncdQdWMU3LRAXITFRh3wsLfJ9ceju+RRZvyF6zDeyo0tGBG2wUVzlD5m7bDqxmND0JM9osK
LL9J+C3Tlqm3Kj6a1UzUlpd7QPN6tdt6pDs2m59ZhVQ1pZ+rvrcZiAGLRYjCuQO7UR+lnzAxuat9
BSDqNXyr4hhwWXJmeqK90FsKh4D4f4z3ARvtWXSdQn85t4AOwNPv1WWES8LH5+81GyC4cY+cOzXl
FKGhnSOTIT1oREOq3kVNmCCOTx14D24B2EFfZrZRGnSil+HqYFO+1UKM6hke2ZbJmrYZ9fUkf7iv
d+DParHbMK6mr4ppreM/TDWiTo2Br1gfVpBvClDzwwb/Gsh2wTQoK6fjt+GHDnMOI2jQ7ANFKTok
SiO9F1VhfXzIhaM7DS7KXf7qH1oMFPM9cDq2c+SWmTY1VKBkOZ/tSowNyXXskR2GL89N+9k9hWVR
qPbDFCn3QtS7d+VkYiM+TmoLv1HO9Z/lZvkQMmAn30onJ4UC+MIwVJ34IlLc3nDoNPY/PLr5RWQS
ilNTN3DrkfhlgQgGQ73hXxEsER/uPpYRxh3Cw+vFeF269Z9YcqpsVwUO9rXl6Ihs9XUybGi+dysd
Ez8JFWPpQ74WbzuzNrPn6I5hv8WOerq8vN0INaxf4QXTxkdIopytj8FnX73UJjwQ1ltvQTbZjXzI
1oXXh4cx1RnxV5cItOXvd1rIQUqGpTbQ4oenR1yfm75LZ1XFf3XQDCPXSuANqcVIVh7xKpOhUK7k
hUV3DgZkrL6icOc7dyoenl3t6EXJVmdVVQVwXiiZ7JchVooWJU6YzLW9ayjPK+bI9APmpw/VO6ZY
nH/9ychf//g9KEmsvVY34wApwLwomaD4HAHW+/8FBX5IySlLrxnuhGCb1hEZZaSk7dHy67Y2Uoe6
dAU2ty0oFTjyTS8D2+IiE6P8tkI89SrGUV/2gt2jfm6gwEbSdJ0Y7ivsstEpe2CA/nn8S1FsAjM2
Aq/I0+I5Ns+FRiCQucZRNZx8IfwAXAZZUPAaoti5cyTIjfDqCu7166d1V1UuqLOwGtitO2hqq3CD
YXxSrL30VNNDX7PPNYxGohyxadqw4jxLMRvAJijMyRRje5gtZKa4k0Kqw+3GF35kDBk2BwTFWYrq
I1Zk2KEusZYl/o29kOaCOhfuUVGTeqzG4iFgJbdMdl8bpUVEaP6JD3GtSKenrH0MirIEW3X4t2O+
nYSGIsS4S02FSiwLmBOO/9TZHXhibKOqh+FnmDMFnpaKRR9LVIpPqlmiyL091f4YeYnohLhoPSLB
KXxQQNBLoZ0Yc8DoSfsOBAkU8bO9CJGjxY9GtY8ZE7FgLlXXmR6ec2qKVIP6ukF6krzd9VRkPxCU
nnjybW7PZp+gXnB33kjztYvWKrw9l2ZC1Rke+skQBR3962mXckCKl0woCkjUX2oZJ2+/9C1EHYmr
i20QVZ3msQ31+lq+c9qhkOtmJ3ssC2/06kGo1MOqJ8ktJa0J80JnQyR8qfXOcrlTiq+v6A0oS9iW
NeOm0qJD31zzTJzZUmi8b+bEqUOpeYBQ3tCkvQ/TFdhuS8O1Xvgvd9kLcm0UjSz2OmmBn8a56NMr
ukQGzT6VZrx2X1oHos4I+tej5bBugAbKudxNduWIzPGN6UWFPYZlwt9xtNEbMCIEtE+gfIc3xsOe
4TEqgLGoqIyCeXL7EcfqnCzDuX1UbTTzUXRf1u3ya5j+/VsQw2YPxwOSwWONeEA/NiJPkG2voZkY
0Kxr1+DnfMwXuutIIkyGiwGd+4q9ep1c9+bECJi7f7SWJ68WmH5CSKZRtlY8piyIwFDCQLBHeRaj
DPciUUdVWuxrII/LuRomCeYLsy/BjYKyCoR0qhoK6h8XsKQQ3jrbUyeSwNx8D+tLNKsL2DpnOlh8
tB/HBm2UszCirbmfxNO14QAeaKOPmrX6sXqrjL6hvwUUP/1p/ml43D3j50M4JNH9eYBzgwoYBnD+
fS8seRh10aLc2/+lY5SnoM4nzwQl872txP3GPjpa6YwvlnO8xJOiQGkp3whv67HPdmY17YlZkGbj
87zbBfCKy0OYg3urXnipCM/fZPa+MKROswdtbcr/HXT4DHt/tcrfWgztUYEZCgSOsrgTcXcEEg9v
zT9ld6fCPPBeHHDBf+ojDWnkf5Nyk/eBdXIo5sBnWy/hKvjH5pK3snhhGt77OmqMisZJDvRL1BvT
QkTV/w8qQmtpiIHamm/cpaHg9kOaGZ5K4oJpwfKzIMHADcCcS6CVBwZI1WvK27ngefQOAF+Le9x6
SRl/9uH+aTlA7HmQKoT5LrZH+NMbu2Fg7n/KFUCTTwiD2hYeZFzBJDlor4Fr3WYQN3KVdqerrfiz
HmAtWam9YcmJI+7Y82XEyAQkC+eJ+ROAImWwRGnC0TmgfTXv0z7n9xwcnNtXuimucDCHFrlmCZhY
ts+46tmoMogor7d7qJNFpnTm07u3kZkmZRnCeKfOM9mGLTn06/28X1UsjEq9WCNvKYYH2yIfv3w5
FoWrTLphT60ekuARngELZssetkvag4M6qSOPVlcI6Mas53EKMXZ4GVxzy/k+u7AlRjdTn/9Q5BBi
UpHZXEco7qhAitHG03QehZ1XecLdEYB1ZFJcKOpR0q8QyVyXUXi6nMQhQwzMxj1GJ4AIfh0yG2hR
jWg794JR9s1z1QUC24npOazPwKZ9sXijO8kVNYynmWBVJYA2/45xIIYH79BjOtwhb2dqKDifgXFv
rgpHWzGCy2LUrdp/wBWlc4VVRJKQe+wyUpSz+3MHG06vkpuIxHypdg1T1R88RDJIVJ0NVJAwGKpB
uruvOQHV1TOstQCfF9OTdQGeHjvdr4Z/U3edRMsJKHynEHwqqrjRv3K1hH6mo+0jOX5bx875QTWT
2cApDG5xlCJ6D944atdA3+58zgDwliwMp+K+S/JMej6DEg1RmgrWwOMxkUPwe5Q8C009PrN4AVKY
C/r7KkswFU1GmbLeQgfTP/H+ZJmetzilhe4Ve2JA0l10AffyEs0D/uTY3eS/Uyojt83Mx35Hrjsj
zGAnynoFZTxa6F6BxlkwH538laYB5NHtTJYb2VbZZnrD+KxlvLXQy/LHJPG8ylGW4bwULwzvAz1V
mU8asYJ8+/wiMETrumElTk6dzC24uy+gzs1VVrJ8n+Hmy4aZq3lrUgtcCGJn7kI7FeJLx7+etMPx
EctjJj6kOWmTuGmk2soG1DPSwFeQf0eLkOwBShFcyaC8GAwlFHhLniA/ainhoJeuDB1CU+lsemDj
D2cBiIYAyC899bM0z10XzUSrcihnhgR57lNP+KO3FQU3hPOA1Vd3mAJ4d6IJD7dOJQ2fnvFvplVt
goThHyUirgJ43qb2G5AV547E0wRrdkb6l0M59VfH17VefcR5peCoiqJLIm+4Cp8YQ/XdgOoEW7Tx
oRk7Fo/q2jn0N5Mci4IilUDlnYTw5FfvFLmjkfwsIAfvSFRJTFi1lOjpMZCvtYOzMIowwYj5MUvT
E9fPmi8OE24IwSdXFrCYKrwx3MFK4Q+OckkXabhb7fV0XDmLmo3lN3RfK5tzW+WDIeCg631Dzvi1
TnABUVWR7iHfTsPCsRthCgdj6Xkvi5aZ/8VDBwYOYw9F6nYrl6dDMApc77n4oaNcs6tnAwDjZ42l
iti38C8/a1ECuRc4CXfY49CjVG+syME5KHNu+bZFSBAdiEzPAK703THkIK+T8iFqwEy9GYKn+SMw
DpiwNuvjype4EQj6cE8azA/K/AdaDe6pV+bjfR8AOLEDNQZj2XOrHMWjq3SHAGCLtdVcmqvDTlPb
MTLXnWqyMxheb25O0haBSUwjJU0M6NNjUZmCzqxsRHfXBLUfR/bfsNV99SBTgYCCpTTV/o8yTESm
PVAXUw2ymPpyCY2LDaX1Jwuecdpp0b0Q4Yu0r1STFPk+VKwZPdTfyG6FBXH+STQnhKNd81jyO83C
xE9JxPZbd7pVwBE2sLHiFd3VPiSFc68e+q2MJhdDrTSMAao/Gq6OIrELg9y9xWpNhN6sdKBCO5Bv
GVGml7sVJc7Qp/NO0Oi8k9Qn6D+BJnIeitLnvjVEavmKT9IINPkYpUCuUzQ9wytXX8pVb5dQhuQ/
rJ1iLOBNMrdUMrfY1oAjhjnVRCfgEZHaF3MFeP0nShym6/zn80rnD8BaJdPuUmfjolroZotZsPiv
65/eYSi6cQN5W2Ne+8yBFDrNswlKRF3N2VVqWqdd754XoeQ1OLtIZ0yBKjgr7p1zI3vyUV/LEmdL
tQXdxdjaEsGKym/3HECFpOUCZpoFnHh0rLjOiyOe1mLV7Zx/qL2DTXrMcmRuSm9vdU9TUESX3pjD
L+dtIMTsZTARcnEapDbRo3fnF/07rYXB4qOSqjRfRTuJN4BU9kdjsNJyFfzIiT36y0KftIXqxXMU
iOJ/qhXfn67xElWYeIcmh69F+TY9F5bkHbme2RSrPSpoSwbcbwnHycPVUEDhvDbEWXNBh+pBN5lf
GsQ1s9rd194uSDYDQvrC3P3OkFpGWukG/lUduonyW/McwlKhQIwE1DG8I2WKLOKDl0898rq9CKv0
kDlV6AxS/1Qn36w8hy5OjMX/wRDa2jKF6xyfeKFWaxp6u/0SGvF1TRAKJnGw5xQ2ntUXAXxJceLL
si3y7+4N+bx54XHF8FXyiywaXQjvrnHEbQEE45FuQ5A+kUicEDFvZuI3iLXZVSdvIqQvphgU5ua0
Sl3B0SP9uagnEfB/AZxBWOGI7Gh0asf4tWKpyZ57C53gTLYhx+HLRStZHoBd2D2ih4g4wXR2hywG
SnnpTKnHIE0K1OGvAbaVl29J0uIv77d6XJComHsD28/taq+0vnq89cEv1Hre7f6rRkLu10J0aRSS
dWOPXMLHF6U1XxawnW/PXFkoPsP1lMtO+IL8uasvShK3BlHsEI14BX9JiDCYaPPpaxo/+R9NceDh
XLR5irvvDvpAYTzu+w/hsl9QkH1W/cRea1+hXogIz2dv3GcyO8t9j0LwWKU2BRVEvLDMWQMDw0Pm
RsVweWPC/RF+djJ9Kb+6R16AOcw13W9jrSCCDxtpBnKcoWTgTaF9sR4qOBOSwLz2/EURdG7xG1qL
CYRBZ1g5Wp0sFWM0juUHozUagkYO/yttO2qN53kw6NvHz3LxX8Ast/heE2hG5iCRMc+28My4GJtq
xgyWWDG7r9E85HGURvCQcbOehls/emEgpVZ8heVML5oRqrUPKqlxTdirg9QaCEvGBRjFtKkJVvhe
Wa1kIEjrLBaceAUJU/MhPSFTExHnJjH4mq4ZwkfX7nnz8J8Znbon+V3Zkr5ciukrp8d064G+yS/U
m7Xh2bKIv3eHk63XE/Zo/3X/BEGxv8YOKydRYBJYgEbUuYzsOSJQ3bhcEi4wdQhboWKtXwCMTPGx
uvuNXnLghxb6536vjnc+VOPq/tNvocA8GoU3n41TRcGrTAol29E6qbJqQ9rV5I58rx8QM0SrMk2W
wnYPKyDaKp6a7iMNNYB9jPkMzrTy6LcJeP27Dhih/hiS0JdQft+6ytBrWSeR/p2NnGMgHhP7f8Zh
pf0F0/moY0gY/zfQlv10m4Cf+KsOaF1dWHdqswX5bPh8ZLq8xnFJYilv2GMTOd89/iuDPWRqTG6M
K5+NilcGZApcY+64ljwUxxKpJzYAN8A61CC6+j+Ehm5w8aXdb4p3VpZhxFM+d4U3Qfs7udQSPm+b
pj8ldADmWie3I66O3EgiPMJTFk/y7TxNkD1DvHbdRCWdh//tiF4X2j1/4h1tNfxrvFHBzlNbR6cE
sbT7o5H3HSKr/rz4LBKx0B+G/XL+3Tha8ZDMLO5PCXEjYRq4WAVY7RdeqaxbqO6Q5q8AwTT7Mh2k
N3N/ayv8cwL/cWW3hY+yyrrFq1sJVqPSSX9QOmcHwEayUgtjXM4hv/sJf4eCZHQ84a+fByVfvBRT
XYkn1XqFmHgRii8gbgjEmSEhC022QcA0HZeUeU/ovJyegk16aYXdc2Vl+5oWS591o2IkWejULu41
ft2gWioaSfCgVuJRKFAgJBzfDdZCW+VP325iwF96+UWoIljL60fj8mFCR26ZJnBo4shl0xeA9vq/
L8kUCbrMpQ5Sn4JG/239q45wzU/e+5nvJkEMjnX0snA0DGg2PkS0p/rruLY1CWvBO09vW6C4CL1H
Kut1UZLq1xMJiDkpqkksg+5TNpSUKftdbdTe7/No/cIhv40vgl3hmBq8IqQ3Vj2zN046MkgYpGfY
plB7aTlXpxOMZlR2JudObwVH8a7glmXmUwv7rr7/lXwFZVtKGuhrGkln5xpSUhiSl/jD+yIxR/LX
a/MqZ2g3AyVR36aXO1xDU1H8nHerz5zYYeTtd3JQminQOcGQ4IWJIIzUTydZYe+wunjHsQ8vhU1C
EGikZ4AONzzwHofTF4jrEN/owkTPksrnq7H9vl6s6XNxXzw1w3Uv1bcbi7zG/cl10XI5c1RizmNW
eXzYbdDLtBsdn1xOorOrdNAHa7wAMaaJcIV4mIkqFkP7Ug1RMwx7oioXiY5VgUOceiYbWUsIbaQu
jOFmLDcTnkJeBBQ+AhybrhXeZ6S18xuwsclE8oMm6V6BeAcy9USERJn1p5w9JEjxpi0yqDS1p/vL
GVfHTrAf+QfaWne5uX4LE+U6RcU9aXE03GEahza4qz0lSFZMimgkJi5B7RKVwdEMTc+j+JdtQ6Il
JBlMieKvAEWxMN0mphLMz8jpfygqva6t9mJuCVAiWTc5SLsf/AZqxI+IZN0W7pjFmHcQrF6KzqS4
PrUQQNJoNvB45hsFOFnb3D1EddsVmbxOHQ6nsMdivRAjmHI86WZlZIA3vqZ/FHMwPfmlG7nvUGT6
1Mwq5G9RiCiZBnHrd31nSncrzN4oeGeQMOH13XqVMdeIBIbcAhR5TAxWB1k17yeAJ2AB7diaknLv
eZ6+UzS5EdcJpJRwkqT6abGN4gEPUaDijyBBhgxKt+zC0c6+/DR2rF8QmD8IVfGn7WJwuovMQX5l
DnLzml266fo+MecQy86arvizCrdDR1KY0FJiufGKCLRv8eYm2yTy1pIG3cAe0HTBTdKDAtNtyQIS
5pR5JG8VddtcuKrtPb5SZQZrwJ7Vhzwun7Mxdxmv6xuE2HJD/eWcRc9+8I5310jCZFEeXNi117Nh
JUMMjUTj0qSv7jkf8Emznc+Jc0Yxnzw4drkjkF3yNfXy2/RbbZ82G+OindS8kUkgcczDS9LxXQt6
gKfy69EFhaudcAE7LK1XCJdI/KNQoYUBIlrsKuD0xMKe85I7hmdytPltAd5U6U2mzKAtMUlb7Co7
82EPAGcrqfWjHIkeX4TCjlHLw/F2v+p3seL0DyRT3mHvvLX7vqwJLTC+1X1L246HuovLt7sLJgYC
bj7G4JKG9ftA54i4EjWEGTvHloHjxVJttjn1d8LGF/46cPyNj7iCQ24V2E42vx9U/oyHFFGklilR
GOM5s8aOdIR6fGWObVNbIHAsfTjqGXtWiCQlH3I+WMWEAnYdIlq6jlsPDmcZKS+fdMLCRo3M72NC
OQBrUgnQXmDkHL1KA0/966SXrsyofQRopxwTY/nBQKNg/qTb75Z7zg8Qpy1/hjzoYsv3jBymxOvQ
NeUfR+3mi7zUMbQ9GmrlD8q+e/mtshoewyepFupgEwPJ7n8ETIZxj3+yIYPHG8TguhiRSle0h72c
EQWaM/wtLJYUfQLkJ0Qm3b9ms2QRm8FNBQPxCWJ1Kb6YJfkvxUwHb0YaIIdk7fkio+K5fIbRn1a8
LMuOHaQOYj76ZTG0b1D570bYAp4MKlleqdR6vFgjW1nx4OS4RdbCGkT20o+/JqSyExNOUOB20Egz
JWR0HLKQjfVFKTBqsuToJ7hIjZ70v1cFfi74hs/Da7a/CXgFYNn4a833Tch9EHOVpC0XUi26tCuk
8/7dICXYohltHnDIWO67DlTvg9DuEzVviPw+X8LE9hp/jF9QZ54Be8pI0fKnfPGDNuW1A1JRLIsb
B1001T2xAw2HRDBuX7trfXJoIhI01pfLUfK9U86472XYrYntEq333Q7kjEEJyJ9d8bxzyAzV58ub
nnMbkr66dGaOfRS/r+YraDC7MsR3nhzpU6djtLF9ZigMYSVCxinibsdD2VkYmSq7amCtNJf990go
7yB5fYUVU1sY0E5qLBAuF0zRYvly8ITrzZ40tyBpukBPHt53QzZcs+X6yslGkgohpsUBaDHVkR97
vYzlZAqQy7ygHknRWSi6a+KAMbsA4tHYVEgJE5mEwTbMGjDryuLrB0Z7e3h8f+/XIHmlgKOOvEh2
//fzYnxVbKFQp6t5uOFpLwvnXxktiKer2ruDOZob03vCFodEarERMKbwah+vrXoTqDMljILiPRyY
Nw/hi8sqKiD9w9fXxS7FZ9IwcqkievGRns6L5SsRkV8QRMdWYPtqKZvUJHnz5+jYsF3dpK7xhZtv
mM4tpfTJ4nnWwgts7yWH7EVRy1V3ZvceMTDAf2qKAvuqT6DCtP6YnpMGQzSWLuwF+tYwOSPHl4n1
dtNcsPz/FN9taraoeIIflZWMCIc3qIEm9by1VVMya0h6t/RoiU5pGwLQcGEL77ZAgaDPNi+pAgHL
P4kL2SdXOA/tZqtLkqkHKj9ysC4W0UX4m+/HoXOG7w7Oc3QuLSC9t0MvuGKvDJjuv+2OI92vNTSI
1rgym8sEcaPmBRfV0j+8JRBlfvbx0/4EpUBjFETQb04fqIV6/MqiJ9hu3Y/rFY3PzFpMmfMpxnC7
vZDe+6UQMTUThQYX+xSp8Dabg6rG7vYoMBQKPDKbmtu0PIaina2kWhP8q9l7diGWIHOV6+7b4gnJ
5bUhdecRCyIDyD9uxtS2A/9uXuxSfjrYAxLXpk3EYOhDPgoVi1x1UUnNsbxQ3xuQ5JJQSTkJe34U
qDuvcsNEZHOJ63YSBEq78cZ0ir+r727ny4bfU8AU1y0Lktdn0hEirOiiCwCimw09jPpbl7yZjJvo
eOPkgvdg4ICALDppbKXZnO8z9B8v3/NSYQpU+x5Zk/R9hnMmswevXvoYkZ4QoSEAb8qxx+lRxD6q
J3FoHRkHLtrTY65r3Z7VL/XdKdVEJoJ7zrKkYYlV37Fv6mkg55l0krpqgVa06AaVH8/enrFtji0p
1elW+33+FzWtczthe+mS8a8NtzRU8Rb0828zKEvxS/poqgA1NjFuBiiymoSFbP27GrKWS10sxGYy
gsxl8JrztorH+7fHhMsmc1VKjuEqjJ4vtV0TuifnYX7rogI9qm6jsmmc6TXy+vU620A7a0AvFYKq
SKFhIqn35eqA5yGAWCSW3D4evibCzaVlscTeRPBscyeMCeMc+h5WEslZ1CYTO6IJ552GAksJ4G41
bHs2R5ROFhmJxFbWhRXxwVvSCc+yYtAu51Vh3PpQow6TokmHFCMbdf6sfLwcfeBKkhqdmEcHcdh+
qMYeqcU6VgMEavqzFDCDgO+FzG6j0R71JlkU7Ccow6mNAdgGbF/uvEO/RYx7AymPYXHAWE3RCv4H
mfxhX1LPaU7Qt697AOui942f5QteVUbs26RDw5CvQTXHm3zgA6tFT8PypQ+lboEDKIqtPfeWloS9
uokK5IkzGkQsnJ5wyTXK+CfMF2UnnpEY1A9cPfLyLVheW8WtEdSqjPCIrpxWCK530nI7UO6clPBn
fZJY8pynG9P3SIVxjTLnIkCetcbA5BDsB4a4kkR0qIMEVHIol7odEMNkKTg0AfFBGzhwXlGctikA
45F2kSWbxYCwe9haqv37zTDwi8f/YYD46ljUD2ccENwJ7BjPUENWmEe4PyNOBc1GJLEHF62DXnok
c69r+6RloZQqtFl2UPzDpqcFvPn9S4VkgSWncct1z7tzmGK+SEyKpqFPcc5T6vlNnq3gpawsWvw5
Incxavey6UEgyvGm48pJ4SY7lp+wqUfTAzBcyeDA3vA/OR1ZlKBxNDe8WEyEk5GiPlPYDUot7Mex
AowSxdfRLocXa16971+wYPsfQdtAmXNEcYsIZKrafA9DKWzNTlQ2jg+LbMhXc9dZBersGlPNMsXL
FlRputQH38/zWbZuHLTtyAjgfY2y7V+O+UQUWXTVB77e/ekZrLZ5/nTJ6LTsJ5vQoUWICoUmE97h
4/mjrCK8yPSvyu+Y1ySmEqdT4Kpg+Oi5qo4wL4oc3iFVzkn6n8HPyH6MV5S71j3EA1p0VMDFr9Wd
lVo/P7ALF15BK+4XAqke37b5wKG8/ZOyyP5/nBevuVZvSJMsr1dF7IxzH3Zi31HLHMmAVY33Ez7X
iWWv0zYkvkvAeia6lL3oRIH8uIqU/MZ4YTuloW9NS/QjvZDR4aYtU7cKzBljInZVOd504M6f73Mb
HS9v27LYnI9hPuqJA/UVYqnbJa5YVViNRIinfXzmq+wjuM4DUzY2Pa28SJPOxF71+okzT8OvoDfv
Qu1jFerO1+hs3G+7pWSHmrywFuo5UrTB2p1eY34Mn7ZU6lPjTRpLVmEkSIMbP5xv6pKyVaGJN5/l
64a3IjGwvFU+9ZZFpiwgPQZuaGxUfJQc3dIy4dIJj8CWdsPYvIKxOpE2ZKMpxvVER26RrLICXJrN
Er9NK9IGMWCXSU21k+gGcn8gknE4acZidE5gMuWMdeh4cIAI1Atv74zAc+MUjCObp6gwzy+DZp98
RXZF7fMwmSIQEon/dm7pAbnI2DFDORN+BOKq/9221fuMQOQ8L6TZCI0PiXUR6S0ynO5ur52OTljz
5D68IrqR5NR+fvdlT87i7N7ZX2hWqUL/zGdQVNRnxk5xnjzgqq8fjn9jXZkoDlwPFJyHc4sDRe+5
Wx+NhanrPG9UBsjTqujvnrHvuYU4Rq6ghzT0yjE04rdu1cMsuhowiC/xCjpZm1O4pihKN6+f6Trs
RMZvTe+Q5uvEacSF8jQCZHbpXJ82G3wIUDvvw2P3NZ48jpfxXb0TyUyZv+26GPxDtlhWU/1YndGv
uiNsWkey97jAMMPly8eNLsT/oFvvVWhd12mFMrh4tNnB+sKseyyIwJuae8IVJ7itH+EKxPtUou8j
cNoL/N2gGInwO6SZNCbcIsLQyRS+xSxwmVIqfr+pHY+M2uuwrobo5x0V5TrkMYvq8ktRxXIbnd0l
2qE4RX8oF23CJCbBQL36j8cfVIvdQWEj7Yisvk3jsGNVCwyfERqrsP2jX2qBtuC89bDEw4MvKsZO
NymRXA31vIXe0hU/rvaR6vqfwN6VAwCvu8+70d+SJ2X6/+6DLcBXWsFYhR9ysy0yDUFl7x9yp3pp
D4Mxjc3EEMIQ0RmDkJx2h54gx3vJ2XYkUTwMjOcKlnFkg1pqrR9Ii8+azKbCp8kKzKguc48pALY/
2FII2rx0PY0YGEPazhmwfb1lXNfGWaNAIxpa76uTkVIugLTqkzJBouKVnQW2aYcikJp/5sfCizcu
fH7DkuiH6XltyHsUfMSABFrV6VT9gY4FYW1dqK5P1ySUlrR+8dgDjDl0budxKivvm+m90HJnUKBM
miFYVxoAXBjEvwhpcKXZeiEh4QCfBpQDZHy5kaOjk1Zm7zhf0DN+4z1C8gKwieHZkZUNgJ6NPrCV
YecqM48+9cDmA5ZE3KfqBOF3TYfop+A1i7rvp3TmiXSiYhGcboaCGEKxI4tPbnMfAisJGbqUzFpR
BnPK7vUJgHAh6jyWC4vwmZ7ZICArQOQbbhKo+AULQQCzLNXmfNoD6ILOrM10/N1Bz14aXYh5+jFt
MkqhDNG7bDuoX1EYVC72yo6ioINw+NccW/UeSnQbZRpHbEfdYxjufxpwE6t9Ccdq6phYJ2/lg0gz
9B+uwa28y6wRhzTNfhP+uluwBnK6LIEsUvJte28JbGj2S4zYWjf6a6qfTHvFAcV0c0DbhPuAVQib
xg/+2sgZwrXbIz0ZpUnemxBSU5R92Ucu6QN93VdVL+dMYAk21b1lIyigm6V8rjToNF8932KQIu2i
s1wnAcwbhFtKTBSbVRkCTeDKzOR8HdBLT07Eg6Oj27uTx464naexwX88Af9l+HJ8ro9ba/WjDMaS
NRdWN2a2FqYtCzP3tkNmpz1EWR1ELHhlJw2yHbZZ/RXazxZLjNDcJ+5AHV4AqyIs7HC3KS/pnKO7
/qciBGzRhoUxDEunlUfxsK7ZG7r/Eg0VZGdTygfnmp9oXOcRzXFjgXZzJa7cE8sx/jvy7U4qFMvS
rVjIYUoh0G78Ng+ntL5wzfTNYM5PrMsquqvXiKI5ScduWC13PtNXOgp5LTSFeoNX3ot2vgdq2V6g
h+ytwN8M5rlobMPrF5V+NK7MW10fFy7/AaNA8UbAJ3e3bWJWmyTmj9/YefzdKYzP7uBg3ClQvTpL
3oDRXJAho9iTz6srAdZaln7abrypAUcYGKCr5hfkgucvXp75FP0Mw/WjiK7Ow6kw8EQYfY50Nbyy
aozZSaXWkCd3rJrNVZf4rNjKMcyDMGsEhgz0r/s9MmEFXHnKIQvRoeQ3DrIbPvEig46hcglmEElm
yWc26Dsl1pcEcVybRfkbM3NGRqCjeXE0eA6r1Wxodei+Mb+QNyYhawUGgdbCWp4eVDRSRs1ZHQ5E
uhRBjrqR7y2uhghT2JSoToe3SjdjVcSFF1Gu5g8ogdcMdA/euR35Zdfy9CheWFQEhSW7iSf1fBZn
p1CE7XWaU9Z5nPUNYS0UuuJWBS1rU8wV0FgM9w35XLLDxYQantXUwgJU4OKTw5O4uKIFj+iDKqNE
a8n+Cyl0bpxM/JriqBFNZ0IUXWUM0dEXjxQH0jwhkO0fac5xhsrLxlC5SPnthVR+ZWdwhOo7y3J9
5EM7TgDbPX1MftUVEx//vuJFzbP6hgjAYkljKS4nU+Zs1W6+89ere+Njh2EkQmF6JhbG0q0jJU2e
eN1Pm9eJiduoRJ2OUyVB4rnlIeCAbvsg7RRXM9WldI2+9Fl8L2+J3EXwaqwdsKU4KnlLM8BjIEAq
+f2W7+PBlirioM4SYT1v8cIl96FTVccJFbQzv1u5q5Gqk4TzTXsbTBpUr2ba8DdqLILASKozVTZx
gOWhElNSEOPbeJCnoBqvsyEqExsTXtwuFv0wDxEaJ331hjIgUgnZ+a5mxZnmCFC9Usdp+CGGoGwF
pn+PmM7WJtgcqx8At/weVGZEY8j9PUYs4Dkj9T93geTRLnPqgi1+SUpKtRCw0xMNEp3+wuMdJIzo
Go3EzntbbP5IfU+Vu1SNHBoPq+eENP7klECFIHGNl2N6dKnVfZRHIJLi+r+xBSBNCiLoTGSpm0Kz
0NryK5Sm8nrlTPS8xk8fwESGcIDQcVZLljgsGLE8ctsRq2bQfNy7X3rBajsJmEOzeUIludwtZ1Av
iIax2fZOWd/AR1Ox8xAcXywJjPOEL+pnClQSqViitXLfQmglbEuAfEzRBgo1l/l+B26dIfR3QfX9
VIwQ7Gtd4ATNoGiicFQMmVVUO0vYGlIAx2+Y1WGx5HMa/BEyvgRH81JOx/SLt47337JAYlmLz6uK
74kJBNmBuTtbFIpDfJCfNttJoFoj81WtkNx5krMDrkqrLYq09Xby918cWUat/1jyeeIaXWXF9fcP
YOTFRZwUQ6T44OdmZe3NSNsWwONemvACgkK0LLuAXfggXC2ABTIsUGQ+cqD/XP1VZsBww5yCtm95
JAQDHRMIFaIZ4C3aExHszpUCHIlc80G8ekOp1AsW8z7Br3lwCn85A/ZT1929fX73ZSpSRYoMWLuZ
rMV/2KCgim/4ITzszNldFebVY8kCH8a04qUT0jzlJD3T1dU6Zyc9sBYG+UdkbokJ81hBgtinllH0
vX161sU2la5yGg/5SpKSZAmvDy70Jc6Me3HOe7JUgCBwx/olu5JQkBbxEEJrfrHeliCl49xHVe1D
5Bhof1wfFKXCgCxpkJxDqgD4bLWYsVOJh+7AO71eoE1+KbaXM52g81YKAudQHzliSx9c6s8zG/BO
CktwZjPxp88u7hUKdj42QQxLVaXcajzKK/oBDR3pEEDe9ppWDIeKlbEsmsPaMiWEjwt1WYrMirAX
T4WB5uiLB4bkzMp4ZCTamgKH3KPj/3rxxZj+jgwYbfvYXi8rdE4qne4rrJWIuwVny1KuXuaV/n12
RZqXYIRWTO7BTVy0PvoMNkeOA/8YCPe31g+iJFUij8i/JWbJJPxp2QgnVtS5ucVpezU7PRVAU7v6
k/ir1s5+apSUhukW4FmJmJkY0DUWNjIGhGxiRNshBPeDn+/w+n/C8CH9urIAHjqiLNoWKQGu7E7q
Magc7wtCvzX6/AYUg/ALMo+kjlnleMBwLw7oKlFuTwrBI+nsNE7tgrL0Kzy9fLh7GgqO9VzROM46
5hvG2IZTDmNCjnw0y7epnEE/YLAkZOjpgTqV8cWc+FL3sMIdtqGAAsgfztFa1L12i24IcAoae7AY
L5CMJvEotviLCFR/uPuHlYZrm/DOsNsMmORIBKRjayokIMh42wDyy+duNaghwh+AnXxWNYpIHzbJ
b/k9va2R0FhhQzd7lHzgHlCpPMXGXgL/nxU9iu9C11ejvAaenfvgigldYNFr5nr0tN+Biy4d0Sv2
t4LXfLYJ9Jgq+oOGaP7HjckQDYWGDoXYyuMHO/hjKtwV9ZC7ykNI9hETGmY9qa2dqJiBE0y7XV0x
j4w3KOd1ZNoTRai8r6S/e45fC/7pE+MH8QvHjNBwFNlU7mSv687zdCKFQ139uvDH4Ogm+olFgYAZ
rnToqwxrBjYWkvY9Cr3OjCp+InitHLT/JyCdB1MrZcYbqegeIxyKSt6rsg9j22LnC7Ht0r9YmG2e
5Em9ITP0OwSeVhrUJN2ZZTPr679wMrbn2sAIdWzHzcBZtrC6CYJt7TYv7oknc7RteKoJxzwB4WGL
4aKtv9KiWUom21+GIkbL0hEYS+i8iLxbM/CrrSa6M1vuCf4DSOq1F7O2a93CObdxXBhkqdVYSQnN
3gOK/QeSOWjmlpe86wcHpS/RpGGYu2QdbMYzvCH1LxHlE4ptrQWbiQ44NcXcfOr+G1Bdm76mbQ+2
YSwnen30N+LDpUkeh6Thu/F93tFZhh2nauszbi8cuTos9IHGHPGjblpP9V5/T/3Uzz6eYOGyHjl/
H1OCeWu4CWZ/mHHJ2/xa9a+J0KIV9KB/6vrzXBDo8LykJedO1keq70yb2gsEQBs+erAqOE66PJYY
v5tPANBr/+/0lqvcFzUsyMGcTAIBpGpuGaJhZ2brOz4flJGw2ieQGcf+9gSzF6qfg3M6J5A9Q2Lb
SmpC1q7fGCPZxBGPlJ6wjNEQu4Svp6YhUfUlHLEVnMepa/cLqh/D2M6eLIIjGdJspworQ4DcFY+A
jM3fJOJHi8hmnH/mmdy90vTechS1tXRIeimWn6W3FFzyJThEUBoprNMwCKpBUGR18w3BGt6xhu9L
97ZGSg8p1OCvOSK/+23ybNgQgDJadmmt+bLh14ysXS0zzeD/tzpH4iv1NE9t/J9u/2gwYgCHPerN
VzemL40za2NxVsf/pXiuJ9iMiGA+bdCDWgycssqtY8+dMeoK5diykMvrCKtNemTSL3WlxnnsNXph
U2TNAXAd5lCueRM8LSdifIc+gt3Y4h0FhQ6W/oFwAmysDA41CvKiQXiIVNzvmEXGs2Fa3436va2j
yiPBAh93+jxBYZ3j4CNyeukXSwjZTYUb6jGTgDOaHCV4lPtXIQGKw1EutJdMRzLAVM2hEer6au0D
fWVY3tqo5wafO1cTujcvug/foLDCEOqTr21vrNjYV/bAJEqWj5fvl8+b7a3sapXM6vFwNNDlJqye
gZ7NAUI92jiSEtEwyB2Sox5bbVDJcXEzode/hse5ZUsoE4/uWOhMvsk18zrtkbNUM5yeRsPt90zZ
7TIfPiXPzx5CvEkJvxTfPS0vPZbOHmlm2vM/kPd7dUzrzinHiOkbifFhqNVJzDVF9FDve1A+V7Uj
l/3lAwqi/CTWUqhO8PLWTnBeF1XDrncBRIHEfJYSKyyvnGcgqRiD2Qg/c960dyvPeUmJAN19fRKh
iT5i9NDpM6mAz9+U5MxMorHRUQVBtB0rdRe2GSyC/qZOyn1rAHorwpusnqqLqO1P6SUtMvSHKide
qjWaPQfTthsQ9+tbjNAoUTQ8eadNLl8NavAXK3s/XafxrhnokiwMzugbGNzr5HiFAAIr3wGx+2Hf
igjThm2WB9LLa150n7CbGuIxYHO7j57heujyW7iOEm7LpAmrMc8w/0qSauLCa7VVfHqptgA6GtEk
/yGet5Khe9XOguJEoSK1PrSQpEAOxYMQ9imPjwg7LRiXjWY//qIdJvmHoOfs9vVlNWISuSywTE4H
Uhraya2ZvfoiRZCLmGpMAjv4AHWvHdUZPz7HKuv7TwIbPqNzk/g7E1eSmTByh4yC0+vuepRgzBXP
0suhmzqHSg5JGe1p0IPXa77oSZ01TAaZzG1rm+rSo/ILqlzlmmY6XDPkYXi4TqB0UkunGwGo9Xb5
2F0+zqiT/RwV/7XkHjX+2alrYRLMEc7EchPdjLOvwrUyujlz7EmHdrCdHN/LtgTE/tk9T4gJ2f4D
66nNfO8gatmQKILyZHPuXvoZDUAao8wau1xMjyIvmD3D0fNq3YsCMutNPawP//iMnPbKSp7wvy7B
DXG+P7qozI//wzQabwRmyD3cMmX+koMnohv0wqqgFY35Ltt49UcTcWH4fV/3YouxRS6xplN5fNqS
RhgXPcjhBwMQgulhMQGdRzLWpdmO0AE+QMBoyM/gI62eKOLycpU+D4bX6mf78vzvlaVEvtiVJyHg
L/nEMUccQcrGKs+DwX3BPu32kV8fpGQKwMRx7RhaxG9Z7mL/V8dG8NEBRA1Mt0WYJ0PZSX0eKBJR
ihg2ryrUEemiJ2JPFcYNG4apWLOtwHNziQrUlX3K/ZVy9DPjxlRABmV4x0aeCEed+oIupcWtPfmc
/TPv0sQ5tF0Lh32VnS1XjSj7vkEwvtgpBYIs5PR85vH10GjJNG485zayQmmXFkPdLxRypoz8Edx5
Wc6meYupHXnTtBEfHNANdaRhwLSsTUc+ypyWvUjzYu4Obns/YIixS4Buq9504SpAJT4K1VgoJwVQ
aqmxySNCwWLZZv6IAQEh4HVynhH93PLQDHlknZeTKTgkgzi/3EkuVcu+i7Fi5HbuQ/2Br5752J4h
8mkRYKhdIbHymLIov5tPCV/jPFPsxXbFlTfj5M5rnlX/ukT77wDTP9avyTXolGoQkSyO0CbxvrJU
QTwdrhz5eDtPxAgIkB5pZv+3cteaX8ifMOJESuRnCe3WMzeBtc4cP4wX8dCp3D3ztdL69kp9AXt+
TXh8iHXtva23PMHxCDmTG5bh4frE6tqXG8MjxHZVjrp3RzD4fwdcf8OTy7H9BXiEn+fKQ+xdE45m
SWVkAFGTfWmvPfnVAE/7jgdnRq5DOs3deeKIBlRjz4861KGlftxWk5WIbAdAoJ1vtF2w9JjUV6qm
R8/yNF+eJX/e6gW/NnxrmpMiEa+lvHkijiqh4Gx5qt28G7TzhkjlgZlQQnhK23gHNfU8AMh/ut9g
YLBUOUv/CZUsTpXJ4OIDZQ2G4Wa55vMQjOFkmj9PGo3TaohDjlFf+d9imCVcBgi/vveayBiCyxlO
0Ub0fPGgeSS9nL24Zf9G96/V/HdAZE2izz1vnVSpATiX3WkfSUl7lOzzJK81oYFyF6hSRZYF9u5Z
JmoKewY0IlhCcCwwEG0ke8dhAYJ3iHqAzYzbVyjIgv0/hyVGJknMbHF3vJ2J3trwslvCeYB7aiO1
tIZxgFlBckFtuTYjiuloff0J2nPO8FSH9hUo+nAJ9t4At4GG1fyVetk3jcgik7u2jZ6sRGJloUzU
GNPQ/5VRDKUlxSV7CDiiKzuzSX/VV1J5rzzEBuaKRAwaZBm++edgYJmNUo+2SaObwmngUoMqmKzP
WZZpFNdyoJN852Xhl+qNqtW5+S7csMPlz8uQYZvSQyAmUs+rlo0iFWammw53x7to41n5vbA4AqkG
LSM2kxbrEeYgoWz+JVl+aya/I722WAznhcm9DWcjMhfX1Klu/GBZzd0S8FK+A7+6Ee4Skmcm2lmd
b5sLxycUsgnF9Nz2TeWNwrjwc7QSKN/8tfXGzZMAwzfJ+nwYNLfIiPIyTrcyWvGNastUU8xAbbOu
8xOYeojmuobr0cKx9llxpEYLHxpr8IWByrKWJmkCyp59AFXAl9mkpVTQTAif6GNtgjVNH9KW111I
jxc05cUH5Hn/zYiPEhaf+qIzRkoxPFTmHAedKYVnmH4TT67m/an1Gpm3/Y9JCQul9s0tAgQ3O2F+
tBpz0gdttkjUy6X+QqT+vPwbX3hlbiWp9phj8qTLOjga3ZGq9oAaFF48L85pC8RTHuywvS5BPthH
CaVn42fmdJeHf89uR4IWfMalC3/tAD4W+JMcufLH4dBMHp3iR+00DfEBhT13Mva4EnDA0N9IOA4Q
dbXo5y8aa1Z87yK/383Jaj+4JUpxyppxdfbT0eGV1F10o2bP3XOXbHXeQCwjN2VvryOVhu+Teon/
3E7vntDRM6lBnUeQ3cjKJ2Rx1sMlTDL7Dkj+5KeI1N+buLhdMg/chBiUZ6qf9X9eeTXO5sAygtsl
bm43R/20bvVThl928wHRrHklXltss+tjNrz+20FUeRzXXWJ9Nd5qzc6imORFJLc2+tSG5bdBO3Gd
TgjK2vce7nEUPpiYmoxEV5V3V9MzKKfoW9mp3PieTtZRvnvej3WxdMnyw12ypD95VU2kMKEXFOWH
PwurBdUMLTDKsZNTGAs6hfqHZSy2bxr5Xr3uQH+Onpu0ZXnkufls7yYPU8S6qw7wSFkYAXNUrOL/
2wXW5NjOG3bFOpVWA+qDbxX+hKkM0uygZd1CfB2wW5kzIiS1vdxJR/XvIKXsOLIALJ72e/TqbihX
QcHFRwbnR5RCiWKFZYx+qrktTRzgTVttokONbD5vUDMpIRniMQ+KGVX1jeqk9Y7TCpBsZDqtWKY2
2OibpYDHWLnUP3vnbOLMwSjDSXLEnzhX7onkkalS5WfTBl1KT2X9EvJA88gYZIkYHZl9oNQnWnlG
ehAbugQpPBWsFoGtKAa5Jlyx87sLS9TLjY7a35UbCrNYTYNpDjzuEW/rb26GnF9ABLCbdSoLPoud
S26alp9br0h1pPuwogYn02Sr7Y2HpHi/ccmo/t9S3RFsjp1D5mlNEJKayevawPYuY1OVKkCSZoX7
Pe/np9FVRU8leD79ghIm2h/myElhQkoRDgC+64ioym5KxqMsoHUqHMcjJRveQxCBltBcUx3/4rXp
6hXRyZ6SUetSGNX4b2dpUwoYdZzs+6ZZhhmem7AgJ/wxz5RvH54bsGjxC3feVI5Ngy0y41OQR1ff
3nXibfQzUYyF3ihTGFzRIPafWhbYmnxjbIDZwBzRbdoPoU/HxF+Jq+8K3z6FrZj74jnGyovoOrSj
1WFReTot7BuY3d/bTVD8kvPVmVgd5QwnKwKLHYjn67xkJ82mFYrF6QvTMvixNB+Y1Atl45LnFVKt
kTaU6C7edyzpnvifVOHvZt/P7EprXi+TQHGoIWYXlM5jkNCsB0+o3tfhPEHW6lt0Mw9fb3+px0Cy
qC3gLjnQX0pdysmxSrcw2qDEW/h6rqN2e1VoyXpKgz7yH2l5+eeD07itAqT01Xrz/0fLWjR8cYl/
A297lkb2bvlA+UW77sUL+iFcc6VxzpbYZ8rB6xf2h7BVeLK1/eJsRQdVjUWBK3FccDcuWimYzmtW
J/AgussU3DyPqnFDredPWbpL/Fl/ggyOu8Ppdc/riFCzA4Fx0qlikFo28iBS4FvuXeYCFvfEQqD3
OysR1A9v+g9eW8KFCDy2yoN3tsbukB8pmP9ECYcB0+lF0bAmyvpWAU0iTMUBw6xrJPCs58/w475V
lvVQTaYt5C+f8zpKmv7QbqSe/W7yLpM4T21xla5P2cz6sGwkHeLBn6/Jst9auYOli3RQ6fFnCucp
1jLLTQ2HHXmpT/oBFRULMvZn7lUGe4oHYkOzj20i+93HtPLUdTAVW/wJ2mjA3TNeXMW6prQby8BN
cPxYE45CFYVtHZhxDLbemDAWZdBRfeJ7QEzYA9zFVXq0C+ewtGVXxvZkVEX1TO2RrxCXRZpqDQxX
b7594ViJ/3vaTZdQXuHllzN0sY78ODxeUwYYeK0S+1HQpKbBVzG2e6DH1/niwz+Kmy9gX/2aoHru
prOYRGR23x+QHp/3ECgY2iJ/iTKxWGN/5BpD3mlArWwrS8sdDe9F+DIvekmkDR02+kc1gUUiTMvC
XcHqiVDc+IeYhzIZ+FOh0P9yRsHaGFjaJGJ/w7URaRWV0dk59zxkCQl7OYHQZInfAfljDvdhf4Zx
E8xjh5SvRezDpCm/23SEwYNhivBgxYYJDNTBDu6QSHPR3L+sldWq9r5XDt8RIra2LRoufP8re3hm
Q3IVEHo0pZ9i9mL8gsyoiu8vL4vOJqBLRFO5XgYmKj+jGCpo6l4BRty0wh3P+JNKuFDXMiuDpnWX
7OXOQYdP+ZzvuUnpCqkhutpFQRssjVfBs/NmNhRbUUWeFX5HrihASvyCETucAalymMbO0sFOX11B
zSI/a1F0J2Bw9f03CpyxpZxFLh+0spPx28Wa/Y2BQuNuCCO2AcAgZR0XhH+45UxKq4374/vkJfpV
LfnrNCfr2nY1LdjAlHlGG6qoMx/vu0DYFJ1xke9GJePbtpRZFb2nSD5REWg2dYzOB7DjyfHVAAdq
R3AWukLoOUF8vvbFKmva6ivPzrYuFbqDNKlQrCRXgmN0M3xt+zGWeHJYERScxsjgVgXWZQA7QuY9
Wf3Uh6KjwfvUuhV/n058sSa8oOF9ZoezlL4+9PqG5GXojsB50vcEc83fldlMnobCteoOPXoBFxv7
kW3zXzp67JdE7LGrS+45Lqh0OUPh2L1tcV7pLTrlaPGJp0yHjWCqpSWViPOLLy0Wy6uHgJrNWF+y
q8nfOlD2mM1oGjMaMaAwXFDe/RAqCqYdwPC3vQazDxDouHevsKeyJoFOG0WdTXWwJiIHGMzsSfCT
xt4EVHspMg2y+B/hFb6O8fkibuvMnJeGz0r5fRhJon7VZA0AAcDiWqfNjQHyDzFonWZ7oDM4Gxpc
/FAZVANFYNV3LqaviFXcv8mJ2JaNytW0IDVwZozv2VKzFKLH5gXOkN6eg0xKcU/hXEmYUgEkvkBT
xU5JekW52avwrikAnRi7pXYDJ+x0nT5Z7R+EYqokBSmNhjDYOO9htNK90cKBZhiuuljjo6KkVLtR
IHIlNah5lMVGM6ddt3S2fbh+yfWm9j3O/vG+M4Hk1oWjMbzEzcp3H9kQ6qPAGzJIMBiaS31c6eed
FsF9yUiDClLxFtZ6cKIZRYhS/Tve5Ft/Yc1jTXkDfjmfSBo1t62bX5CuztCO54BSxALmzBhxmi8s
wti++duSKUzdUVaeVXc+107hAlnZRUPmADnPXQ6HLmCDimRav09fniCpdQQrm6uo8IBr6Jc63ejy
vbuZzYxubCKj5Or0qng4WApdgZrrGKqkiT8wYQfHyj55GFjpB7IztIxE+At/JhRji7BAI0wEB/ZF
gRsgSkIe2x2fw+z8EyzNeXXKJkV4Llx/P8TCiAZs64gSKNDeluBC3dq+8DFOrbYrIsd/FVkbQS4x
19yZ6OvrgeMZUcCwpcsVsrnSW/RM5+MuRyzgjJzr4tGf+GwCHxpMqn2EMdezbNZc/RiWzRAag+Im
iU93RgkiSfI/AynmUNS5SFrz8gpieCdP2GeLNabNtovbUtckkGzv4l/LPoiooP8yFQZOvO0ZHtWg
ZlJ9n3GhiBN6+3M2gpesuBPu4nLrB3gGu3Cp2XUwB8h0ZCFo9nZr28MK80u/qFuKH/GAVVQmG1dG
lzjd6LqxWh+lSdhdEd1Q6JNsIWEwxU9tf9UW8BoKXM4pzbKHMPfTElVL1wUxAqBryW5x/QJArSAq
PJb63uGWUyy5rSvpoCuUufzUsGAAQ+xeiQPGuDjRYBarzrEnvDXxaHqPRo+1iNt2enl42N1sG6zZ
vJF/V7Lmajm2EuoCidyErmwfoAa2xr4SV70Bz2T2e1fX+VJG5lcZQMKQUVOBhmEt4lojaZ4zjXYf
NQwzYCRbhu+NF5e6GVuMyUNxAThwLErjuwlMpplmW1Ch80qo/skTv8OfX3Bx+AEwseRLwzdrnt29
4f+fpBbtk4w2MzhlsFfrfU6HuNHQPf2fDfMKnRfuLUlUK3zrZGp+qsrUwUjYQ9XEO23otIQXBZsr
eOQeeu4mQDRaQn0v7BI5xKjprTKk8SVpD/jJx3wAm5CoyEAegMtLg9ejF29XRQobfX5IAkgIgAPx
IsKcQQLeDBooUCDqR7mN4y1elUdSZgBFeO33JDEIjC23PljFauJ++wqRfx+gGWv5962ag6N8g+cJ
E4NARct4WWZxNioDWJ6W0E6Iqbwp/a7Fl5HoNjUOiPwjdL+I3LqteayK7XC/guGTFYRaAOZYX/Ov
g9b0mUURI0vaooVNXlz+dNSVpX7VtkjM3Ove+1J74JYmuR8M+W1y0WHT55GaYgbFJMXDnxBzrbJC
7OC8+QEotS0XDdfRA/HNTI8R+Z3tYbZTF1i+vG7Ant5kSBWTxSHWjn0eiJe/R1hRKkinz5Hozwvg
qbUMCU9G3FcAf1hV1C5aGgW4WADqp9mGZGNXsicFz5OiH86onKjFkPg2VZPrDLqJdHOlb+iDO78e
uOPvSQegX+WS7Rg6HlxQPg9mvDYbsi8hsgH4nOOPK8S4WkTn7usC8bVPvzHclprct8EMPnlHcdaM
5N1ohVGotDzfNDq0A3040IOA5iusE2sdn7mU2ugA8hIF6alNHUzWqMkafNefdg2LGoAuTMS3iUdz
Yk3iSyEL1rPRzG4jN2lh6hl8FhgvKvytEuvAtw8iEGMGYaIHGja/T79+tPszfJfbYxZHIJK2I76y
PctakTlVGBmrHOy4PjzLkyskMzo2LwAv+4Q9dflMQeRR2vhDGFko/v77OJzgtQ85sDjnk/NL2K5n
5uvb9uglvJaUnA0+mC4k3pRSWvhb8AjSg/BUex/lbJGDajw8e4tzWUrFOS88xJlrxMWXO0Su5LuK
+06eU6qsXUVirM+ZTNNBygicWTtM7zJtTPpCoU72PY4Zhqkkqq3V+k5xnJcY5UL0/9CtKS8HGW7Z
nzGgShEcb+ztm6CIPeljO+kVYwZLGzhTOtn/P9G4laivyEhHmb7TneMSQEgiRXLhOzvOcUfM0f4y
pY8IuW8gGJptLQMmOJv1GNVdM7VliEliPd2uCP7ReP9YxP9kVdPHIeeWyjQ+nfjovTAY4LB2nHrW
fIYi6PCCTYjXWMjIxMlHVteWtH+Jpltu83kkMggyQdYo1xQFTmd0Wj+DnK336laz0wkXnAMi9FWq
gsVIvVVCJjiRwAn6FKFGC09p0+IgFYBBExq6tX9pnOKzUk7lVeLiFC5Djc5Ry+8izw9t4ZIeFyWu
jl0u4LZyDbyeYasi0cwLNak0d1PPkbQoK2qYvqIb3JDJc/GfQP0CiIfUsLmKCmNEK9ZV4Bk1NWrL
3/Hoh+YBsgiW3+Shq1yPGYhJuMpqEdv2iDO34RGQgWUD9YP4BE/A2G2dzsMqLHMXUmm1ZGKZK2R1
XpVEgonvCXyHulVBSBAhKTeLbtmrkW/p2q8jakLYzCeFW16OFM3uJFFKogjnPUGh67a4KqENCUEL
B3M8B0d53ouIKNupxc3RM7vCJhklYZ5sTHWLC19dshWfZ7Hyvh1dsdZj9d+Netwj9qTsomF7x6hF
RjFns+pzRW6ka6G+NDGEqb8WAhBZaJQgHiI2oscM2d6j36QFfD6xopFkRo3JTHykd1kSkVJPtg9B
jJuv3xbbbdeg0PJfnB+nI3cVHwl0an6W3REM5K1sGK8HPlT4IRJHrLUKZGUKoRidUFytbW01Jgqr
EpaEnb7jIUwNHd//a+Ug8Fjb57eV2zhq52K+qbNkLjAVy7rEE87aPm7GhgLhZot8qsqaWuoXNnAp
3a8kIn2VbPOhNnmXPwA4OBjUTWLvJnEuDDu8EiHY7h5pXj2EUl4uyC9+r5liZIosq2z48jqbBSNO
nhX4RTU+8MfVj1yEnZfKDbdZxiWC3+SO1vDupErOpkCtIBrAv/EtnqGpoOwB1UhEHk78si6JbhSr
aj85bQfVW31+3bPkt9yciqpyt8HTzj2WIy5LfH4taSsR4CYSojwZYJZkBQTMPW515UrI/9/KhO1G
yglXdQhSNXQcTqQMTedaRtyTH703Fq0ncorP51tfmK6ZiZeiaeJpoT+ok+aIiEAY5+LWhaUqTcx+
1+DMWXNTI06QeejN0MHEIMsWVuj4o0sqlMFjR4pCP6P7ZmfZ3YGRNDHVsbKYvK5REhwVn4oGWpdv
Nlvgrb6QXvTHCi2R4Kpon4uqwKu3IKe6ksp7anSdUlFFrDhF6zhOIMjM01FMKGeHungsnjHIRVgy
ti8VTL3Jto2HiFdW46BUrpN13sl6dJFN6OU6hcKzjgwv6ddEFNUegv5CiGvApMmj7M6qBbhyCrfj
qhCsW9Dq0YVwBYy1CEVvtR27xavmKfh0m8Ni2tix9hwMeps3v9Yf9Lns5TlI4vvJC7sqz//Rf8I/
aB+T/wvTBfOlUFQBvnL6SSsSfy/i9OecqnvLJiKtqIE1CQcIpmBXJN4qT3ylmHbCUQt4VZuatBXv
x8dCQI2DRoMyhE08oKe5Efs4S5tffw68bTUPtbHsHieHPvqF/SAvoNhOL7VWLkmQaetBuPp7jkRq
66vzX2/ohKtaO3cBzJRe+2186jwTI/D1SfuearcQcRzEtvpZRWiekX64wvyQX/Yp4FRxxSAE9M/Z
/Qo/mXPzbh0C7NNUZGRwx6CFBjFYj3fyUVv/QAy0TTDVgeg+qwCAVYDbQJ4+Vbcf5HKPWLbGzLYu
3+Hprdt6NG+9l8MZqTwAxaYc7aJ6hfUbcpWZofFnvD/yfWFpneKYZrD9qY6AaKY05E0gnfyvSjYO
xgiIV7h/59Nivj4x0ZL/J0x6hmyNp6uYD1/co9Ls0eQRPMwSUI5GmToxvHgn3RJEZ+KHSRt8FOWD
E5fkgC6B50QFiPpmUstjl7emEjGeSRJBEJVAQaLFUjRUsLuahNXxSo1Rp79MGMTpSjUz9CsvUNzh
Cysk3tQU5Kqw3bnx9xl+7XM1rRMVfhP/hKsnoegBKwrpgFx8/3xRoTzwzW4GZrw3IefMYnKvSHmK
QDd8iUQuKH1GI7HKMG3KeHn+hajfPaNZQFV5pklmRrNJtgmO7J0zOF7HyHfMxTwEoUhUfaPpG44G
QRkZD6XIn93kzMAf9wqZ4HRNBGkiLq6AbAtHB+YZszqOYfOPjVUltiG2JPA2UV+6BIj/wZBr7sBt
DqcH9Nr4wvBYcW3o3Rs7L2oh/7kHMw0C+QoCDuQWpQ91wEaMU1TLt2whJvHsMe8Gt99xXFSDttWh
XupRdk7EAcAEdsbjnJ09+0uVDfwmPvdwaatb+stSeTT9VTguuZMnuIXfWUoTLTLvhgav2iiP8UT4
96SVogRbsANtFGxQxkLFerfawmUIoCxTbU6wOjj03s3XsJogE4Ri5iJCtG8dd8mz54nNVHg/Hcsy
haJVBrMKqPD+8HvlP/b2NugaaaxdTcdsjqDwapshsAtSPIvmYKH+wLaPnQmHermJSd+z2U0Ai7Mp
Sl8On/Bip1PQTnUt2jXzgnglO+cvKed3J3Nq6TCwLbzGs/myxSZQ83b+MnlurnqpYc3o+ykLcd6b
wG66rXC5c26LlHfy2gHdaZtmVis8JreEWPwex13Px6KP1ryRnkjkBPLnliDE5LE3xsOKw4MKHe5p
P+vm9sOtNGxZwbPB3rFCAS2qxyY+gxG+Fl+14zq8qUCayMSADshaVg/qcoXX58CEOnAYS0gk7tid
6mRy95zt/DKetjQhQE651D5fHuiFvnoxSLtPpfuKWXpUXlauew65DI9dmxHw5CLnQLu+rApdeHi/
HjaUtaDurtUKh1VYl1KkzgP6Vt5OTKT1zlmQk4TcDYrCaizzzM/wV7Qy8T5ZaLQ5owiITDFH8iZY
27OmieRQFCjYWlEPcAerwjo3CNLhsUa//0Vik3R1we1q+TrwzHhvquek9XZNX5zkhe0XIj/zPnPD
iAAtcM536ySnKEZ6rkCtqMOemDX8iIX8WsCtMI80QL8XwDo8I6Qo82tfXphndvAclBZQdZuBBrYx
p4BtifsNu3BJCHYVkk7QJ0q7VWPDTUlpnFrDblSCbOAuYA9dvs/e1eBpefnZURqavWIzRSj+dExP
3he8ClXAll53S5bnBMkIiy8AHFaUcHNNVemOpp2zslkZs3OF570T/Jw/fFjcxiJSamGyEGZryrwk
tpuRX/GON4nnNOJ/RhdoAKWpXidQZ3QQ18EKWuX8YpsXaWNXh73iM/QvtXxe4xB9ZCbzHDYVvO8a
ecIg7hTMha0C38T9IOsdIH7L60+JjQdmRp9GlBHTaeYpGAcZ/tR4BqWTxZ96TKdF6b2/xDFw3c0l
vBNrf1GyhGImNRHgTaELaMTrWrw5MWbGYI0G9qoqCZJjjJoltvyhDcT3Hm8e9HSoPJ66Q2cRKgyc
dNs7Yo8T6Ll0eGxYnOR5DQN8qI+QsHjcmbeD0H2A02tiFifjfFSuTz2N1t8XMxrzAjhHfcT7Ne4/
Y0KHyuG8T+hsoVMd/h46gg9p+GjM5fUHT1OdK0piJty3kr+p0wQA2Ugfphwjb15wvOk4tD1uea59
rEduRvvsWwUCOamwM11A1XPZ9iobp3KU862lvtjp+M5I52ugiN3zke79FNwrmWNkyKGWhO7wdJry
rGzvXsAPFf8rpTpvijOLdar/blqk7AIMsGjMqYqckEFP2sVuDotXhKH7GhZRDmSyOnIR25AbURSg
316TkzlHezu1L1y4ZuZGFsU6MuqjG4mjaBLBrm5QVYvGoZnO1ua47b+84mFQV/OM9oIXA01n/Dm3
YPEitgOZbw+vkN6pPJrLCGom7Cg2kJ7KtvCNQKqFthN5qGCaHjexmu/9CIvn9y/dwRcFKwJRAjYA
XBSB9fSQ4hp/AVuzgqy//Rs187mPwQ2TO1YMk6aRj3L4WfgOvmyplHnXYAizcvw0EXlDFs8aol5V
WZJ4I3wkTyaSAZnCY3p6wfvEhd78c1ZfK2hdz8DbeUmMcrhE6L1GwjhSf+GkJu7e4yeKA92wjskD
ixcxY+XO7dgrt5qZ/+qqENIw1lUcCZb4c4uWJibLJRbiXGc5+nOL/Lva6qa41+aTlaA4d3Ht4v3n
dyTxLQDnIARoaGs8AsDlHBMq45V/0xx9nGrrdvS91LB8SQ2vTprW0q88wF97Q/VE6EqjTysMdL3o
FUpgkWlQQ7p2XCDuTne7Z1Cp00hwSDU1BSg/GXoTvLBUxYE1144yCFfyf1UODliSLTtUGKRfYUR8
NUz/D5aO5cqYTOSRfNU4CRovkFydZfOHzNsS+PIhwMJzztCQT0y/BDrw6CTXL9JBWxxyLI8xW+mu
OHOVtpXqocMFtuf4wxy1czkB1Vcvi5x1RgPbRzKHUohIpbDdFV24w+ztzQ2TH1taYEFFxpk+XyBc
NhAKovd5qEFqz5IxemEYRhJ61/+5sXyTorFvd+kaPSIEQFxS78Iu/zPPJMG49qCbxs50oFN/TpJJ
r9ydenCydy7PaMs2wDCVte7TpgPxMadwHnmGLfywJResvtlD4tkQyFIhSitqSm5vpavRcBVGmJLO
aYgtXyvLzxBtxLKG0MuR02i+6/t9MRzq8zwaI67HvvlNzQsLvLnvtMdICoCSEX+uBbX4fvvlyq5R
mnlK88td5P24PVnmlU6QIEZVbMjaYL/GJKxAJYDbIK84DksI77Bxjv6UA1WnDi59OtjQup+SuEtV
mx4g6sgjGo3Mj2dnVdORTVB/uAaAcpdpilQcegFlIVLHGY+/VlFKJdxLXayYDbEqCAePXbf/U0CB
QJq3kE6fCI85XucJjR88N+Nt74ArsTEGsA650E4QF22AwmdoV6sgMhjbjuVPaM5igNCWfj06N6Dg
SRt/yuTvMUOFEL0Kt5aNo3mZbH+kZuztSXoNxEeQqZoH7OnvqxgxOjkJJG4v745vzuaLm7CX/6C+
O2n9yCQ2qKqF2fJNqn4lSCl5dW6Hu3bbzhbRMq0IO3I8WNvLA9eAE0VlCGG6ssbNsq6FYuBcaEiI
qrqaO/7kVbr3j8bLyPJayBg0kHW6ul3e/NOeljXVQTNHT7PsipkJyVPbd5UxMKZ9acEe1MA5WV8h
59ohMlatUdB++Z1GiHXLhmJrsbfBOpmlFife+7X0Vp8sDirsuxBK+BHc1JB1+Vov+iqwE5F7fN+v
71U94dKfMpjMogHq0U/tG8DrNIZp/UZ680B41ghdIqeDY5RQbGMWv2iFi9on+KEY53ONjOOZy54X
Tt9Bu+zmQFKpXNijbIjyTKdLLo0ZUx0Z0CINeBShu1vTzWN/aFPLLrMw6IOhcOgAGtqpLTHzUCRi
CoSozpDgyElkeicgCwDCQ+2WxwyJO93n1bIsUp2KUDEDcQ4FXYWvbFKxUPPbluVPZC5X1rmeAq6q
o3UATz9HYp38bSueNlal3SEuVmY9rvrAOf9pjww4APbRWKAqkb1fpSqUXQTACGyFgu0b47UdNddc
pYy7QZ9EXnGtvnpHt8AvMnSUkb5+WxdKotIwoY2tIGcQIfu+OUUJI1KGGmT6FiEEj0GlwAfz03CR
ylRhlqFhXUqy3u9FEYfVyExNyMVSsl4bV87u2U/KfJSpiFPetqZDmcgqeKR5IhNoy02ZDnUtF5z7
tk1fOctizAz1tPvT7E0Q/mGsWXTeTjHxRS2eaedCYtQyRq67GbXQUIWP/io6w6pkIjCTW/+80t5T
PSyeVrM2aK5ZP+RIPvGR/WmkAXd/Ywzn08GgWr66II6tqFJPN4c8E2dXKYC9/v92C9Eh1NIfv3C+
GyQTY5gYNQkU/qJcCaZqZWua6npJluBV17vyq8BtXPS+GSLwTNm46C1X3vb1BTK8ofu4fAwJdSxj
tHrEf83Ky6CUCZs90EZEPiQ+44ehUQxl8wk4JWM0tDlYlTuBkhIzeLv5Kcgr5eNl/PKeSiOi+YA5
4bfaTx43e9SInNJCw2kPNfP6pdHLwkF5huTQAbhPGr7Il7iOm7phu5KwbKQLYCgY8EL0OV+fw8ck
vcsARa/bBQkSHgEfu3goJNfx9VcI0+aWeGKvWCJ7Yw62i+hy7NwZL8bJnCcZ6njl+Z1RgRbZpNFr
J5cthUUsTFWfUP2qIP7Kh+iNawqLocn7xmjcGsv86Jas/ZeRFkTUjk3etb7yiv5/TeZRWQMs+Vrs
BJJUq4Ek3PVmZ8gbPDM77VW6e2kS/gD0bZmq2lVnm9oSJGvKsg0W0EqRSLDMRt88Ly+AET/77s7c
TntEJh5Nehg4sK8vj8dzGxcAuRuvXkgnb2P+7gt7+SrsDMzB8SSO8K/rBNgI3pdqDx3hho8fhZEJ
N6+3dTOGSxfyxoYDqZry0G1bcdGOk88OybfjE4i+JSfpBfaLf5KH+sfxAoPqz10kuF8kfXxjaWEL
GBU5KkrRNRTead48txy/yYgSeRQHQnYgo0IHeoqA6eCCZWwcAaG6s1kM4Ehz6oMAzMol4Y4WNAel
J3LEu/aAXa8fSH9qjHxw/NdxcCk88R3RN4Ats2BOqMhd1Qmj6xtln+7CGuWEiYcSEwwigpfK9eI9
HcfzHzxdjaQ06CJauFmAlc0LrzIGzTkZB2tmx4K+d8kdp/26cABSzlRXjboxxbuy9V5PDYXhDgfi
JSgMM/emmIRKi0g99ooS9f0nSLE46dGfqZYEs5CVGy2VG70uJKC5HMJpTkDaKhLZdJsjL5L1Cmgz
YfRJeuAVxvKdFLN1d4ATmGLX1FRTR/dCwhvfoYeYdQYLS34bENWSOMLVDTyioPwSeC+bQjwqNe6x
+eMJnf6k0+PIBt1bO8oFLIsBFndIKCvIa6ihxHG5Aun3xYEzktE/G8RDTamqtL6k3YO0k92KLLq5
QVRuQrIEAPd33iRGGKt2HB5M0wJK23Nj7j9YmugOLIehaIfeKZSWGBiZYL5YwSmg5pNWculEdZQV
XQtgoJLySSxQ+F4PLz3cyt4iAZ5nHtR3U9P5uEW0mZkDHREfzrGvlu0SJETkd8aUO1rZRgyqnrJe
/gLNopAmPPp7FVcBNsxCzo3kqJHaFqG57UtDhmtOllJqMNBP25Db7Kdha7E11SxLvTSpDi1RFdbH
BpE5Apc2oTNEOYRvnVhkvSyIVERDz0x9uUjc/a0LeECOw3cjC8GQ1cmQFc6T0hIEP09Ifva3hNHZ
xRUp5WqjCgcg+YJO9E2yQRxkVI4DpTShGx5x2fXt3tSEByxwUwsD7HUTNrmrr+K1bdlLDMFURx1N
dKw6FUjWVassk7ZJdCJcLgy2OY10utFCB3vl2ocA+hlM27T0QX0lhUthaZTWPRnJzR81VLjkgz3i
QBtgKEsc1wDsKbNc/yRBhRqx6i6JFsKz2yIrNys8eUEOHSdxWhhif6SxDDfOt49JrQpBW8lq9Qmj
AdTZLdcNBCZ6pOQE5oCB4hx5Czp9IQaMqhKxCaW9p38Wdpn5MDoKWW79aiWkcqpohu/FIBAZe6xb
qQY6S6E43trPJVWwYtaf4S+lQqn02LkaOBa3vqyf4qT1y1n4cvYmv+aQg6njKAUxJuskN2yRMRvY
yT4piqPoXfHltoGQ/e3w5Y74NxWya5mqA3NVeQx/cdTSi7ai9ZnzG1iwEGMYK8DJI1CZhCkNJ0jM
GnXfK2sSSwKabkDQFo2a6I2jckDaTDDHMUEvZk2QL+UjpQ4vjcmlPq08VnsKPhHGseV6MABmo2S7
f10sDv40A71UKWaH8Svq/Ok5iTw4e22lja5h0rvKmDCS+OBFWcnoKbmNu8/PxCf201dHHzS9AdpM
UEcdAt/4NCuoTH/d0UU+5Hlm0Gp0rXAVWz2fcSbMpoEroxrm984e1UC/DOspXZngtkv5XpF8nYd2
3Dx3XN+SP9kPo0UyWgR9nvmMI9Y6sD1w+vlzCGpo+b8ZueD3/7SdcHtKcJ7I0LLHE1OOqAqZDC70
qbBc/AxrfhDphKNKw61WRATUpK4LFgkcZEg3QBaUJR8NK6LMqZAwzupMXa+KaHMTHr0jcZ2/1St7
nT1iGwd3ntABzUXS3kNUjdQnHyZOl3qsT7Z8M1uQMPnuHRUEnbJ8kmS0YB6iupIBAAOilyWs8aVU
kHSbjxNw2JcFR49FY14LEqRyK1197TfMwHA5cNfwPK/RQqLG6Wm3efSqemYu9HOAP1r0vO897R52
69G75gu8kPob/qkZPaDRogmYb5Rs09DNywIG9trnGLtf4XJ3pRW7wdKGYKTlAFUW+5Ck2m5k1eIS
og3wZkBMtt0P61hs1XCrZ27OuM86HgPWdOskYRXS+y1p0ITJBF0s7qBVsFJS6cPE2bUIpCiCmRHY
G/nrolWrBV34ImraGc++4yzVsgIfe7t6ewCj/CahrdVJuWa9loPXEdR/ZFNV0/8Jfm2tZJf4G9gw
rIagnt0Mkbxd8A40B+PZ+MmTHfqwz98mQQpX98bRf2LJAvgqyVjZgN2zzm6SPOp7acFdA7vSMnWv
dOhKvyHKDgeevFE9A6L71rZ5XkBoqp4f3uYr1UH9Mh9d2egyjoB8HnqrsLcNl3wIbDI79hWtFOQp
R0GnIjErvUf3Q3Q96MjYl0qYqEmHZMG+aZteQxdEHqLtnRkjar56W7awrzmkdVYSfBEQjg5Nj0G8
m066Sc9waNKinY6OXQwxMiT7LhWLX8e+hoPN5IyotMFrtMieKXmwD+4eoA3Or8vcwA8C/cCP+Brx
aJIybEr/ZVGL1HPAXP7UzXSOql8ievdyJgvS8eQKsAaaMVNUoDAIoA3CmPXoxucdcxOTZCNG+4yG
40jS0P2ZKd9D6dJOmJul+ZfUFmrlHEIeqFEPC7/05jm8LQIJOcyhZOXCCpV7/a13wu5XvnNUc3df
LLK5yfqGxBqjIH74SiWSdfRzzpXU9FRY5/n6dP3p94JqLo/mSFCihtpkmwPvrtJx8j9xJeS+Nws+
EmrXiwemDHSOoUqxZcFlzmdVmo1k7Tz4dz7aRdbj1SA8TysVmUv18ETw6h52UTwjZldrtwxo4AXw
YVrJZ/b71YLoCw5cTLlDrqHzAyBZL1YAHaOek6UHi5dNJiOqeQ6GPmrK18wWax8sWpZtUsL6nxpN
QmP0a5xH+1T7rWkKODTwRbDDk+o6tM+Fc8hhPNL2pf+K3fOc3gYJdLurrflnjsHifjBhQ3jis/q5
URy2HFdKUkK6YoqxBOo/AJauMcYhR2VLYzOprpR37X6snFlTe5Np+q9373DaqQPtdn5qT93w3/2K
fZOvpiZKo8G/7uaShpM+bLIPSYFIUkRKD1CO/i4epKW902EHvb2Wc/rVIMhqywaWAjjw/QuGLsMC
v6OvtFgHiRQQW/rqlNduYGh58nc3Xxf80j0DNxBpNeiG8N6wFWnJIJGnq+xFBPqaxJ5PlVCYfAZq
P7D4I59ExIfLTHH4kRRrvX3q97Mqc2CXumTEfTfLRUNkbubMHH5jYu87Em7xlZUubQVI4Cpz+oUp
otbqPzPe0qRMWjiWPpY57uPHv+cxq3hUYQHGW5n7TgO28Lqlj+ZdXmyLF2xrLJEkidqdAbQ4MrD8
XsBWEKhCO/Xb3f18RaJYS8wPIgFkKX6fWNzbiXVkhdIfem/I7BqfJvyTUUJ0Im2WM6ayfvFlhDcx
7dYCKm0SA8tY6jAtcYQcmab9hqIcM/o6tYO8hF+jqleVLvRBBRkx7dCgsnBPnMDngcQ0NCPmRQFX
ca4tR1q7KXeODuw+SERk2qN+vNQn5TrdIxL5zJVSATlbIqKOuRR1TOu9+g0uBQ2PmweZkv8NYFny
2l85eVDl+NKrY9XmOxxgaLZC1ur2vmLLuVTL/lCGM2sLUPMiuTXrf08B37164FJlhLKB5/Iv/uJK
pHxbCQPPE0KqxlpcFvCcUPtaI3t/l4VvkfJKMwokgUmXiRTfixPRAOV8CvZlOImEtUJK30QF/J46
gzje9U3H+L05EIQGAph6FIBb2+SAiLRC2pnEpiDABmd2EMsin5nuDJrxuDA5H/3OnxoJaeJtdwE7
pcypWeLdS9EHkiF7tPgVxhWgDwYP560uzGiRYuPikrm+ZrSfyQrqPLeSnj2C9MgqQqNz6krw1D+z
PNwKeQ3kmLFn2KZ430ulaG95mqUfp862WXykLjfUbXCKdZ+PlHfRaeJtUDVf02kr0rhumhuFVzAS
WMeCCc97Z+lLskRyHvp6RZiAsKMYZhlzcLNxikZY9+z+YsNla7pLwu3zv8D08bZUycOUkpHwl6su
YDZInRBYASOzcYvfjOlSBrU9jSiXHBvlASMUC10FULqHL/3+hRKQlH0oSHYhd4WbCcz4lBkSZJjM
PZUfkVCbVKOD+tNV1ajFwZFuyRfVypBnBt+V3XH8F/Wma2Oa1LOKPmqUv2X+eXRiRTNe7T8jYxuL
tVLbtMP2QijkMYqnh9Lib70RQSRqXlqysGF6kwuAToV9FwNpHItbkyJXFPZsCvlckTilPVfNiNUJ
Z7jVDjwARMwEVvBhLPiaBzuH+Cj67DF0PvDWg3shoHA9JedU5B+EQHVS3T5dUpAr0gB129eKvzlx
YC84IDcD5+anfaUuKSunCBC3mHMX1aBwgdU8ItzqYu+7wCCGRRvk+dqyLZYDWveCxVZNVfR7r6x/
TBSVtXKtKMDbQHqhkN6IetpFdmbZ5lNnhSUEW7zE+rkraWDQJiGGtZO2KyZvLLni+Cu08D48S7kW
ddl5G6X9qWKoMS9lAMbTn56D1byy1h7F2rTNDhvfnueCD4WGnuMhfT3U5g/Wp5OUV+dm13D8NYuy
lXxv/fvOGRvOM762W/pgMVrcKNw3GkVX4d0TIq6vR3uA0LgRELSp2fdRr5IVwFqGtUTd9TvCi+el
eUHhG4HcpAgje5JrL+JhzVJzPP0/wcmY03Jujrmy7ASG2dOhqeQzvO9TcFNS4npV3Jzp6qkZ9zJ9
ThC/8SyxWLzOiGLEre0W4iaNHawJxU52eXpSQ6NPO25LZu6KWFjBMxv8P7Lrh6ck26IjAuyyUtEz
DnHsezfGq2mDMZBFIF23UIoknB728r4PkSymPuYcHWi1c9yFBdI5AQxYvS6ofKTcvO4U4wDbljMx
vaAUHMUKrFZLAYkp+TuQ85gOy/MJOgPWI+6sR6Ixp7Qr/a/ctVkcp4P3C93bvxrFzyyX0IcLnatq
pZ6IYKMcEhkTPNh9EFRPtAYK0FrgVHaVil4Savelsq75OeOG6KOx2UBUh3HjKgffLYQgkM3KQ2Z6
R8cCDcqKZG9ue3rb0HtnxYO7TxhNrkyvKGaoyCVEBAJgk+1d0EjuxOyK36qU7X4hc3O7cCWmnaLc
hNaXgdGm9QbPqTmziNZ71Y7xSBtS4BIVcZ4SYBYsO4HBsbRjW9KWjqSj5VGkIxfpiQ3YJaEJaXnR
R/G8lztdB6qpkqBpJLHnIjPN41+MK6ntTwSkPqt/7eWs3Rs0RzHnQ3VYf3RCqA83wJIEJAysOEo9
TpmAqHOH8FgUlpAeKAZer25HfvzuWphl5b0yjcRWJFEymSyqHDappKK4PD8osXdu5M8A4mHvpHDU
rVhRSu9kzUmquPRm1AzMBIWyJtPvJQysu66Z3Y0g3UMe4FNUIgTN9+pQc1JuBQNZx87ay6rQ7Fhb
KkzFoWfEGvD3MkJqTexOBRSKAQOQ+v1lh1YaS00bzYS0MpaXrhLiggd43FD+S//9lkwUsSDMF1eb
5lF31W50bRNjDVC1whAtDDv7g8P59CuHb6MhvXoqjoJuRxGIXjUVWMMqMU8PlFQMj8qlVKJXS/LF
Kzf/IUWM4pKT5wNYMrHxNwTkAXcXdIjfTkyQ9ZgBTMASVUaGqomV/Lqg2K4Lt2cu4s+9A4wDTf8U
TSJllDoQV/bDp/rt4wCs14yHPt3UdfAwOzd245EUm/zQaqkPJxkUIMc8hgVPtQ+INUsVcc8XXHEh
6y8np9FlQ01tyEdwIiUHWqJqDTt3xhXJHArOGPbbTfUzbTS8FKT9q1iIDoVEa1iTYuvFfxwiO5Hd
D2V81rpqhgm7AfA0hyEDun5GRlMB7eVZnI0e6Tlb9KrZm+gw+0TA8U4gt/7T4aPD2wFKu5zm06bZ
sK1xxXS0iiLcSBXdnE4WC6Ah4x0Al947REmTQToBcpvJVW9fDfS6kHUig785AS1LIxC79sqHIOQT
DeheEzMWvtF9Lw0sZXDQ42x9ktEL+qMk1fdWmcPNvs5scouAMByNhSof5/RVhxLTHpabFUUIrU/X
UH8VFjBM4SEjK+lT6ZDzzMr6bbjLmIshGQ1XDt1wH/41mxrbMjJyTF4UI0vdtC0OzBLrawnyhWEt
B5uSJ97ZxOZOA5u5wk9y147zm+QKnee2q0YrSmP6sBzbuGqt1Hp1molY1PO6fqE5z5vGQe0f5NHg
mQfGdtKM+u3Vo683OFtyTH4JXDb67P/mtvlr739UM5Y27McB0GxmGyjHk52Q22B5xrFv3YyWwkfG
TxTkSfyuEd7VuNV9H3w/eIwidONZPBzxIFxQ22X5Hy7bx7ixf82+raw5+nig49cR354lNLXTHofr
fB5Wg9oKZ2LTGbaVTAuW1+gEfFFOk829lcN72jC/G02HGU1RTxvGlMXCIlx3dr0hP2ml2Pi1Uf6N
D+zcs+yqTd01pKk7ezlaFFqV5dzaqmDdzIaH540ZzzDDHqfhWNBIjrpf3+IsKK97H3LyUlDKylIc
C0/FiMCTUzqQpBrytowCd1qF1EGXkk8zdvdYwN63UAHi9J1qOR1CwVCm0UYQ6jnOg4N+Q6XnkciP
OzPuTmWalf7thMS4brM3Oi0UeAcqFWOBFQ/d/EF7bl/yXrZa3TRZbolX5lKj3bRIYCEBCPlUstFS
c9mUnMDOlQM6iajiqdzZXLVckcFOhESyxa7x66KLauyXNsynkbWBnFlvtEVUMgiabjy/K/XyEHpO
yP3EbwZl7yH9AjA0hcPnxQBVn+CFZTnaDr8i+a8a1RojPNsspkMrpczKa9PDEtI7aGEQ3xSJZXdh
06rD9kWKHVDwwa0LHm3+okJ2jzP/NTfmLveB83otQVZT+DAi0TzajSDstLcfVWVbZD/X7KcXP9f2
K7keH2BJvO8J3shQWW6cUh9GlVEikn83ybApikh4CVWqkwPcmPcxABsLIDxmMpJGDuehVAA1G8/S
i5ePf2eLpl9dJU5FY3iCnN0jQTuok1sAlglV9IS6oJfmrrIF/gOfFdFT7MlGP2hFDol9imBaT3ux
R38lQjkz2owHhZCwVCvFlRJtVOQljX/wfmH9OjTZwDiM0YjwelUp+sToQnqHA0lSevmi3pFfoVUK
WIKaYdf3mcmNywaA8cn9EH6nxiJ+GFsJbIKQGN46ybSj8Q7oTjyD6t2Z5BfXZv03Ba0A4G1LK/If
EhVBm15bu39VagxkonObV0r6c0gnl2yTbxPbpSiswhWMc5a3/akNhv7ESMjq0dEE5Q2yCqCcveNG
6/aU3P5gjXB28AhmwHg5ZRkDJs2Xwsj854kkMGLDXmI0ZuLUt0NazkgNBGwDj1DErYT6zn7GjQY3
wy7fvH+ITj7f3HsfwbXyt+rMVdCMxJC2lD6PkBYwZvfdYtZBrjB11liiyGdMKjEx5wqOR5GjYjcy
RN/BDyKtzJke5ETNmeU8o5hgSJB2MuhagwWZWbxRRZwyzb9yjo4amEXPG2fjswa4H+utHloOUZoz
0NNF6lzA1yCgHB3oZIS7mPXjjT4fwL7ZoGvwBS5Cz2M6MYlYFsN1Cgjwpen17UfUGzDncWQ7dgsX
oLTJV12JZKUT2IDkNTPidVYgjyEvgC3eC7S7qLhoshJDYDEVHP9poOn1khK5eRpjs+IEKIYWEXLP
oLmUMTBigm5p+XRTvUOVBF/k8xG4xxigaH/r5BsDmxYvDD0mQeDUIsvlA6h3iqAPa4f9SlqvSAPs
rurARi78+6pvKpbBrdBXDeuAlDWDSandx2oKLEH353X47TADRx7Ln7MbIywWIQhBl76FlJY4d1iU
xrDu/mleT5ceOdgwwJ7r3UrYUQhovh/STyfDTSKMDhrK6j1AJe0kcrEizpoGH4uq2SlBc+wyRKZQ
h2yiE3XrtHHcumS7rTSYm9uqigcK7xLqCIJzU/ov0gLAMg/4bcOczUv9HQPTdJFtLBelj3MYp9tm
rDDNiH9nAvlvMaknChF/9xlDdoCmcECyS8qtQvQHQJI3SWmACyM+XuyGUbzuCNs44jZwEnRQifdL
lZObTd7CELEpmLbvq/C7qZDOIbmMEOgvxIQAjfAKyg6b7gU3zSeH2+Nwaclvg6+qK/HldF7tKVK0
o4os1/v5A93mpBEgc5cHc7TEZevogu2TFdZwF9U2fk/U/Z1Y0roGkay7FWpEBn0AtsKzxQaPEjqZ
7pkF45ED8MzVpAsTNn6Ss8v6kY5l4BBVCEU6p+fwG2O4fc3HNopituoVm2mR5LkgEoprEZbJikk5
HCK/4dGBkMyRZpe8khkqG4iL4U9rsvyZrM1QpYue9F+kGrX7elaHcoWX3wvTE75A38CSijCV4uJv
IWt2H2ExmEbfwzsaRQ1xmUp3eJpSyP/AYj3VZSAptXNcCWKU1J5A81WwBIW740BaH26YKu5kmwGt
taFt4YE1n+/d8S2qG6R5kAfczDNqgvkgwOBzTHg5VBptfhPipRhy6xvEb63Cvm1ycyiQSk+/BCjL
oao3CK7GlogvcoOBD524VZmRlvU/tCf9Lyw4ww0T3xKeU8ulRzgzrHFo4uo4IPaGZZym4MpZzkJF
rGosg31PvuzetZ33kVNKghy6rmpRq+J1jea09fF9rzpMQjZKFMqZXWsw64/t7nlhkdFUIT9bDJMl
TnMLa2NCqgBM+VcM1Md1BmnpJRKhtyVqUawxNRZyFnB8VYUcnmVRoVI8MP3YK4oe5VkcyGrnILJJ
iYPU778180K/O8M4i7KJOMer4oKp22uVpnm7GpgnWlD55o/RvEkQXauK1lt4gvHW7UxPxDiLh+wD
s8CZBfG/PljCMKRwgj8M5uVzTDBF5mHk/VbxRXEZ4dAB/TKtQMDzqxRVPBiTwKIz+0OWVgVzTT8e
DdOpBT94VL0XIeEN3gC0APXFNQEmA0ae6+EvMQDzBIagVvhzufLWjdHEJEefs12G0cGXUe4cJhkD
HBWEW6ihvP1ZhyGj9QD+ZaQxGGS2QnSlPs9Sa5cQzlzexprNSZe4ItEHFxcU+2GVrwtdqVNJi6NR
FyQ1ULo5RJjZ/FMRStwJh3b8izpgzBvTOM+3RKvaJSKcYodLnLukJ7gnrs6I1bVY9f2Q1/Lo2FHU
jUYTsiX1mYUXpn6AKRCIdB7YMxQ/YGCCpwjJY28nvpFBgbUVrjfSza52nRoD+Ssx3n40qIXLVORK
ya0XlLDimsBvg9I6E7o+Zvbs5DkSAtcij3INA908pBQng/9PrBTipX98TSpEPfSDW+uDZ9IRhP7p
UiBLqe6e67CAUwrjnrcQfm772KmUwsQVnY90DNeglEhQ+aPMs0BNCsFUyCCf9Iq0FyQjAUOb8mqi
sbr23eJ45JkFkLeijwBTN88unOUu6fpNM5Xcbvv5MfUIYGRljqMO0MOgxWUFB11tjPuZlZdtNPF2
MvTcnn1npG7b8XflnFPWsiccAz7pMDaDX1bX3zKXRSOyl6FRGKndiGvNq75kz0yN+MHryi3OJtwx
l3Kig/25pg+XPCS2iUKiUR27nCl5lFyFlCAUgGsFind83EI3Z1irFmlz1lu81q/7XvDYuuoZG3Nj
xQ6QX0mmex2MR99jn1qa+T9SDOLBFH1ntFy4yIA4wDaOsbapZonlvkWIZinbcANHavxzmUEaUPQR
wdMWXlK3B236s7aG6gQ8xh59M/XtzpTGYt4b9u6mvBc8Bn9EY4W4Z8IBX/ebgLnIq5TjIEth8tX2
shRjsWP7PLRnyEwE+seaWAJeZL3f4vy8vek7fAkj8SWd7RBos09Ib2V1DKZRju9/F9Kk813G5Yrk
hKUlyE9nHUrilrSlHavmcZKWbcoiwVih8MoRwYO/aAh3OkfaJfKV5oOLceIPNXbl7Hmutzrq9xla
9NijyXM8mbH65M1weHHq1ZrnGT+31FbuQBw7CvFTIhOYhUoBa1OMIGSViO8fn92wEcIfF2AE4onT
iS0jy0poeUcK45/Mrynfq6sby4pykWFolDmMGyHYGEU9QICdlwjrAvGACyMCQJrS8WE2V05Umnqt
33KhFMkpYr4jpLMkW9FPClc2W10MyJWtMLc06DQlSboDOB5pdFnlj0xwbqxKt31gW1f5a6vIOz1u
hTk7pMOWELkqOIs0RCy1FO9Mx+40vfddeMZKBfrjMWeRAuCt6ALTgn1MyipggLVussFRghMWsTGz
rsqoZ+QlcX9o3wdVMEww13rkUai9uA2vhGWYUUKwLvML97GNs8Ul4gF5vK8Fh+Sn6xX2yFCaVg/p
9MGoxFT2q83LJm9vvI4DJ3ofmn7w4ZFpghPmgxq9Bb8f9waS9pNehrj6Sqi0o6FL5ZDfnMlsrXyV
CUYKNdAbnGA7mnqq8BgQqjFPdXObA4NKaMgmtGkjF3pmsFYL0fFH0CMHNGNwP/tW4Gxl6vpA3TuZ
7VM3TpLN/HtbFWFD18kcW0fSvnDeH/i65eFHc7nPoRG6KzfB2x4bW+QK/B8vAuTmrKGCvi+biu3e
mTL6IG0u6aswVrDOq2Dvm5JFUJT17nQ22wG4iuGg1YWTMsRBB/10CN+4tKFbJjX769yXPwKQzqXe
V6vGHMC/WzSNlU8S4bYegR/HWuEz+8XovKPockd4uGBAofhY2ksfx1f1mwLbJDWLsj4NIN9YaZMc
D2t0PvZ+o/HJHVn/9be6+Kw/zpQYku98O0nqkIk/5xIul0gZ75AzhU3d1lVe39efUtMOAmdGo4+F
q2i/PKFjM/2/WeIAEcu+vMwRDquMJftc802QjT4q7LMuP61/dohvV0FoQbjz7xL3X7hZHQQdE78a
p8vX3yJoWMes5g15+JrmZDO/wJ9HpFsCXX1bkvqGMx3wJXDY+Yx8sl14ZsdHWCxE8qCd1jiI2A1Q
CRFcBS88K+H9JWeNmFcFN13yfZJobkc7D0g/NBXxw28zoNSmgcUYs58Y/dENZDiWxTRTT2ATY8Zr
g6oaIzTZYsIrG7RDkEqSGLmeF5sY6JCXY9UtN8mnvgSU6i+C/vVPr7aW+72QXGjHmX/Xqmb611BV
xmmTZzazv+ffVJlmUYQzJhtlE/gplnrHEi0/BI+jFB1XL1C3SHqV2iidLozCa7RjAqckBFcLGU5x
EaN2A83v/Ng7RymIcE0hIKddgx8t8s1Hi9ryMrA78tnz7IPMKoGy9RnB89+3KlVJpMQRCNq7r7o0
oT7huK7RZs5XxSaPF7UCOl8uVQRY//yXePXsGSyJ0/6o1NsfR+VonBhww1PR5zwykA7G2vsg//f8
LO9dg8hwhNQB/LvEmmYK0iR9aSrOpe4jlTHUKn7gyUQq4ZltsB8jdQxef/ylbrgfYDZmmngdU34m
hSLcT7YhVt208KyQACGfeGn2yH+jg/a/WE0KjHnPGM7RU4MvUZNIZZmYH/nmdHl5+ChcVgqwiH0u
eE3ArBKY1JZoO9QIJe7NtC9P2qUdkQ3pk9OJS6i5FeY89TvHGNx8XwBWIoSuDRwYmC5kwCZTlBW7
zMORoEZSxCsjWbzLrg1vW7/W8RJWIYszCe2ODtA1D6SM1FJ1SxnkVHKRatH3Zi7Zq6I8VTGK5Ah/
wH88KSqt7T4QZLvOtu89Ua/XfP2F9BddCOQ7SDZTf61ldVEXwO+LDYdk8hFwh5qIVWUBuMdeM+t7
tuM8XMhcYFcPxWgwm8yGx/NxkUVr6vSfYy08S6GzV82zfQ+CZ5RU21zEwvzOQD+7raMhWY1W2kJO
zrtKiEDIeKHLyrQ+PGnNzivnVPLygGg56SY+qDUjOt5fmh3eaKX2naxmXtKqraxquk/TF7YpI89A
tselo/hqX6jxHX1GpuN2FISbgip1YhsOo0rZOkpVB+GndY7AbjGCQPhJUAlT6f/YdriZYnaPTHWM
1EqpCJseLT3wBz23+y3NCDlk57QYrfmQrwDgoOG8VbQOSXa0fAK1uwE66hD3s/cwYkkkfHH5gGC0
ihPO85G47ZGqTeGsIPtjJPF5vEauguXTt7MQPSRh8/cEzAEP2JIx4U8jYr+Azhlm26i5AsoGiNEW
Crm4pfn3uylA+79Vwoigr2vcGiyoEAouEzaTx0OMtlAQ7n2IAQ63mmJINKn6nRohTFCljfl4i8P8
HtGjZ0nKhFAPTWu3b/9l9+ufaqgeEJ2Q5+8D7CWwMzoC4vm12shfL4JTG27wi80V93WokLTuxxjy
wzq4r+++gauh1nRKP/CxLwlQLsXeXM6ihKAA4ueZwClrlPfxr5RSnMVXPE+rjMJiDcGgijiu9ynd
Zpt/tw9aaeTanMyE1Huh9RT5pIdLlXMVEnplOGN4MMZgAK4/qKFYEK+JSDh/xx6nZSvYziq3AMgg
x/giOEOxsi8DWdUPcRVhnWteFffjL8Sr3A5BeUJmZxneykLWMEV3IGhb4q6m00+pgUkOhsCwRQ0K
o6aZbpDnnj66OMfBKQygq7H3uw9YE4DqgICC8I4IoPHpjgryeBKz3D/Mmb0kCUldIcFadmaHA2Si
WueGnpuwHZeR+Xu4SZzA0aYFN7ZpcvdYDV3iSJjJ6ES5NFFlVt7UTBkrp6YLKXs7d9wWVnzYKsS4
VSsV+QJb5BUiJvVuB5RRnUmo7TmIg3DjDOKB6KU/JyAc3IZTEjMnGTp11D6ioUjGrWrtVNQzKSFh
hpKcL9ms8fRI43F3W8nye0L7I+T3xkAOr9oYfoSgSS2BXtR2YKHdvT10XoMurwIS2X3VpguDfdCy
TzRpsD4iAr2jyDvMjtZYJGYupG+P9+rO+t6CqLsInF1ksGZNOo+tJwMTU1xkE2nxy0cthrnGq5Rl
gc0ZOEQi4jzDecfHkOY51zRVBpMMzTUj801o9ci9Hd0DmmOiPtFvxDNMO8RGFvgSbw1flgzyRXmf
2uZdYSWO12yh90PCavWe7YTeRY/Dm2m++meHJpvmDmKxZpIL4FDOXfSfuAc4wNSpvgi5fddjUhmF
heCmIIcVzf8lQHttuUmtt6ANqHs013UsF7jGyGMMh7qP582PR2RPBsbcj6Q2weEslRugzFzYlgL/
j0VngJPx/aMojohjocwmM8FQz8EDlN3SXFjBKns/6tgA23afIDOnEaxlot0MxYfIVxtmbM1XjOsX
29TalbnA7R+tMvQCliVvxmTlwkpaSXmwsm0EIgrDAtTZUmdgB7TAyqrsALUz30aGyPSKaof5F4mQ
wx3gfN85soGpB6jOLNATjIWDgVXWGiC85vvQw5VKuI4iqatAwaThXX8L8bmQOKr0JcpIO9KX1VrJ
/98yWiveDPYG82NvUGOKJmrbuWfH8HlMs+NJZ2SrmrCRsMVG74eh1zBhHHSv56FjCAwOB/tmuGQ8
xOKhwcU3UQbY1PFESJFMWZkM1P9jI2HRWD8x2jh3vG/hXPKIOMGNBwI8362rxG2ButRC1YdXkF++
/7pGmrinZTishgaVCQ2xQJ8+QYtyke/bjkIsDwdCOsqoQVEipoOF0ex0VTONKW0ae6jaI6XtS/1K
01TkwvJqPUy2Z644bxGy7pmSAZkjRDv4Sdy5SsGrkUzZA5wradxmB2YzzfsIwTTvxKmG7JCkG+FB
xZA19nKvT6tjK+Pll3IMSX1tM96D9k2Fk6k7AdVjulHSzi2GS5r/jqZIcfi76MwpsBMsf6xE7E+S
P6iWTAT4d3Rs7y1kQmqkJp80k5nkZ1woXySHZSaLUQKBgYR4wl7Oh086MnKbzEv4EjqXa5b43nhu
24bh39u8PycX6HxF2vmt37aO64IROVU/CNCOYjI6RxIPO/k6Eik6xbdNYvxCq8/T501hbapMRD9o
ri036iZ40Y8QtJdRNsvDbY3Ha3NElU0365nVh+pUz70bGE2QTpzocoa7pyYcryYe+fx/nFG/pkLo
E854aT5iNomaxNBnnVq/ecxY9N1aY7T0DF1NzOE/0Qx55Q/bNd2f5XfetgX963bMemwV7xRGtAeC
Y9jEJZ1JX3tHxWfb+7kmalYZ3Uobt9tSwkNVmRGyn/xXKU0xOUfapxEr/6HCO9DD9Unb0HWlT+Ej
FmFI91bnfCG+YGpPPFpuyzOmCiI/mD18OHWMGDXyogPuB8a8gjKbx/n11Oiu31aniKU+QG1cGa6G
0Yp6PEeA6BMP8XTs73B6twGeSilNCqh1wYncvGWgi7EjJoftue+G7Nq/4yElY92ETWFR5Ivs0km/
rrZQ1zmHWQfdBXlK97DvU31niBcDjCOmUXHuxrWQma47PIl0Bdwvd4KLjbzMbkS4Rcwrjt5S7ycw
2oxuGIIzVBvs/t5Kkdmy/LqEvKNtzjSBh2ctdZ0SrrwZTHjSYBR//S2yYiltaoYGl3EsyRzx58o3
0DEzLFF/KDzGfDygtL5cRxPS2KQP7t0ZbGw5/I6CWrQXHYOGFymVYNtRIcKSwgFUam30i0aTTPk1
PdfnP8u5Y9KqaxZ5rHqA10A0enfZIPP5o2XjlPdErc/o+YLUM9Ps5zSPtCUEnw0BdZ2V46ucBPjB
mnhyw5BjLt7SmgjDq/MmudaSVI3eqlzw2ucmApxuJel/H0tfkmvd3L5Du0an0MFSAyft7MCB84r2
sxOJzSxW4aDujIoeD1uqbNbpAB0TARqnv4DCCwQ6nsiAProhyMMLCRFO34rObcEyDu8Ter+FNnpE
3GbnS+VKuQwLxw0wDRflPBoPE2N7VsCN1s16yRKkzlhea70XdA/gtDvQRMsSY5RJQcOSvbLhZVw/
GO6iRWZbdrk6xuzdtrmu1quvtXpunHWtn/B2sle9aKSQUDYjVkrChaOQl5qbTnyeMkFqYDeOjelq
CHRYcpns5hxUoQ/Sp5CP3kpqzA/2wlCN9acaUcpD4hjqMCHOr1AQ/BQqL7rKEGLyuaiXYKW+HMGc
BpYw0ebnLEGAm7/AFHotfeqbGluKGNue15Ps8vf7MGtBL9ujjy8GcMvb671EjyuCn/Nyqcy4gtb/
+5mY6EfyOwbmRxvJVBokCJfufHoBArhn2P3fIojJXy5H7zC0czNRz+BfC6TNcOGjvQMnv69VgJAa
0cZ8Br/P2rIg2jka78boceQpxAUfLRjS8IqXpFf/EPfL3CL3rW020VLDvGb8+vMaTSGzb53GKhUx
omTWtFmcYmQorEzteJCCdFmUhOtrBvtmjzl9qta7Ed5icTOSHWjeTfFgW2rXh2mI4m+72J90R6+s
fIksunLy3MYYjzb+Yw3PhQjV7ZvWsUccez8Izk9BO4k7H9aXjsRT2jiGKhOnSmo7Yr3g0VSsUMxm
T7kedpereIPqLmNCS6D5g/sXgjvfNFJv7Ita4UFJMwPtchs4LBd5ZeROtDoQZ4lN2dO/JUpUY9v4
gcRS+LVmVR1iHk96VhCZzuLUHSf6TEzHVzgm6zVR6bEf2R79RKtcK1qAtGmPP0Wf57Jy33F1rjZk
2yq0Oxm9rdZyKS9u+0XUsR8hXzOvccbjxzCGL00iFiQxThAubd9Gpxqh65601uUHhTDhs6co6kfH
t7gjZezzof/9oPWKdL8EZBDHnXF8c1qNwKwfeK+15jo8bLTddXpZPY5n7MQEWLZoHR/2+BpZw/Dz
hiL/7/iFLCj6SrFyn6fuqwBQGV7oaafE58ZPvCj03ixCvwIWSrcAkKjAozbo7dALx74jDA92weYb
s5deveVqyV6l77RYdRVt6YmhmrCiXT9Av+ykYVPESp1ZBVcetW6p4YbRddQQ/6/fS8QlUvQy3iUi
d7X+igEkdZFDEmSZ+0A9Q+AtJ7oPifo5NYB8nLLgNr2I8LkTOj7/AFUkZ//GOhdfxQzIgqAxGk/+
bpviYttB/lWK66xTKkaXxwkvNcB/JPeTuVZdcVSeDEaA4n8lAAtcA6Nk+C4AO6MlfzWlzw4FmbtT
kGuIJb9BOzKz2POpqHGjAqbg8be5etrSWv3UrcUSmBxeGG7ZwW3DqfDvjhNYesopdFyW8eoFaGL4
Mq5cHzd/Gjh4qpJ9Q8PqgrIDqJ20V0u905F40QN0qQaVOaSO5zMAv9cYruXRcVv9pTuldXfhFAbu
cz6GW5xpdIpp0f7JIjcPP6kWDrkDex3tQZ2SAZLZAvtsprp3M6oX2nP/QOBnyRfVmCJK/W4+DYaK
QupmHh/3he99E2qhzVc/4jtx3zE8uCsbrzqDJiOUmi0glia5GX4MkCe09q0+CNBbCl13pHCiQDDd
yWgzA/QLmEAHhYPaZ0ZIZK2JmhptGCjDuB1YfLTsvFEeo+RSYjwD/0S43NkPPTck7rhQkSyIvzzX
dRnLI6X8bKNmHRSIUXVZUdKT6hMSYgV6BxwfnzAtZIVBS40RdalSqGhygeUGD/zbf5HJCsQVUpCM
LlhXeg/3ONfYK6r9iLxAvkODPvzyVHKVnXDZTNE5PSRSGqXvsFwyTHh8AK0rAX92ZboPENfXeke5
oVHZRQgncM564Ma+0ZFhBtma0xvhPw/havBU4NVXZ2PGvLJ6vACoEDsUDLmtJHgQNzJHZ0ZW+cX/
MLAXFf/aU5H9z8p+rmwYRaaKR+h518OO0/benJcmVZoetsgFk22/axhcEb4+GqyRTBpUlGOptGTK
06ly/RFY8eO34UQJbH9C6SyY4ZRLi/194nhkyv49b+yheGjMosXIsaNAVelh37QlX5mA4uqbMcbv
nMGt13lkcPBWPsimDcM3+r2x5wNKdBmyKETZcfrL2Y2JnZFx8PkCQxmb7n4vdY3yjg2yZJU11Sqn
Bw1G5U65czGPwZnZkuAeiadzwLrutvFE+jBbazmioh5C2iWjfbcFQbJ1z9XCCZ+9uasYey03wTwT
iRaH6F7hYVqog3IGhPjpxryMfAda82owbHbFkPZ1I+0ukpxtFclNgyAbfK4CEchczBVHDgrkK2ch
r3i8MTj8uW10hJgLwxDzn9Y0AFr+gl6F2fNONEXS0/YwMkAyDJwDZedywejGRiDQYtf455hTVCX2
7ELjPPjvMG/WdltGvNiP736Uu2olTNGwiC2vEScrcw+HFvb6gQOM4n04tkiol5QVKAxN6CyiQxOs
jTTRcONO8XZyNtHG+1opXgdAz29eh9NT5Si4M8pWcoUoEtXn8OKVwXangLpMjyyRrZNNZ2hf1lRZ
IijTVC7WBhmOkDtxaPBgkIMYWOiRpP61jtYU+VD1mnnUlWkV7ZS65tohP8TeydKPUtSS1K6LCQWj
+A6izdVMgMSMz5+iKBVYLIdlEAIChtmd8i6JuAS8JqNlaPE+EKZxL5/RzqnGzmIFNPi6ZgiR1dn6
wkIiolFM6sdE6uE3RBdhuv/JO3sb0/BZiLojaxJMVy7sM64N1Zo8ksaqKaqfWKgpBD2p/HwfQwU/
PJKNIqQdA8qB2db6IMt+Kc/qKShxzWjtWNtZMlMFfalrcOmZdkceif3Uc9z79Cb0sybcioYU+l+w
EZlBmuSSdrzhwJ5EmdiSv8QC1AdMN9S7VJK+n5C2VUuuolb1bhCfYiLQG8ELq1r9iIA1BY3yQy+/
Uz1Zpe95w376yM7lq65I/16it0lDMasEHQP53rDpFIlyuq7hPabgtKK6PKuuJ4HkLXDVZwA+Wttd
knsJonMpd2FocwF+bAE8BhbHPkgrPMJ/0EBD8CRIhhKhDPl2i0htN+rechj0A8eTjaRt0Ah3ONIE
oxxoVtlJr316WDyN0BnX9de3h6thzhUatipCynx9A9b18rWAEuUZ/F/CKF90/ZME5qceaYv9/4+k
EM6uc8Gav/4qTC/uOmOTYBogS6PbzYIEQmK5Q3ovtMs8/jB5GUVTeRL/DnjmRAZI83Th+U0anLFT
GHo2ABlvnZBGJR0ScaesbYAUzHMmA+x/ybpk0PhGxnnrFepAU57jh2BDKIbnlmuqMkj6MG+Kqml+
vbEOXu+O7IBqJfjZyGhV++/2B3DvSBVyo/EDDP1fFAgAY4nb+0RcosyEX4h5ZffBlhgwyWlyRuYH
rhzSNrDPOZmPzYjyhqCC5QKmUjNzKu9gCeaeAv6kq7QqFY5xpNzx0hfAS5DDdtH0dckTb7c/cVf7
j+iqAc5AyOL/L2Nj4bfIqANEjUpx4Pjbu298v6wxLLYYdfzt3NeQv0sPmS+gyC38LuOS6iG3T5uy
IFGzv+d85uEZxsR4Az1eHEFJEO5a3s6AK9dieEt8H5jhXxZIc9+SZTWFiXaFuZugaB1/llkaJ28u
PEJtXDK/aQLIrofb2LBa+MLFLYOQ0zNoUfF+vqwvdv8jjsOHFtP9H1ayjNZyt7xLpM9m8f3A4Eon
izZ84PXlVa0BWArBu13LOTi9Wl4zASqN7YwR/BmxxjhoeAqQK/+yKDefZusY0eppqh6AMv/b8wvZ
a13Sz+ZHhcINxPnt5kNjkPyWrfzGdnElWU7fn82ovpAgLXeyVOVn9F9N8f92XzEKYG53+MsCtqfM
6ckJlCMR4HbFup+EWlYcDUinMwE9Z2PFdS6+EQ54bMw5wbBF8ffJNUOeRt6FCYJj5YDZo8UBzNwV
DFVdvL3PcZAqL5Q2rALbvilUkl7Vwee6YiGiG1Ai/v8O+rU2e1wGXCqG6nYEshgmN1tu8LCyOTgJ
qyPZK3ZkOo85sxLoMTfXA59RiOb0+gnP8RzWBoexyEvjZ0LT58eChBcMaXNSRR/SF4DkeZx7eySN
UVBBVP6NUxN4YQ/IIlt+85ZdhHRSJsSE/RhjZI6YYPvP5TGYO2ongKo/yW577YNjiMOs7+SaYRX5
64YRIin7lM7x+bo6t9PRI6qq9o4nhndwYE1/MN3+4GVrW2ivXzMgVtWn5S5FtyNqlsPZMqEpJi5z
71LjtaLzD6Q6UAsSTruwc0TneD5LzdcbiWRsu4nlNEaOvIwAf2VOQxhTmrbMeEdMH1+RXZeHAny6
SvS7mv3IdqePraggh2zXcUx9FbBtLLQvrbFolvhfXCufx6yHH31sbwafUnlqUWLpSjCdgqT0CfxM
pTVETk0jQCxOgz2QRxZiXO3R4mviJCwnMtzf2osqfMIy+4pwEzf1BF4iXEQ0Ddx6W0j/m/73HFbR
W9+9XmgIts1PEPb5Q31+um9B0+0fnlZQJJOt0cniYNnr8XadGLKhbb/lCUyJ9ZT3QxuDfTnlk4OX
gKPLYLuxR6FXOuJrJkMFXR4rsSVUnTPK17Bn/KtkGI9molmUcvpKyx45o8sePZhbutP4CckKqsH+
vQjB+yjaAqSb1VsP+3BL0n3nzW10DDT7iBPSmqd0V1UBVL8QlNH3ZGsVU9g6SIaXpgDdavXUyEgv
OynTvEJ0Q6Mx1bSTlmiXbCwlX4bVPgJMWNCs/s0R86tyMRv7YwK4Rkh318K9vy2XdugosojoT9Yl
NrWA976cMaeK+BeA25dQpioMi9OuxRGTd7qIovcCBSMYWymOeEosSYI+ZRsiYOy+YPxxm2PQ4Aw9
AJxd3mpbLBFn8JsAa3dnMJW4TNUg0gIZvHlfGOFAJT3g/Ct4YVw/MEfekHCubTGgconhCV0TLRec
P7hae5+RWfPNm8ceS1ENZQ7a5tdOA3IME92YovBSa8VurjsALfvbpKs5qL6zxW2AQ8QBUc9OYMG3
G4GklwT6x26mM3PKZiH86hs6kNjY7rMMScB3tuvIx3z4oIhBZLUgIsDMM9fR5k0lSwp+d1Lp6zdB
wKc5SIfhUkrToJEKVVo2gZjgBr6yvnUD+0M+KLeA2Al/tQEhI6xWSIGEzba2wOxSBeA2ammQQm/g
NH/8eMEzhnJn8Bl9/F/rHOgmef60kBYFD1B2FUw61Lw/emE7RjeVYFB6GFHhRbcU633OaaR2Eaui
0Xkn8P1zCRrAHFtNhlmBH7eOxFJ2M9cAtonsp8RwWyUU+xrEox25dcI5SnK78x9S2NIef0PpLNe3
0ZnW+pfnJveOyWI2ABmRMQ6WlCAkBsN0w1uIpLecV6mOZCJpeVFJKNQTUMd07QFU/KLhGjt1JSF1
2V/q186ViZipWT4Y406aH3HalsPxKYMI6UY9bGOs7YBdgND0MncejMuQBX0I5GlXZ3kJjgW32DaH
AD55jKteY2m93b7UHv6Ng+DgOljaEMAi5jNUUnPXudZ+4uiH11753Azhs/Iv46lCVIx9Vicf3UO+
8NZAusUWfJRh7gqZhQutB9vSjZl0tVrh7Fgn2XyigeqbrJNNEj09xKQAVE3gian+QiKjc5VAgNqL
kO+upFPpyJfsqMPSortQk+ey8ELKpg22rODa8udisiLbOmvNfz7TI+rbCmt69VtdFbatbOhVJw13
MpLXV0zv7P6RdDrRq1QTsXC0ZQby9SBP4z2w2SNYb+WYE4FdDXM0kI/AyhcoAQ+2KX7vA3zTBItF
bfhEoiTDJfrX3VOyE2qXXYeSiDIvXA47FJQJYyeyg7z5aZlxoS8FvMVZAPs4lLeUKL6KhVa1ORCX
KL/6xzfAcomRTi0NDvQkXKvSOzpLbVNsEaLO4SOX9OVAOP7cxk1i6N+s3vN0EaWMD4Uc4AX9oFAF
a6VONlJc5Ks14LgL/ujvQSgKoIWVdEeeFWKIKd5/GvQquGj+EiOLjqMTqeJpb6GELo0PJmVSXqvf
88T1NoycCslFVvLsmpXL7ASIUPWnE+kxPt7b//LSLrEJRStjIDvJwVmULOb3Hf7laL6dvP+VDNR9
Uh4pfv1q6kEh5xWeknZI8JNMjc7Isr7TitvIA24v/TOSxOX6lF+sVOeEK5oAvtJ1098iglit2Tup
xyga0Dxvy23xMGL/HSvtWU0cHzBv6kOjTwQQnGk2fY7MdaUSKG1SJSz+7NVCuqa15S73guGJQfLB
7YLzIJ3oX0jAHOxla49ecS6YqQK3WFfa9qHjKG9ObSuUhJpCsobMV0D4IDFzHr+zy/FVmV4hP7W5
r4USindzeZOv8xy2xdsu0QqkbvIEaJE2fbo6WEeO3AeRjv51piSs6FGxgcMPxe2PBgq44zMyeHiZ
WAKVh5vIDx11EljOEChV7mL/OMGGWvFoKjMoHnfaGZjpG2vjX/NOfsAYAsHSfnUFq0teCpdVVj4V
dhjdiBA9baI2QAFXQsz35OrD3YHjqeNORPm4p7yNiKGzOq67I9nvn5/HYBpG4GIym9lyXH12zczN
oi9dgZP0LfzJybCeonJ0eeK0Hg5kpNtXPb9tLNOdPqW1VD6kCNALeVIKQD6/mxAEqFXTz8ad6ZaV
diTZg7zZrhWqgs/Nj2WyFh/+8Zw7GEU0CKYbzs6m30OcJ6MSQJSLvW6RWj8SpFPOHmhH377PA91q
C61AeaWssiuPUdERjNGK4xdLOW+bkp3t0+1boO3XGujdY+kiH8oiCht3HaLe53r6OmHXMUParNrr
+HQdyaI7LeGI9ML/o16vybpmaYxmRAT8QOlvuAO6eGm1XuB9jha26DfxeGIddnnCAOiK7cQ2HjH2
gguPEl0IzhQB/aG+riJtDI99QQTMV2NEq3aHjBmgxJUbq2h/SzCkxK3bGPH5uTarEQDYWvbRQhbv
fI9m5QRmdaTDiHz+A3TkXQ1QyPNVT1JqdDJiu7QooUHFfWluA8CNJpG/wbcjmGZHoQdeNx8kdKKO
kCBwI2uk2crHRLesb4H1Y5Xk7iqxXPi2Vlt5G2XDwdc3R80cN1jA0wWWjR2kGyE1ctYKzUj8fp3v
XpL6iLFq12O2jz46r6EPe4GOEm+XEjRwNupdFHKn80Quo15Cm13tnYFqUk7zNUCn+6d0ugJE1Sp6
PzEF2iUo1mpiOACxyktlReqg7g3eEikT3vZxkUPxVMnlJI70eO/wN4PIIYghEBFCx4T9Ru4hvzZ0
u6Ue4V1UQNJLS0Au0HyVSHA/WEPguBreqAN/rZ9nmGZE0qJ64PN5Ml1ovOrNCHnGPhmqqr2PJZY2
sgML+UlDfyKNLxKDsBtN2kFZJkwoSmPU7aEwb1G7MJp0U9ylvX9axmjzOSTRwVYuxUPrUC6dCpWR
ZHP15++vD4WYz+nehoxXEVpqO22naC+VdIxwwL2PvxXA0kvODRuOp+z5sP361URrOKVpJ5EjrFde
CPv5GMYQTj+DPPJJmSOd4B6VIkVjZYHia4cwK5RbeNb8zAaVvAkt616glVl7l2b2xrTZToNwN7Rq
YfNkIuKx9sXDXXuu3oQG8ht22+Yg5Duhu2JPjLfUnoPE51/k2zJ3HIzlbP95meFH05Aq3ocjZxMC
ybXyJcvWtd43W2JPyDy1VRLHeJ2CcYBDt8Z4nhbn4o5tGXkErVEchxegdkcX3hrFm2C5YDk1cxa5
HmNBx1GOXx7+MfiMYBrUG3uAjJXy2RD9UrUn5QJQDiQazUEJTUCDy2rTlSJC+mK32tkspgmVN2S0
/3Xzj0jAR4v8MeWLSOT+drp/CAO8dOl0ZehKW+XcS+IZycn7orfnEfaoSuW8T4u1k4yAXWkAY1di
nq9U3noHuHZ0lgSQb2LhY7FRmPTbDonu9FOM6YNevmm5D/HPEKhgB8eoLl/0P9VPAxk00XYzSMb9
ueVv/ZCBk+3WnveJVXByWMhj/LJvCZ1xLxmfw3yBGdfLgUHSoPHq2Vt+IU4So8CfuWCQjE13pgTY
rOlHkcfyqHeYm35FPCrXsxnsJ+y7OmsJDRTHeWOk+wFeOkXiwsb+1pNFldqlS8v15WBhocSiLI3+
5fCH1K78Z6uH91bHnlptsfk+ub3apja8YFisy2vLZGwNw0WHdzp1/fyf2+ayQvGowBs+dheY+ZWU
Y89qFSTYH/tx6znWX0X+HzV4lIgxb6NWOGdQ+We/+ruXxzQ4gSgpiRs9VXhDmeS0lL+8OTPldXp5
wLFtAuRrZCT5st6w3fItDbpJOwnhl2i6woyGSDsGOdWWs5mS+WEoBDcvK+Wt0letsnVF7y/kzW6b
fcfmb6yf0Dl/fzVS0efR+KCfhwYxvaqvDmJ+iQl4VjRcAGIylRTCqA/nziTqtC7jUMSgT6qVa1+0
08X2vwNsXC2wLy5LTer6jwjnfD6kuWkhY6c+W5McT96bJynLj1ov8JRF+ZnOrDwwH0NPQCZ/D8lb
Zow9LYylW+I3HK9TGbZLdFzCoZueVxyakNZsNyuThbDwOKwgQrgC7gkghg200d3G9fzyqNsJPrcF
1w8x+5CDs2UxXLRf1ZRz1vvq51JUVeKKbsbyyn7k5Fzm8Ji9wGXAU61eJh1PF+a4LIe2nN7pUqwZ
WYE62InBbNNirxH0f9v60HZAOOQMBURZChupNhBKo0lSY3fbLs+OGTJ9c5p+2jLTVfC4nwcd/kQt
nRbUz27KSkQrJjrC3I1P9EqlyHwR+STVVOt3caHHIaZ67leqL3q//paQxhVWLp2Nj4519EhgtfJy
29GqdIrxQRyFNgdbh32rCdgzfenzu9U0C4sWOHZ+ZdF7FCKYE4vho8FAwUeC6486S9PxV22OY7d+
baMn7YZ/j5cXwFdDzBgAj0ptoMU1XmUnq2oT19F0Xipfjsc2AmTRn4CeL+ADfxAJ4SKUhNOOsmni
jQPGKamKOl29fLmzwgoLbNYvNsAKFEYVhC5t8pLPaIcDruT6vp4dN9QICfYaGDvsWxX7YTh43rop
hEHzc2AWoJYIXP1cHhD55KQhpZdC7kE7MmI3pLMeZEnp3XkSUMW/t1CPN/KMMFZhls0tU3z2d5fK
sGSbQ4lmjvhyqZ8GzxKd5yth3eDjZFM6wKNAJQX51OhjVvq0VAqtNtrV8fOSpRPQNFsm+ScLrce6
AgFxZMVFu2iQ2jlPmk7Iz58wQ2J8N/4i1ZRCc6HLu9sTMHQBeVj+EcxWboDJQV0hN76Qlk9A5hTF
Lsa0jARvXLFziJy6wADdWKdusMIMe7me/r7Ajo252ifsRd+AmwPvo9rzA+Xaz42aiXPddze7EELM
7P6h4j0vfgc2ZXM9OrxpRwTmdNDUIqTvml9+dieQ6nm976mlaE92HBlTdYBq+Q56CrG4Xo1ik2Bn
/s46pDHG1kwaQgqOSpgSBPtdND9BKP51haUFshiJtzjxQrj2uJxdRfpbUDDbMfOaH/44d42H7CQx
36mAy/GKOXPDHrXcWLGgaBXL5UeBAJ2nmf8JpVwYOeDh7sBp4L1UYW8p/L62rpTpIMOHJg/iA++W
mL5gC94862Xfa3H4uqqRAihnfCbeDZY0Dx6rjrOt43Gux72PVWijf0aOuroV1pvosJX3qzPbYvTB
zml6C8bfUchcKL9FmrhUONqadnjckmnDmdk67kEY5GRc55mRmNsHcII7Iywl22XBVDdYoEbtyMBJ
wVQtAPVaPFOh2SxkH2GNbishPVcduMd3pVOiUoehRn/7EvDYlLdLDRB5UirFh2CVGhDm3pSXvEnR
zzq2Pii0NFoQynNNBbNvaRAUX2CUaGcq68gP9HxxZw+Wdr7B56TY07uese1Yw+ryrbv72godaUfP
T86bkd8nKiIkBo4vFVWoUYIgjWWvIESdvusuUQ2PtbXJ0CrvDnCvUUT8KGuu6CS4U2EkA2JH3DkT
9e4NV25Nk5yYDhD2drldI5mvY0wdz4526oekwyRDHbjGraW5ThreEOxcc749+9xn2685HMS1sjdk
8kK7dzsmcVDlWRJc5yZ1CdCx3FQ8/NdfBnuHDiF2j24JxdSofZt/9iXP6CHY0J1jq+ZnFe29h8L4
JHEkUJMv+Gx3GnJv6CS8Rdc7ilrHbhvUGXw5vSjJRR/9y0PwfgrvImiA9O0tsIoGPYvHCOmIrGzg
LUaTqZMc20afC4Wq7sruZnKgtWejx2TEzsxX6/a2kE6sr9WiRc/WkzWjkpmZIXu/+pYmRxO4m+No
nm5r70xSHgwsf0yG/t9t2oHFDxv4WVGDZ5KCl7tSHnPED6TnR1Y43tFGLM+I9nK8uZNumdQLVlL4
AYjT6rjJzxAX1EGSQLEpKyvwNv/LKFPwH/krrK05HoQfyOfllyEYPEuMAEFtcBOJdZNkXSzrp5lr
DeE0buYONkr7+WnWlBaZW/WrUaMNLWdHCe3RMc/Tt0c57wolRK29NQ62u0VXd6rvEgNaUITBdO+m
wd0Cs/PNZMscixnW3sKMuN37gjkbO5vX+iYDRKoB6Ntg/hQDiBRhxfW5jtMpifo1w7njgB+d4W0Y
AH3KgBNHS6xac5Z5gRRoUuZ3mR1X63A0UMYiMpTcfxhaACQH8OI4b3G0PPVauouiavYZKFNT5IIg
XczzPCnzxO+5ruRozt/UhhiWb/UdNWVmOmvPvMojGttXF3vsm4qDJjHVHZLiT3LTmNzOHj248Ybv
RT0ZabRxoR2yer4EVbjrxTWawCsLEh5v6qyYmotybHkqPcgYVc4J23bzVtAiUD9CuZtwwksn7j1i
jS5uabaK2BMmD7Y9OtOBHWv9cpuHs9QXUXzMT9C7etSel7U82hXUyEOCIKRlGPpPNaKgzSfIrT23
depQmn5I/dchm3IiySGAPHqEZiOXXrs4Jjj79BjVFElxS0W2w25P70++lJdq9E3IDOXY57MU+x1s
ylP7y6bbkWq4UfXNGC9V4pxBPCmmvg4A933LWWaq0QLpun/kseMt1Fp4rT7atGnKw9BaplqBrRmu
1+SGM1C/5kZ22jTcXLvglreFSCdxIrfbCzp4NIOpX1WRE4IdmLDlH7fvrYi1OJOnZdmognVg9IWa
yeWmbAWlZ/GjNVqZrOaAloG9Vhk1WHERyX97e6itG/fEku/DfssBC8avQQXL+C6DjexPla4srO8i
DEI7iwC6qDDBw/63juPri52jyoCRADMe1jF7RmNAWLNvh1XGzeRnhr5yqFMf0z9e/xuxuZGe4GX3
obV9sB84kMyV0F1e2VQJdoFNm/RJe69ZvrlFvCeiFnG70LdTVNxYkQCKFte1A2zzsyLrKsP7J9fi
LIYp5sTW6XvzMJPZB9Wi9WVOP5soYr98c991tfgpBe0qm2z3i7//oqydv32AqUUSvMLFfHSEkxba
2XU7HqBmjGcW0pIjXDXWdLZ27ONKz+HUNid3dx5BDpiRj31VyWIbjDuW2RwIOo8lLBtRCY9y7sj2
ltdYRAkCMLbmYsx1zwUjWrDzuwr3mkYXsISZUHPaKPJFR+zEah3fyoQcIMzGAOl+lFzSD23UmzC9
gBJ+LMdUrZYrhkncPGLYUFLMtatiQPKqJjxXz2DCNHtrbSJ2f4exaQ9dOrbZMgPR35K7adufar9V
Wp8ggEQjle3QY1USYCeHgLMICapUFPjzcSWD35dMMrcsIvT2etnHg/qaHp7zSdcJ3clcWOoS67yd
3gZMTyogGTH3gsKcA0sdr+f79ixKddeZhy63p1XAUrOgHRwcgj+cF/1fV9p752T70uUBgUXE55kI
d2wfUhJDDsClHPTb4ddzRoLilRqE/g8YLjElFCh6LqC89OPUq0O+cypEj2PAWW7gKZV8N+ac7xVv
57orIm7L1kF6VT/dIorWlANobFyrEOYhgT0RtbDZ/MX0amildXMc0rSi4AaOhKaJPeqapAFtpOpY
K2QZZas+fMxCXTmsztzALedpmxAPHtLR+wYsJJaV/2gwe2dVpHR3A1wkUu27a4KhMbdCruDIAZCZ
lGkcnZfpdCbNuGydRNjqaNGf/aihOlyRfacw0Zf1o1fjIWiJ+Ofl/KcU44xx2B8lR3osP5Aoammk
kS54mpmSIBIfhISD+6K0aJ5qnIDCSqqTETSd6YWJft1zLVjnnCQsVu1rZcKR3DN7uYRxy59nE6C4
IY/wQwyyJBPCPaJMngAlRmcO32lfge9FcJvV1Kb0KqRLVNLh2aczCju6xnVtNqebTkXVgaTq8A9a
TaiFeeVQNRsI5OEBaIgTX4x7RXVhBTXY6HGLnzZJ27KkWBXloXlyEVJQdqAbINoraWUMCARe9WlV
7NKxDrBhLY7An5A9WqL0lcMpWGtH3NHMdmxUp+Vi1W23dN71L67gWzE3mvviCEnZHYFgRxDSxTVC
WIcpaNKHuckjoMhUdHFaWEah9RJ1YOlJ9dKT65TYEQV5Q3f1en/koDVobRidHycK98OYOcUord4D
x1LNoJzS7d30y6V8lMomFbAwViZGD7Q1NGKtgnz9hEGnOBMsZEoCJojEVa3O4i9l5I5i8lYvzzlR
YgCgkhJx4HmIKHTJusozxIs1br6fxVprwsRCsSIPUc59ZzXp6DVjuMNqVLqB+YkTC2vJF+eYGcGP
wob5GtXCeYFYgXjim+Kl8F9y7T+EQTUp6Fez0q/j5gsC+1EIAu16kQ5XfmmDZ0fylKdXFHvRtgr9
6mQdasenR73WEulSbNZ/JSD7WobZJdnrPQjzHwXwBlUMxUJhWYzxpB4guP910vsiyZgb4JplxngM
ssfb42+hdE3MooUu6cpxECeZJbpugwW0om+wGLo0ILjqb/DO/sAbRRYqlICTX3cAnyvqgMG7elPI
vz8MIcrCKaL6D0pMVIw1ADUv7q8pG6k2KV6YzX6a3NzprVoi6awqxszuHkEgQb1T02cpGZAjUlZS
Co1+iuMmDUhyba2mVIHqof122mjSWhZUlujXK1afr+LumLmdHNpdk+gV5xMFegKtxp/bHHz7rMW4
6wNFFd5I0SNtyvQ4ZCtc4r5SCdiJnbtJgcDBnjJUH9lEL6gdwVBC+WacXGK2iEGkXDbpjgPPfqG7
h0l+/o98/yVrGwqvEYBThSaXp2R6xIvTXeGuVIXMQn8N6KTxDAgZ/cY+Gn99QvzALm3aYD1fF4X4
oS7A6IyTN9714MtvS5s2LXkCsoWvn5VQ8uk/Plkn5hmjn4lj9pXj/FSztvYVIwNVUZ5L9zjKJ8kv
01LIu4IAwl875mYnMcMwPhlPSdRDVdrVXlezY8Rcq0NOf5xwumvOnIAqbhVZN1LOutDX6RKXfcGI
rmDeiJzkZIjDvjVxnNAAWyAOLyn2k01hNFydXOmfP3MVjpdLzq5Zx6TFdy1lDfnlGd87E6vMBEPE
TdI6eJkLDy7QDhD167QJUb7TIb6+v3q0h6jB8/KJqytlB0meHdPN+JEBK8fQcbC2tXEoxA+rEGL/
kl8CExghqYDvLFMMV2AmiUp5NePxu7NEu2Bb4p2phl37RRvJ3JEoLwFL68lcHFkH/7/4gBBcUCJn
+O0dYDqp0N8OmM5pU5J57I0nteMyCqMNrqr2M4Mvpa3oy0MYDQc+Z8t64zSIohsm/YgtZzy1Sf1j
MHP4iNmqmVSuEH4Ost4KxikbZrOUFcdCx6LdVYknYBQs87Y6AebP4G2Lp2YbdjY41bPyFiw3jvBX
CCEnT48hHZb8P9VcurCadkFYPvA0BUPnasg6L90pH6+7EjIi1lfW/48EyIabhCaej0nijAy9DG9x
UPajbild6OkmuFfuoHdR1Otx6TgENuu8EspoBKMUpG/s8Kz8Ku9w6YnwGBHQ+Ys93zmDHglfx+Ii
AHtmPR4BarHjOW5AROhr0XfHfvDWN0F3KNoHRP+Yme0HsSleLjs+MBSarkjOFVt1PupENasElNdb
lzP21npCl2bduqiF/Oqv3K6UU7u0ykjpJCnV0PqIgUy2U9ElVdOW4s+iADdcmH/b4kMp+1HgPKKE
zvXsJZGTAc5zN7uHau/nvPjBBIyk7ELADxugROEvFXD9YkFDySnbmchFh6WwYKsY2wpYP7aDUI3T
aNA+lH+Hc0SP7JvvgEPisfqV4o5xd94oYhRFJ40GqCXyMCnCv+jq1Jjj4eJgtEDQm41uCLZI5XES
rtqDbbXSONoMXts3xHw4qH7DN7LeS3kAUw8CeY/u7h6ngc9CFbBBPtOXb2Q2rgQdRkhJpNOawPYI
MTAKD527eS2X/0XaK1KUEdVEgfzevKNnVZeVOkfDsmNsTa7DXkeTGafe0SbAmKw5WpQwOUWU0oeJ
NObswnjrIaYZpauCJ6cNv7CDHCSiJQ9eHhU43Af2BsKMAGQcbAzKhm86ovoXJMDEr3I/AfUb3HS0
g0ToLm0Aj8e+NJ8hLL5YCNgFUV2LhPBo1BDMPj2NAu/JkrYzuMsOUReH+W8DyiPBcDthnhBMgLS9
qnCvMifBD1U1cTxorFzfiza2Ux3eo2EIP71fO3lOCibyE6nWTIcn8ZC+LJrTsc6g7YjeyO2UvV3z
4BvIp7j64LZO8Ms9YKbBwm9Lv22oPxwyUiDaabROqqr4NzzPSkVtpdopoARVk+uqUQHbDNuO7K3j
s2/15qnxMjcaZC39XWZiLHaButDDyWMlFe5BjvmqtPHumH2S81/rjVSgqoh6Uk1S07wBu1R5sDsl
00gJGX+NyoAvMMgON1HLTTUlahvXynn0tzp+EgyZSPgayNzhVoISTYNwqEarAbsOwbF2GvY2dR3k
7k3JgCDBYaWLQpR43n6aid3ZXPmFwLAFUjRhMcGJGI3JWm9xDdVfrCtn4l0fel93dl68Zk/T1LSu
rEfVL9eNVB4NYU4cfJlIE402HK/pu//IsZ69LU1D/1MbwGrhDDhQCMYXiB0FvCjKsWb2XmwGkMnL
bIRtPtNSS8pmA+ilA4WqP09DBVfKZBrEJi0gpO3Hdydxx/qBn5FwK/oD3kUF48AoeNd0MqfFZTqr
p4L/70H6JXAtOYU/btRfB3lfNYGlB19P56ojA6MBFwdBaDjlMuL4ePX55w7bS/BJqfikysej/2Dc
qZC/UZXgwwheL+kh66DazJmhgBviAqPSwVA/FPSXa8QGOtVnVGEjdyxGpKeRu3lq8gOG1ixgv3YP
0u+PoCvRr526SlS1kUL98Ay4eXOPBv3Pu6lgVvrQdn89LF7wptiK8f0I82rfo+dpyHrasrrlV31X
4XWlWCwt6WieXBH1W85NmKEnum7+BxKAICFc3/HFpsQSa3jSTa//3Uqdnk8q5msgjK2KnKsziA0W
Q20qGwWvOCfohKhkJAOeUZ5ny2denilnzIlcuyMqgzM3Mo36zBqI2wJvXmnRKeraI0toKh8w1kWL
t9ZFVq0Qftye2OBaMVYJDsmwc77lS7ZAYLbdvYSAAz/rAP1RIoZxF5eBf1lJmyF0/dNGO+hGj2+E
5geWhNiAscdXPnq0crMXYV9LOLECzSJ/9lO2gFkX7OkqUxyXr412zhfO/NELfFIKHppetzFNo7WV
2op1BQ9f8z7XNorg0eyhW4yInSzcqICMDAVX48iQqp+ULpaiiRYZZbtZjTSXwhJvBfYYIjngf2BT
CNR16pFB75ELlbOND1E1bmwVnuO6JBJV9Fse6j1NKbwZfMflNkkf9nz5tVNXhW4dXp89lh774/8F
PWvgZAI9sNhHXHKKPks0nt10fNYINdrHi+Q6ciB86P+LZbm5lwshuXmcGoulcmE+gX+fns/pXbvi
b3KJzvJwsSR06UVScs1/XbNYbfQFszOSIgGg8vTt1udP+amiXuCs7rd4DBa8xUSQDU3SZqQDmqsm
s7jrHvZz1Z618Sn5I4Urf0C37QlXKT8zfM/tx+FoQoaRVCc+y3wE9/V8oBmZjkOWbOZfwvI1pIoo
kNx7qEXxt9RYNG+t+P6xAD8QkhUuCTfcjlK23KFxa57c4OTvWrUKIY4kcnWYBBaaPc0kE0pBKRLI
lcNAVDzjJGlqO9LGviOryzRfg/OK3/R4XrokZeF5gCkN7QwMenEckK2cK9aT77TAAYL2pSKWkJkr
LQOFDuURNcoQUfdN+pd051119ohsNJdDUhlBtRb3lqivNkyNVBng8t6KrU7M2ZqpQOVojVfskLF2
8+gX2nptsZViuBJARkWoi70MPc88A1aMnasdhtD3tpyIFOKC+97R0KygOCET9+sOgJOpxSLEZpOj
LJAKhiU5IpPtgaz2oTc6c8g08zjGPlZCkWBu3uwZr7squhsB6cICGbuPHCPSm15OMR2fD4/BqXZi
aTKQzDhvRAUpnvjbaSnYtXshxbMcYiD+Ix0YwuGE4trsVfFvNqOPnXr6MbVKORb+6DqOfmQAbRgt
vHtZZoKwyo/nnnoh+4ufOYCrT2EAC7Rwyl2V1OlRTJqDkgwqv9Tk9iWV/6i3ZuJBqRuDBSRKEfjO
FIt7nT/HLuIOGlDXF+Hc7oUwQv+Yo/kie3Q8AtBhdpqZ+OyJE7Xma+o4+i2L23Oq/VuPSfwjUVqx
I2AIBVy+tQ6GzUz8sQ9my+9AmNMPpJ4basVCTrSIroGQqT8wpsWy1jDbQ3eDzVaQPFary3DhH7iP
JuvVWONjXV3x3znMyzTTxoPTx011hx5meK5vv2R86nw02gLLNkIaPou/cwcEvT4TdXDTLmQ6b5WA
p4r2urZMmGLgoVGNB7R6B/pnTEBTLbm2dQjikSUkshp1lZRarF8oHv0anPVpRIZie4GmWqIjnSvq
KbmiFdmKhV09EhVuvuHhEuByGPDAfjWIayqzipBJs606Qeo7nOJcexbinqnw12XNm7gT+YbA3NuD
BiHj5QIHRg2QocH7dfJcG0hDzFCNWXaG+Ljf659GWCQbkZLzK3IH999YFAgmsFJkxgXE7WIlod8W
7tKsN0pJZuo4AsKZV36xcef36Zx2sp0dLvtTO+cEcVKtQ/GV9ttXpdAp8yPyEHxA9wKy3EU+aZwd
tNaULtY09+ZYNi6OcSIFlR1FevACloJsmERE+dgriMB4CvccL7DVxjO9sGBDvMN4wpraPxEVDiAc
VWY1yU/sMRyKH1Fbz1/fmXZzq6dYOwNB9citRl2vraNLl+RKbUyrK1vxh+dATn5ZUevNIwWWjp37
M9UowPJ4z+CqddN7cE1AQ1OYYcuBaIk7WxQPIgDl6O960MnbZ0YBlsAPCBxom2DJrG7M9PnmvLGh
YKH9GxhFG4ylcT0+0ZIi5WQCj6Gwo35qNdx17w4RlDfc5lDfSup33sh8inK73KtEqyG2EiJh9Rt3
9kao1en+i9d/wieGlJPtoOkDe8NbwQd02h6A0E5mGa4SmX7RWka3OKgjUolvKioDG+L3axDiZ+Lv
eQu87BgpJrInyEJmCLu1bsg65hZ0hcuagLn0zh9TKzENLklubSYMUupH4GO0AuvBHeJHf5cg7txI
4tXn/J2z8s1gnCMJjQOMked2QcYqnhLnmF+aDCTSW5Flf0zIcFJfH1fJ9Y2odmaS8YXFtN3iEI2C
GCSwljT1JKs/Q6eeSnmDet4btFyWpF9g+nhhtEeFfUa+zsBhveYCqDCPMHk6/po7nzOjCdXL2KY6
byIQ1QqxpXRQp4W0/sVdUh4pA0m+PsXj96HOWhLEnV2OqmhEx4ymzvyWc/8pmtAZ/TNGVWwzbg52
g4/ZS+eqxKeRYjWebeh3vl1clUX+LbA8pejJ5ocxQzmZYwG4p4a7da3zZf8dH2SlKeD681vMQPpC
7NWJ0pwdlc+vvsuIyhDL0nzZK8U72XwgCRZDLie0XR14/sW9es2kPI5HOc6W1+syMGrbgd6s691D
TrRm+rVGZfzFkm8L2MyYhH/AxEOvwCN9HXG36WxkLX7ZsRkcD2kCeR09Ctp5PO/2AK4NYuln+ku4
b2IKGXwJdnK/gENPy0bgegZ/v1rl0sflAIzNLKeFmnXjPLh6VSiIU3pRg6VIk2J5hJsRnLTqQ11M
93igj1Sfz+hdqckOWqxQRPciVQCPaJHeA+lDOXgiR4H0n5PrUlr2GJxqoKa0e709kj0X+SrHBMVO
ilVe0kTDIYbDDGsD+RHj7Wfcwe3p+Zl9XtWtgTwFC6btHNuNf8yw2TOZZ+bD9Rr5kUkGxm4CE4LJ
LXysdKN3Qw/JzLuACivxaQWmYro0l1c6fKkF2iyorrmMfOqAVAJQL5kmdKyA+ZIxu24Kw+nzE3pI
zBeCVTVnAEeScoG3/C8BXSv843CdPFEu7Ag63x9X1JN5dQ4iL6VpvAYHeRh04mEzqVpSAaaGhAIs
NQf0eUWNphjPCOL6tx6iLeq+HhfnUKHQraCQniJc/F73v3cqoBgv2cjzn7JJWtiqVyasPc4ObmvH
a91oz3UrdlOHHTsCF08JYlpPxJQfe09JYyrvG5yp3vDOdf8pt1+7dc2PbXO4ZxRUdgir3W0DpoqQ
O+EYDUr+yv7tgodM+rxIeIV15TwsCBxfrGqgZvOsQHa4BkL6lttFHMxjqWrCLinCu/lx4KrT+7wo
r6tLNsAxFsH0YSS8mTBBGxlQI/y45YjO/SpMbw9/JaZx/H/MBnDWKecUIUEydDtE6k4Yp5yCqNXQ
K8sYnVt4TvC4T7bsGtNtOqi6rVZfzdW5WsHwG3Nki1PeMNJ25p20IQ5OGd9nGmZiAIWpL2xmndTb
iRgOeNCJODf5OsHi1K+q27kufqt8rVPCZBVDmpXQZNlcyaBH72F4vKl5WW3qyupUv0eZH4LxVEzd
T04KRi2U226f9NcARd4yPh15kwLfuV6wpJ4eqKGkbDgXlaFZozqdNZbvh79TUrNokkz2LAJlI+T4
CNByXFz3gGZ7f3M2YQarCSelimdHpVzUMSx4SDD1m5WWgxjJblgBUq7CepvLJaK+C3J1k7xH5KJ4
pClcKN7Wl/T9setGGEDdTY83NmTjRG0sm+J2bF8cg8POaLnn96OxZOKpG8satRvKf3RCvqbnYWKw
GI823DstR9Zn2dwNl/oULOB01Pc6I76R4p+zhnxITTcxlVHKompB7R33jWwDYr5e4m+8bc6nWkL2
qqMEk5dL7NUvsgtZYfXWkVHSHuxMF7+fxAlsBKS2aItiF7J0Q2eYDM5ktxXzGhmw9RRUVz7wgzmv
Zld8qdpzYvqVwZqLjcV5MHtwpF4V+4AvCrnElXnQMcxG17sJYjxmtkj9VrHoN+fPTiCg3Q0Vo/YU
HHPzjlIRoG/0w96CXKk+JN2TMd53S4W0lDIngQlwgM2DSwrT4odfhJeHiqWGMieRDxefT3CWkPV+
Hcv6YTR6JpvUtQyMnVz4AsSPEpjd85C75jTeAfWfVZLRWcDEiO4nPB7pH0zXjNd55MQsDL7fXxKr
rpHp2quqCNyu6rgLfucGe4bmLGau/5xdiZon7rOJgwdYq8/2nDortiMLn+8Y9HH8NWgl+ht6e/2T
mRMGsnLg53Xa1EjrZIKM7JHqRUzfxTccl1UbllQDc3qVULWfOyn9Q5JUyGVSXOVNJpgarrAcfbCi
5VFtb3FHkZKew5eJ/uBfQz+JFOLq/55mvOlYpGXLmZXWjCeyDdPpgXK3m1eFqtVuzT/LWT3J5cif
nwwQSswodIIxR/OkG07R03sq1fi/poSwlFnxMmeaA5XLoT7hmrEA11WdtbmcCF8c/vYruahj7BU7
Zuhl88/6FlYbyTAPYvzACNndDiIoJ2D+rSO3KanrH4D8qyQD/UBngskEVXQkBxDyg+tuP7sRgyYX
6reBXivgpD9Syfx2q6f7gG3Qq38t/US/XG8dDAIpJ7VMugLb27fGvBSCoo3BUAL1vryaC0HpIBJg
1Gq9Xqgo80uRoCKJrflkmfanV/d1HU9I2HckASv+5PbYL4eGJmJrzksDY0JmWL+nOUTzxOBHfFIe
/X8OPTBnM7J8PoA4+sL7WT58Dqi72NADKQ9ZpaKY2DFmygSp6DDjhtFBV/JmHSBa6T7R79+FMIky
SEsfJr3wT8817qanxRa8h7w2vIASw0NumgbZboTAQTDakBxMMVM5glotcPh6izokaAR/uJnFXWj3
A/xGDqJLL+cVNigNoQ+E32XrJ5kjHj1jJooH1cDn/tKhhaEamFyzVdIhOFk1OEi/ImA85TNd8vhC
MOsU8MkZ4k+pf5EEDjZZEtVm+yC1KZSTWPjgbjSys39Otg3C5Tm5/zSOrcMMfm2n/EYReoSuMOKJ
i8LI2HVzm0XcTL6dsuNY39IH8nz/ixdLdK4/DavHiFJ8YNLChOxLs/fEXClbIrVlE99Ha6y+UnPM
Q94R4CgXejtwxkBPOuz96bIwMvrmg6S1wZQA6H+7m5z5sBlxX8bCIJAVDwcAmXCvGFevjhZ/5Kg2
r61EfuCLTqoao8HTI+ycW0ku/DvjoKP5LVMVueQ+nVmjssSfuv1+PSlKofPmbpmusNI7CUAwShbS
sCcqxm1Sr71MQqs29dc+JGGPgeQt24C8fELTi4yOL5wkGg6mgkPwP1mQM/h57po44/FuRvtYUfM9
o0VlJG9i9Y8dCYZn1DR6ye/faWPzkKPw8ZYOUv6tjFdyxP7M81xlZVVpVxHDsZENlKwRti9/IBA+
kqkKYpySzQm9qXEE6xSVb5j07F3PaGpkEjz+aw5fbCKeWTVsitf84+XOHXfOJN/A8AfkOBDWPImh
9dRRwya6o8VahOg5M8pJ/0x3xesdJP6WLVwpnjk9LbK4WP2iBs8qV0YhQWV8nCH3FZkO97RSEDYN
UKEtyr3fM3MzB2FttxXSawfwW00pmTJXZUvS9C4RHO4Wys3JkO9j3PVZYQgOGUQU7KYW0eW9OBKJ
kel+EuNhXT6u0SgaObAAMNpFih/CAFhkui4sXk+oc0wvl6fLvEasp+E0ODZRzRcQ4gl0+mvImddM
M0Be5YK3C+PMrwaiwGJ0weSkKbvMdqz90bOdCp1gONb/ie5xUicOCzzxuspk7psLrd13BQPcaTGs
pSKTiCkhu+okD60w5ClFlLyychLSv7Z9XnSObJOCu5yJTgCGZ4D/CvVrrOiJ9po/poEN44MjhjP4
9LRCOlwvsPiTIMFZnn+Z7PCYuhVIXn5YTHBqWidKSPcPhKqh3uKDSXiKtJcEVn8DF1s0xpXrKcFv
hNk+8K+eRWZwGkM6kVXK0sXXImoxbaSIZyxzo/eE2oaG/RSztjxDkInqsc8SqLspyfVHUUwRCihD
q5zr335ojwtawFnGnj5rJzqC66A6PTbr0mwrwIfNKhd5c8NemJNDb+gpCOmlwrAitnygNVV7k7cY
3w++m37Ime3d/sodNVhkYN/Lsln01fnGyPHKxwLTn2M8AC6O4vsY6bG1uWVnO3YuBZG+MLJcFb+0
AgbZ1Mqds1rgEILODK60uB041Mx9xv8CRjahnM0yfTsUSWzj2eDLBG9VHNv5glpP299VHPyAK2MD
GLiH1rjPdGNxptjmMfZbPTmHFBCz1dpDh8Z+4fMcZudoEEtiiu27o9Dmz+yihlhm1QKng0jiTqO6
4MwQV9JeRGdtmNT3wc4DB3FxnlQU+dcjg7YPPw8EmAO/kc0T03uq5CdTjaTuCj3KNl/KTtJVlzcz
I4WO5z1kVcheGNfIJ0GcLSRUCZXc7mB1Gka1UPI8MEayCk/D69MzgPMJ56fXQYYNmvDhTG+dd1fz
sgbi5pmVfSwqO8UlS/MjJpYR5Qt80danC1nEAOK6HxRFudR8RZJ+1qvmNk1TclZVNgm6Fea8Ci+m
hgpYR9vOiokjgJMyPVuNEQV4dgCtkDG6WZvVcLRUjnc07YGA3hUpb1b8tWAThJ4KLZtQPioRHCsG
pSXtj5KYcfdivJrwbnqA2iRLtF0axLv+KCH0bD2MuEEaPybcFjC41AmnJ3v2mSfneYyc9ptAH7Un
7DXurYfIB0oNe1TIo9WPbVGYqEYgx/SDWb0d3kDi69VenI/0xUfiHcvFcTLytPulcFPUiJMCuXn8
tWndU+YaEcGbj4OWfEqT4yCfbrl1ZHoMxn363SgKHsgpBKLRBMsDC0C322zj/jWFrUNVc6vcuEJS
S1+6TAaxs6bbc66KoyPk2dTzj2C8aO7hOnIv4/AEIZ0OKJsRpz5GMZFGYAO92baqa8cqS0xP3HBt
6rdOG8YAyLA/54oF3oeO6y/vwT/cqVoPvxjmB4tv6E+Y5nvPtLNnlZPLt4bwaOV3v8whZAcjKJkX
sVi8bSxTLEvVL3SeXKxGlsTnLwu+FF2DohSS1d1yZzpPbfjxt4WjThyr8ebg09AZTqOYgvjsG2nH
Y2NgQ6bFB/uB2F5+16E5O3tKbFJyddDW0dlpVrFK+jKUmTNhxVYQ9pOx5l2sXMRdH0nmjmDMnNXr
atBh2mb7zpuXU7M1aD3L+kNXxHwdiOoptYM2NjMCAv3XS+knIwVAUbPzjEMNvMhbMOSBFx5Gr5hE
RXkS9CxG9FAvKOQvX1A/sX2VIInDpmK+O1i3ia1u84VEzQAQxEShjtDhpQQ3Tds0BZrzjQ9wzzYR
mNVAa8PXjAkvcOlnHZ7RavfBWMD9imTEThRnPkfn+384+vtvvKHtgmEFqFoFYPvkVPHTvO6D+EHf
JCFcx/qvVk+L2d4YMF/9dYhvqwLJbSQk5VT8ws+DI+TuVfuDC3/bPOZLtMorPI+HNZ+VWrsqL54q
nL+RgluYJdbO1Z6mbgbBaGZRa7UAWgQ7rvHx/1KQq6FpUh023Ab+HcOW6YSncCaCGaBXUDixFIqx
JCZLAGr85kDtykrCK5N2HBUtClIMWxS1PzWTtmzVKzNy/FwUkdbLdR6jHrbc1Ev9mlaTBk7/dLzG
A+I98O+jlySfkRzwxS21sZYF71OiRWYMKK/WxdqMIEQN+5ketkVfMDq+7pdT9MHcPGG4KaGQvDRX
gyEZJXAt/kQsRWsuFICqrg+F6p0Anocv3H2sh/RMZv9BrhPMuQrjfIkdxvl57prc78qXmsurLnuO
Kg2qRyLdmVD/zKQp/ue7+SkieZLX98b8MYKVseqgojHavEcLX9mV135T45wxG4LUpUsahxh+h8iC
aB3OHR/d8EERJeZnGJQnJcKbV5v054MmznwQRaE9BKRCZGSAjfdx3bDZIR8e/WCeLUUKCpx0k3iN
Q+Gy8O1kgqkLOF2JJovPPjSkkHakhR7OIEgTtNlsQ7FtK3ZwQOalCT/cgJzIL6qpula44e4+gqvU
rN5fBA0ReSfAr0c/YWhe4Ej6QD0cmOl5vrlh/NS+s8lEdKD0+uZgvDWmrcrZW1Bb2Z0+rO5jUFlO
x1S6SUS8gJxWBL6T0YZUbi0ATtjnHXs+P9VcE9jIpfHixm4RPS+H/hGAiYfoSz1BFK1aw+YMuhGA
T8dr+g5wqlxfA6KulMnvx10kgL7bDM5uE/M8svH6Xr1b7hBUmFM6aTadNKh8p6g0KLdHEURbjwWl
bOE86dZ2oEnqx0KbQ6yWnFmpBD9O9vPX150TrMckPg3ygQ/iYzk+RZZfxTDKjZU51g6Vs1xKzJNs
wubwBJgF4YF6DmZbmenMLa8QQ9Ve9pOnbD2Q5jJICjiUsuNnrQcHKC4wS1FltYtY3GNa6/rJLawO
XuWxeqJi6ExV475xYlVFWXw2FTz0+gLP6C3GAMOboiGcYD7ygr8oxn+EU/VT66T2adnLz1/Xg/tQ
NHqMvVN/fBNSJWD2cdT0JzeDx3HaSi+ts9i4/kNNqh+KeXp8Zd6hHUQXEQSweEZcAu2Mc4U27TW4
5t47t7hhObePbVP1Bl5QzkljsgwNGfccmrMX0dM2AMAKzR4sAdVvXwNOulSYtTeYmE+ClWGbqX3t
da4MneziUY67jk/X1fEpsT5NoQXNAoJV8U2Y/3x/s2deJg9FUkkiyni3mVEyrtd/YsJnuq/eoCo6
UYqVJCt8+L6JOhtVjfZrntBVFyuvjzpP3FhIQTiDQmFn1voja872UcOjE3XogOjHI2FKQ4ZYB8c3
aFA20KQRomurqNw59YMjhOzJ1OAXOA0OWxKdiydDOFWM8M5WMyy0VR+0ts0sduANbMtwfPBK0kqm
vqU7HO6haNMAcQ4kzhwy4GGRbdOL8pAmUoCiPiymMUpta40O12jUBEij0znBCInNp1lNvHlRSxl4
cyvA9iBJwgaHsz5SD6wdtInMQPXUDHHaINEV62IXOwvbITs98vIX97iuCdi/GXjfP/6uw0wFMo05
gMwUu2zcB4cxpx2P93AWTwT6aYtUKBA70rklZHDABNnPBEBzKz8ViXMuLf2bH2HNXpLc4hMSDWP3
Uyao+FodbH7yJ1f+1lEX25hoMC1TeliQuMLs4gWTvOG8heNhdv6RUqhC3ezI4G9Iu+ebKJJzSQdb
gTRxqlttT77aPxxsNV1h58Lqjzq29RqFM681dSE3x+S78pLuFX2p9eqt3CISlFxGNptcs+XGW48U
IY7wWuKKq/+UIgh9VmPp9gC85lMQlcM26nParSSGz1fGqRQy6mKr2fAqaIJUbzMW8LrpD/zKtOhD
3ZnLpj644T82yoa0sx/KiO1jZcNun0gCE4lXzqS9y0V9QZaoWLOobROTJR85XPo7TFFuTwUo5aHp
yz+dH3IvzYya6hDOu74MsFFhaOef4ehoJ/ZpnBHpd/oio6duPcjMsHCvt9H1nooy6Q814PeHe7Sm
y83Jm+ml5XGpG01KsNYHQTYpjTumMMRt9jbGl4r9bZlaiCEiZSSHwhYymjN5RM5jD1gaZARB+dSP
i8oHqsjEHwRRnlHWxXzYFs9H0jpqZVbFkh++mYoIk23eO/xtkJB5gToPVudQaIWFyUP4pWezikxt
jfO56Srvg+t+P1ByLyISugGBL4qMduCL882fs+sb8KB7A04Y5RsXoxwr5r0GT/Ddtmt7UwL1W1vU
3aFckJTUz4uKtANX/OpAE8fXTA534kfK9rE6dM599x0BQjX1O5t2pjq139NT7xEYLyjRNpe+cmjj
Sd+IMEDgajEbzKJiT7jPVf51NuCVuBh4D0Xx6jODqQI7fk1wIn4ZE2WMw9tBYnx3CLo1kSQXrszd
fzPlT3S8XLsHnBc5Q199xVr+Gi0zECxJreYEmEgAcrssOwSbVvx8twS/2Q2RcWv7wl/S7iKx9Ndt
jiYMmZYgv6xoWKDpu69QDSCAMOfoHjD1hGIBcpWyV97Wlw/fsxskjuJco5jZwarikN/289+zqEA+
zWrrjS4Y1Y0M2C6rm1i9fk3fUSTykTvcsX6OFnyWgejkPbP5tgfb+qyNAhAEtuaBW/Pp/4Bslodp
yQYwdHAALlsRlM5Tc5b8ivI/x8leG18Z7R/cT51kCFHZB+eQNXaRntGXWSxfcH5kaE7IUMrJ/WmO
a+0sw1qpCriRSy1bHPqmdmVzyaNB27NAoqORP/czBitGnWja912m75YVqMT861MAY9sTyznaI4tG
hjpv+0QP/YVGfhO/uTUXhp3CWKfsoDWZJyGV5oak6wPOjW3lmcSeUEcBhf10nMX3DTKBeN7HgsB6
s4Vc2atStjr17w7eNRk7rWIyvk/BSm0329zYCfOjtDakWNwWSuOLiKXPU+IAasNp6VOA44nnPgb/
5k8GH9JjWZPK4+DJsCkJMTuRZJX7SU6socTqdQ+m89jRVPP4AvnE6H2o7GIjkDingVmwjCZdJFu4
RTkeR+3mli8EoDlrEJAjx+6ZY08cGADXgrwGF+BYabc0kiP3DiooSFZK8Z/P/Aqc6VaUAEUuk2jX
pwwxjTW22ghcTzy/aD8SR2dERjD3kuNkp+cJUkWZ5i7qRS81qIBB9ak6BsJxpb4ataLGSWKMflKv
n9mGTZj4+b2wWG6tvdKrnvD5iI5xGoMqZJW1Gk9SJEXMUFH1JDGFbM41Rub8agyShWFM2oEzuofe
kZFuhQ9yoJSspWOW3ms0s65bo5kH3DeSTpkGnsVXXfHeTAjGjT2EA8i5x7i/sHwZ0YvXFLp8tVgz
Hk/vionU7iIpiwvoIr1e6ZYLuQ/IQI4YefWJAxKgjq2KSyd8fq4VgiJrRP7NG4CPJ4nKafSCY/9A
IhpzAKDNlWENKYDUzpKqwR6jSSx2BBChpE8EVj9Dus8ErTUuslGYcuUaUaQzY5l1caxyCzWjSaRR
jpsb4M3tjCFxF6aOzAq1ymPiKtoOD+h4ZN3zKDCOOLdmcEpRjWWGNuS9ezH4XjtUoH2BDMnF2l5h
6nQAIIyu1QCNZXl72vuQFLwQUPjP+xVomAbLCY8+GlUl6aBn3Dg04xTtTBekZ/jAwJBSjahdRtuX
7j2+GDWB23cHqbXpeLhFiggDr6wnceEZqc3SLL3ZSbTvKfJTrnz2u+UkIMHfbfIEzWg1+akuCGLV
Xey31at7CL+VDWytoB2Ho1tFjmQb8C+xZ0XMxQd2JqKKDiVPD4B0RaDLncJum5N7mfeKgjL4yrMS
bg7y95Jn44GkHvSOsuTRIvY+OGWG9Iuki8joEGu3droZXuCqM+xOm6W5HmebxTTylKjIJA20F2eg
BTQwI0WiPWYejF8thXv+mIXQZe5iUmGYx47fL0AWWba0vkCRUSnxkKHhD3FtPdfrFvvS4npdC5iO
rN/pEJVKPaK0aGrJFBlPfkNiEosj6yywzzmiPxH9Aj8LcH477eqAwXtJXM3I8lUykGugT9nQwYSh
GIMGVLpSLnCRBthpVvLAhsALKYJUJ6JHFbO3AJDIY1QGXs5h6o96vuXepkyPJs0hvU0DvL9mnRNG
R+cgU8px6KejPQ5xwnHjV4yiOrPTweSBrVXqLGJ6uGOk2/XFcg5DSj+sk5b5DCY5GevWbU5UtKdv
RNkJKlkI0wqIiwDD4hqV6ueB92ukW371J1rPHIMeNzadD0LTcurOIgmqxJLX6bE3aLCpNAXX7oY1
LFnjga2ixX6QsJ0rZeGOXD1qM7EN9kA2c+gQMVt4i5sa3jYIaJptZVkUsv7E79+cNsofA8q+Yktr
ZNWxkJESqp7ePM9TpLa7paX3IJRzZePdhf9VviB7PwQJoNNEFxfE65gI9SnVMZZTttFwJiE3Ii3f
ECUcMfHVPQcXciaY5LuSWe3VUSYvyP9NsV3eyEVPOa50v4ECozAYet+B3CfeYzg7jB7+GrEhCsFa
782FDWOG8od5vn6fTOZsjh9kzgRGl805dhjepUJtnx+snSjbIfMjMCKWBvAK0jW5xugmFJ6Mz4/x
GGeewM6PciJ7U3BcnIDjiu0N4Ndil0Wq92N7o/RC7F1/YW7u0JnqJovvfFgrV2xVLw5hriFeXRMQ
i4WAsrf65clp6tsVYOnV2hlCzXWghXQ3050K69uW3ILY3tQPktr9Q2VMUTVSk9061wVtQOJtGU2g
niJrk6BF7rOtV1FC9bdZh6G3rgf1340lS1T8wc4MSgZFG99SeiGNbLZj3uvAxapfeYHxQNxFblYe
YFnrpI440dWv9K6guH3grBHkeVDOPmQhErI2AkxYpNfVBEZaDQd4nFRj/F4ugtGJI3o58p3oKo2B
ZCyZhNewo3Q8BYpOUota6MVnhdwsWYgxTTWM8lAixo9hxRxt0rDBwu9ckEkj9XAtPFFXSp2rzcVl
GQCWUnM4hPNzdq9OMRRTeH+W42/uyX4MSl2cc1uFVphHnHcIUJhHk4adkP0AfmPPhkja61GiokKG
CSPbqvHGQYYznXSUJ1cDAf8O6pVdEI72KOelsXk/l0rWRaQmRjqVjvF5dQWZaAB/554XHvY/fYcu
DoICZ38Be9j+ne9gbr2FIFjtBm1F5jphic+5K2Fc+jlj5XT6LyUYug5u8ghDRQcmv3tGRoa/fnDn
VNjEDVH7BVgE0IYUCuAt8mi35jHvwkhWwd3RUvyemQR3t+WoIkz2HbVVDJx2q876ybpwdj9sTN9P
kcqiclWQjeBl5FRoGEj8qNYsY/SmltafBi90SzDOhcxO11yoOtO+DqLsE6x7eATEwWDiWGI0uX6X
uc75NZpwyC24psV/ssPkPmVVr1wYzPDLnABg/qa9i91BowL56GxCTogR2Wut/joaT5u5LHJ6d9sS
NyqY24Rjhxw+QVY8ysfZU+vgKYNiTNld9qFLWvL95o6EvcjnCAiVh+Indn25Y//MEYq0YW9ZQTnd
M/HOJQ8mySZSuq1HYomU7fVK5jYlpMKeaGqMg6cFgz4f/MHiB0X0BnteMc8Cj4W9PabVGcwh6hSM
zn4OHj13rlmPw2OD1lI4CaEJI6ESQw72ecl1uOzW7wsDdv3CT7JXmLWC8Bw2FYPgqp0I1ybgeeQP
FqSzXYVtiPV2vFwMtafKxpG55idXrjgeSfBkGv4QP1Z21la5QnIWeH55qJVPlDSXKewKeBRAmbmB
wlvohth1FdapHDnots8Lgwyr7wjc139Q3gRrosaWIPxwwb9j5ypQCA/aCIHFodJK9+gm45y2H2Vo
yzMqTk5gRnqIMlJcEoshTuNPnXWd0k2fsm+NVyTACoWdiqFQAuajGpY1vfLQWSV7XwzSVzrT3ZX3
OUOePe3asq5FMuQXC3naaexdt6c20Je7zLjEcNZWZKHWHSuv9oD1evGxOpqoJWUG4AN3xXv2H++1
H5ivwPPtG3mpt5iVr8/oqG4GML8oNFLgf/wDxuZGxdEFx8dzhxdZDXEJRRjm9KxAyFLpULWjA8f9
VIYhxPrfUEVkNXJXEFJwyG7Fi69TOTHCqKb6hzNpFd2N1pQU24AZYOclTySvCNBC1//nMHz0kMPg
HbqoxJzg4WYaLUPTYa/K/ynSy4MQEbrkaXxoxS64rdiFm0e2haWuaonspntApsHXG/OMDAIv+lN2
p5EhCl3ltP5wUWr96RLSA9EyrlQdpyb09JBSlB3lw5sYTRoP947eRl7lsgecc7rOLMsg8bmy8sxq
ja28alDBqw97YRVZoF2Qm1pUPakHNrRO2lTis3u3Z3o+OH4MvRSQ0iJYz61O60vzIB6cxt3RhqRV
/dIAyI/uMv9rnGDKJu9tkGssaT6NIdkdxY4nIuro4LGhlkKLlQa7pd/AVrg17tKF4H9TuWjJA/e+
dhzNu0wqS7X4uphmkQ5SJ49eikcJf0vH8/uVOkMips/74HwMcmDaCVaeYzodpHlm+4b5ufBznAhh
gGaaX+QRs8MzQ4ABQYfFQc8k9b8EgGdbAnbeDrrVO/hSwVcnM7rCcSP0Q2wYpfGg5yVeUa+un8ih
muF0UnCoyzXGZ8hsOLdfV3Q9oJ9dItdh2FNMpEUZ50EKzPLbQ0DRc410rUGYLvzBKQ056vTkmfof
fdpZuaTGK7jXJVmOf/x8SxVoC7KwZ6BGdhZn0BerP3UVs1HaWwkDp+bxO1WnmraQQe7CQPCIZ457
x1TriNS1ht933mvoGNY8DfgESMz2n1dcB2seCNK/suYTQSrfrPUYFRKUYI4LfsG2hcrcqQe9JZq3
rz8LVfg7HeysNDO02kJZEodeetPVQgGjUDb8dpTRQzBaJH7/FMrTteSVEcKAyKVA7qSktBuCq+V+
1Gy2LlcUVEeTWto+KJtwJkMDHjAYOD1Zu6ZVjhPX1WW61wx5wRK13pR67C2lB1Qe1eRFh1VKBa3+
KKV+3p0v6uCddv8e+qw8vq3Kx4jDugJHp8+Nd3J8ObwCSVqcR046uLpCIsukaDgfZoT1MpVFIRK6
EYm5b5vQsXn4zrCg261QO9Yb04n+ILX4iR7vhTDRKMBe4XK93zgQDEi+1WSVONnnY3mLfcwFTssc
ulcqAIQS7QhXy5EZfBkchYEi0Lf9ZaDgs9pnrXG9ulJ+lqaj/5SPQEZLxJvFA2KpgwqHqoHQ7Fmf
Axi2bDPuR5uqtN43Jh2HxcihVBZ1PONELjhyJ/USm0MNZBXNYamQTzxMnMcRr53XBq8jEvWbnXoB
A3/67fhQ07r3dU1Bx8MuVgS1u+b10/nwttpUkpGz/VwHmBHQzwNQ5z2nEsQTFEUp3nLD6I6RXD0G
zn/FW990gs1fL8rg/AXSRXWj6YuoOxcQSMoyIbyxCuxH0Mo06t+bbsKdBs+YZPW18GCIKQtdUy8l
fK8oeDrMmvBGtSrahB2pynJh/Zuv9JQRMZ9Y27MWtozOR/eBHJcRLAIw0d2a6Bdg/o4JPrb0TiR5
UM0FKIkXpA8g89oKGSrNXe8eGWEe4KISXs0A0XnqHrAeLyJVTp14MYGFwjXzrgaQL9ZR3//PZT8H
CJpzWOq3q5GjnOhQHg3vLREs6KdIDu3wOzXBIC4RXqC2/xyoat4gVBhrV7ft4pfgtvBMumJTAmB/
unkm6RYhEpWHDJarPY5ejFhYK2Z28kDGQjT4qXhnsvSGBl5zRLADKWDR1IJTkKrIE8GM6DFpDDZ9
2vEQTPHWC1txPxfZKoEcPIH46fDGPfjjvEBxNCVTTpU9bhApDgQDYocCnJ58YWGnRaDfaY7QyABE
9SKpilPGK4hm1qno7cLunzAKkwHJV1cvPKHaRw8N1hpe2BXr/CcMsGlSzHm/mzU6KBZS4qRVLIYr
ebpY5vLRDBNvrVJFtBLQM6Q+bN0x5Tt/8LTVzbcmvjEUliDh/w8DfVl5r1DVrPIXfnieQ1HPB6Gp
cyrUsBzmmYo/LBZccpv9Vt3JB2KV0cpP5L10VPnlfiiiqPiYzcG1N/O9hiXRVJ7QDI5jbTqcUB+C
uuKH2u6wlMH28zGrdoSf0lgUigb9a/Hy/J7u+G3cerJ7XscZ4rfZpFjqZ6t34VKNADkpk+QE1LGc
zWp/2P0bDW49ZjiwT9bMEERrmWSAhfGLZJZKDae5INCokEBly6Dz07Ntxkb5UHpA9C2D1ihozSPI
3m6wFUctgnIA8akUFUDvypb4kVNI71dG/9BUeNcUpaoSDNhT9uR0jcVRrGzt//v/IlEnG4ELXGeb
feNFFBaWBrEiKgL4eu65jP9f3thqFWFFvLD1DewuOQrHOlJvHfUpddyfuOKoknf7xVN209blBDjS
Yax2tphfShiaFWLwSt1io5J/loSwoZUdXjJwN2b/CS/5+KufKBf3MInu0vBYiBLLAwnzdxUn6+VW
jH8alfJQ3Kmz2ZRUoEXmle3Tx7jCdCUJme5KRkbOTW76+NR7sBg8UurutTcv4tkWkoKp63rnTx0M
KKqGY9IHsDa7CMFhiAzZyqIp5dN616kJuabomNmPjD5sBQHi7lkJmXcjzGLE/k2hbnr/09XB+buR
HL9xFEnHmHAuvPQiJXqIMEK7SS2PhEuhrTYNhJsA7rvKGOdWtgITJoe2aCyU6+3mTaJu4dCka3Lh
tp6/g4rJhIja9MbxtVcj/UTRmtMJeghWDM0Xf0C/bKJ1bfjynYiq1C1wbYGI62ybHM0xm6EAeBnI
7aI2EqOVDnu6zN94QaqXRtu4yny4c9X6nyqhsAbUZma3YuIjvIk61i5as1QZfIYPanDel0a+c2+v
7Vhko56FYB43pW4l8zZ4khis5BWVY799LXsoDPNWkUFJ3pZf8XtXOrJ6FEnlHmLh88DVS17ikuui
MJJuXCCNY4TJfIAVJYD3RTSj5n1XMxOZWIXcU1wxiUX9eute4JtUg3oJ2dT9/AHs9da/5dRz0B9K
A8lKlZcwpjiJI//CeI188Uv5oKqUvuGjJRR1ZTJxp3n02UO2CooNjRNz6C1o3p9G7pu6/IV6xCHZ
n+YLAywaaksV/WlsCB4Iubm65iN5pUDTO/hxJuWj3UNZnSK9NozPYx8KLG3Fv6tfXA3qBcN+aZBK
gLu1dVz+ojGfcGiLjUXboUIq2E+6SM0OiS5qkBTAkcaPJTtOd7CnfM3GoO1WBSTijBqbGwOXrasP
1Vg+dR69NHVS0xuf2fzwHrhRMJ79hZK5/Uv5nDnT79ldDONG392a7uSY0KHJl/sqb+jiO9taC5Yv
GlLJywZ/C3emOj2naamOqqVWX1dtw3mglZZR1pAF4u7PWs64Tt66PxKleG7gFbDWrAZa/FiE0WUE
dnn7yehySuxEa2lr59d/T1VD2IDGZJDAxNKnqrzFmJW/DfwBecHS3XXZPbtzOpu5DD+6sKkBs/QP
mxl+oLZpualiuLOANYuXXOTn2NDKKdF57ZXzDD8ajvFpPZF1ra3iBRHsScX57AGA/Xapo0459pky
U8MvFIT3Qqnt2a3dRDOENFV3FYS7Gi2273lLaYTbEVqbBlMdJSZLYeE3WG4w8L6wldCgcVpmzodj
BzU2zNEdgLpoBeMIhIBG8DVcCRq7f+dSmYDVkmueMRdYgCjNH1kk7lF47Kb3b9ORTTzQt24vDG2z
T+3y3AlxOoAMr+llbshCILiUvOv7/uLs8wI1bf5rWzH40JUau2tuahIrzzaacwXN1l6LCcC6SLz0
zw7If5f8LY6DdgvwSZtW760DGAior04ZN03btjziC6nbLgCuJAVg4vHO6O6M+asM9PzfpNpjt4BI
Ep/z1jMivda4KmE/vOaq6edslCi+T/i7LuKhuK2WFbAUYmoRYfkiTwwjIWTyNY1D9qE8ojVaXsl1
J8yA27z4xDB8rwOgC8DITiunA4GHA4WuJDvLL5nNWjHkE0jTqGMFNsKPwszcOsHtPU7bFjG1CBLZ
SKI8K5FI0YmzPXVTqBFgVK5KpJRnnkfZdCr0s8lGzkAK9y07/6GSH8IiM57ei1NpX4MAs5KXK8AB
Xln+7BlMxleNerrCsZrLSBpuOABWvNDh3FRsKdrSHOJE+UIe1RAszJLTj6vrHXt4mkM9DFNr0vf2
HrYjehx03xR7C5AmEAWoKaumJTLtw1kVq0Vc2L9XU68CcgwaS+tObO+xCC/a6dLJu6JFBICDnNnL
sJxfiggQN/L6oyA1YwqPP9jsOznsTkihw1rpvF5G+JWmjwP9FQJ6Fm38UogCQGnP1/7hVlmeM0qV
zZ1x5vSb+i3S4pvQudmuDfjUW0sM+C+9gzUSDJ9iERv7gEfR8sa7Rd9VJUMy11NPSCJzlFGPyXVq
vawJ/5ei27DcX4qfc1xt/bOwFVXuGe8BHupwodfIIvf8A/L8J3/G2fnx+7uOKybdDrFn/gUKNa06
x4kiZZtssTL2HgicibFJbi0i31dTy/3j65sV47/ZT+ukF+cekQRWt+01yGOy2imZpgh2zuPOjChu
R4eBR5mJfS0HMI8wH1g8Bs8sigWLzS0i53k3EU4dhSx2mM7xo1XOCJo7E6hzG8exjBRgf3j0DRlY
6ZD/NuLoLHyWU+5P3mIUgoQyGNgORxGS10ROA7xVF4uXGx33cJPcESU2VCw+qqSWkq90BTRwBzW0
8GC782/NF9nFitkUx0QG5QqIry96Q/K3qSYZy8kktDyDZ6XeNJ8tq4SR5zlC0k+VF0d7yENZQwQL
eOtMNQk7smE3O4f0xGbMJ/XN4WugfgNGy4UzytRKpIZPYAykQYevy+vuI+fiixcHD37y972olCnj
f7/rkB7ftdxO3mYtCnm/DacxXFIE4BxgjVrI3mwFwS7YB0OsctBrNpzFp3BCtB0/5FtJC7JXSTFy
CJAmV9KEi3FGmIEL3JPtnvFv3cuL1XaOx675D0L4bjnYT+AhutBLqW2UNgwNgiBeQB+U7t16iwdj
CEF2n8T1/uWafY44yr6dTyJfDU0DcSWAPFV2bZ6sva6CMMuq+Iweaw97aTmoIT+mYQpa+7ceFHqK
Q6a723oZktqwnKkSYksJ04lhvVRy+LNIEYKvg5tCe/aLsFm0EismBppPTSKlRwIlQReYlBPjPE7O
jkviveCMOp9Vt38tAxcmyfE3FxeeIXVa7pp9MKgH9H2Up6OvXT16XtBG+dGa1mt0b4iYyYqgCsSZ
aZpWF5f+0t+nS8CJEDt9KJhNH18/ex2G/zQo3d1XetQ0sdt7xW3DRx026jZa6X70m/ULLQtFHkMx
4cHK0aBcgsPZlOu4icJom++4JCDgcQaUjsxmOA7uzfIsUWg7Oi0oQe2b0096AJ70QVZ5Nhu7U3Y7
b0r2FX8LvNQ4zxS/Hke9VU2lQuhP3zBO7jzpKwh19+4VG8J5EzjA+mnB2PCfjjQvG2wQaDxh6Lvz
AS94KElO5XdlDYd8G9VQGsRbVSIPgvh2voLa7fkGsTxxqPJR3kMGwaS4LzTGXwl6VD4G1T4wJFuk
y8yfKOi3AuiA+TdDbICp5nymoukrjR450dl2scRXOuQvm+gb9spIwmJxjRrIY6TAuDzRsykx6yxx
Z17mWYwYomtDmHpiCOOyh/UDEtuDojYUDt50+WyyCscFZx6wfQYHsJ1CzO7mVSHARW469OcWTfrU
pfk9UHSEE3q7+QZVbRCfjEIC2VYGUPkDw/p3r2UKvbXbUZ1EMzSLmE441AGDi6RlevO09bXVcR6e
KAqnn50DhF7LC1dRjt5tHh0WRxYuxVoKx6p/fiPnkBxxVeDWkUqetUbugduMndsrfzAcaxiafklL
09sK7/sF94PGUXB1TZl3FUNbLml4Ge13oFbwNFqFp2oZCQuxTRM0U7SWOJwxsplzd+68KkHPlZad
3/rqjkW7wC2vbMQauLkrNECAMr4USK/KXlZi3aDwl5Q/63pdBJW2/9KMWcO+x/1YKYTW+BR7oBKM
tF0Bv2lihYavoz5HavKeH5FxMp2ZQxg0CsHlxJGIJsbe8inhC+mfdWtfmv3E7gJlx/xsVqq5GfI4
y/F7zAm4kY13zaHbvipJfuJze7qmf4qklvV92c87n38Sr8r8U7fm2vPD2X4aP7gNpyZYiDUReO1v
bNpQpwNJ7jB+lT7hdcgIKxI1Cn//llweHiJwWF4nfpIzzF/bMhS56vQs3fTdEM+L9N9ZDBACJUjM
c3j+QfZlDBaC0aTImBrTj9UtYAbVsg3Tn34tRWEVl+BME8Tyl3eNfVOqC3dOkBlzIMO//cTLMofu
cD3EbRKHHMo/j3EFWNOmxpEpbyCaYClnv5L/wtDlfoIpxIR/ru3VyMx2z5MLJSNFtGxIg1ozMmn2
UGGnhruH+sbWI7ZNFCFurBhJN1UvOcFpSPAX9v+mpT3YBz5heNkyEpc5sSQiKs3CAMhcbFX0Qd57
k9fWmkcFoiEMAwrLPrthnzC+o5poRgADuc579V2huyW/c6xNbLQh+smgZoEqU3Mi7zdAau2eZ1EM
ttdVyEE4zCNytdbzTlr1AkOSPlD4//P8U1SvetDx9ITrU2DLYrkTI8kSH3ZTiOoglb0uBM1+leFJ
/7m7ZVjd79buNPQF4LFZwS9ed3UyEL6s0DJpJY++zQ86N10oNjCAmugviFPatCEyihFuW83QQv8H
5+MiytWYURSY/8ulYtk3ZjV/nBIZ19YoyptXCL0xt0PYf1A3cTJ/guRlKGVzdHXBW2yg+7jOGGJ7
lKcxl29HMS2VHvQ4tQDOQyVkkT74372jzIj+pR2Ec2h/bqqlm8vxc8t7YRL0wJOL+NvDkY6Eujtv
u/BL+1nACjJADYu+4VxRDNhvGVB9pHjCSRTJLmAzbllbVj0+lnwTzsud3Y9a8HtgWfV77RBh1kHt
WzRQylGXldDlN8YIPsbuSVR57QE7bVCwcM5Gq0nIdYtfkqfmSXvJUkNOAf6rQ2fgQ3jdF7q3XdvS
u68ciEUUrnGQT+dg81Smck/qbfvLDPODlN3Off6jjGW12jl94xu4BDtjttXRc4LNjAXfOc1d+Bz4
yHY46ItsD2H18NUN9HC3p42Ra6bPdRmoosmgk02D4T9/iGLpfB5YIAJs2RQvgAAqALkTOMTQCInI
vuNvI66yl5A/H5twu02ASMu6hJeLuRA5m9pj1VyFnWpr1p+CBay1eF/l/NzfIEmg5IdjtslKgsgc
2NFvkJTCtYedRF4/eerOg0z+Dzt7tIF25WxoN8WBTp6jeTfoX85lQtWJUvNHSFu5J67tMhKMLhCf
efoNxziGeUhkhcKy+55qT9uFVV2ETMU8vjG2b5lIGC8tC1R7gq1C7wYtw8zgIbEEhHMzf7XeGaJd
QR8UMDSfHTbTC1R3VPbwa9BElUHnCXqp7XM65OYwbxaPcPFBWFoge1bIO6UmJwfkLNgnyzh75SFc
FopHaCzOCHGMC5Ibtvs2WS5TAUn5WIch7wqRXt9A6evdG0KIiofZ4m8/1vywsxm7Jb8aK+q8pe3v
HGmmVtBrSgbzdb/nZsbDpLqkJzdfgD3myu2RX2g9VDyaF+ehzbXY/Bqu/bgPSe+iX4HO0yv4RUVA
EgGszoIAS/JFvpNixYNMuDu4V/x1gQvGBZhyL7tcVmEqkhAzPnX37PMDZYJetwCTQmboK4KC6GbB
tZtN6rDWP0FFPXUXf2nQFfD88k2kIRenLLhGeGv8Pmg8QPmPOJWVOE+jhzvs/ZJJdbpvPsjy3gJE
kubN00/xLQ4nS4dwL99zON18nndgLO4jyRob2iVAJLofnbEMDwVjPm1bbQIFBVIHE4qddbv3n6fm
SY/MqTb0hHenmQ2YzBde21u43vXnruMKOGtgjuTXth/+Aca5sm0y2gE5bBg10MumfMf5Uch3qvRs
WpF8UjxAO3WaaU2jAAKxM/2Jr6d3ZgRLr7aQurFLN8dBgtOL2CMRnyHPMqny7pR28mdDCjPZUc+Z
wgom8SsE/zEzeCPoBRCZy79Q9Tnnlj/IYegvrhzXvGNcFkKj9UUAQAA+iWwwmYAK+bIrvJ1djlob
zsdEpQ/vH/F9fV+RzKU8chukj1o5FtQ/S3ZPvNvi5j7rFGnJ/hE9/ncUTTmOeYiu2tfjnlbygbss
++YRuUXPc6Eqt7zevCvDaHoTz2O7HbwNowlospx8dUI6z9UUCAH0cipFkBTG5XCsbggBsu67EeKB
M3PCQ2ta3nbZ2SpXmMM7wrF96kvWgaeHKkDuBtUGsQFzxGjxyP1r26oinjpO+bxXh8I/uc9Wl+/o
eP/RIDqquGyJVvd0w+7uoU/git6hW+Vbh4Kz1pdh6JeU3iWEHU2BeMCxZ/LudedZmNEx+KjBPthh
XTnqhZo2EWPTXV7/Scd8O9sHZvoAnWEEdDDahmXA1HTpc+YPBY3uWOX6sQUQGLbdxzm8R1cUfTBm
md3VfCx28qG7gZwbXGdMQ85Ds0wKygRGHW+k+vI/s0Kuia/11jSBlYpT1BbfsWngNUX+adNMZP9F
aDSjsuoSwwyQEhFhEDOgFfEaRd2kw5NOE06Q4zg+i1fYhkwxEV/uT5wDcIh0LYtYj4tTKQVT0IDi
5B9JkjAWZvH/ehHwa6uVAf66dddX0AUcKVH32PlPzRsB/zlb3zOMu7PPHtubK23MQGVWppDjudFK
kqke7XTtwzmWaG1bHcuiQI4AnmD7KMi4Oxak1CopGIEUPLnSaEfLkDVVvEEanM+CEoR16RPOQrFa
m1D2YcdZqtQWOC1WHBJAL5uBNH42x0gtvnKU4K6Nq66Lumu3kEBK4vm4vmZlI5HnFNhX8OYSqaGn
pzapaEalj32jTcIQHsBMqrXaIGTBReHHlab5+cIqHmFb4TXIPCYh0fZPC+Kfl1Xj2ilxEkVMfW6G
rBcDM1gYv4iOai6Y91cbntgX3LCAMClyuXzm9/mojFS5dLRJ+lqusBKAg+oTgStJ7PB4ratsUdhH
6KBP4gLh05laa1hBg76ndMdzAEk6nRjoWUiwpunBthCcLWMkXEUpkHt98lmoZjA7bEhiWgUoYsgO
8O0XleZ5HfYfWq5rGBa/hH2Cfuvdj8xWDKDNePUekqPKAbhxrLCQi84gQemCyF5Ajqwdz/PC0Y43
NGUeNeXFurbET+1agrf1JHm8SLXRRbhBIcLdHKWphlQ23tidePHEiiUcYaZ+JOfvla7CG9vLyQSC
PS3Rw5Bp9pHVdFrmEFHDUmjAM4QvHtUVGOHP6aP07wvh6dgSp9hEmD51n1X0nWmsmV4rVXIMzAP+
s2UCTdzFF8DrOZkZinIMaSvnPYIbSzFTAI4fGRsScW/Fj0lK7wcihsCau68Pxer6fNmEa4GwAUY9
hyrVANExBICtLKzjBO2EixVcgN5cd248TiBkaFgn7BW0fdU27iysxGOqaLD3/TfkimNvmxFOlZzx
m4jeApxCNW0CddOoEMjmetce/IZx80auhFJOBRTlxnztAnqvFs1RQJldOktqEsZvqzgygwPQeHqK
m4wkBGALbz3g2Og11GzSrHZsTJHgfeTjPEs9brlAHgj8FH1DzjjMffiunuZN1Gknj07Oltpimjl6
TmHRGQm4CGIP2mOgP4d40aPSWwjQhWTa4A6os7qCfjCdPFmq2MmI0iBM4RxDLcn2AeJpVvbSq2n5
l2yhmyZUvssO0/k1hvDYUovWUQq8SnJ4QXo6GNTDUwhmjFpxmktGqaybbKogee/Wj44bXh5PUhxc
U/+mOWelDvRbFlhGl9zmjNLS228b4l1MAEqev0xQBi1dAS4XDPTVydI67o6W023I9rzC+NOnCK91
BXVYRyxLrtnonSCNKNnvvdTI54W2DlYhIdINnt5/Ma98/W8noPYODw3tK83xkNNltoDl4F5kbeLJ
nDICZ6t4oIFpXivzrHLMefDnphprdIAlObhsUGCec2MpnxM60U1rndDQTTMS5MuH/2+qu+hvNgON
7ftZRn/IQSw922r9VWRsNpObAHUR0LXJtkEjMMklCBr9FfRFUkJX3P4x7OR+Zuz6a5KYPR2epqBi
7f03BAmgFJ8gxab2WEzxzWdoZntTby+MfuYXYmi4jwknxLUgPtN1L1FQMBKakJ8xEYrRBGDCoDRw
xI5Bqe30S35rdU7SGVzhYYIEbBZDyexTVsUHmlDXzPVdbJhwexwiyDAJaRypYpxOG7E6mnTEFEo3
p8YTuntGcUQw7B1aJNwxE+LPyGUhUzMPsn2bFjLAkZdo/tSDdcUBsFopVROpsWLvF2aBmmZ2rMap
BSi8xj1OUNsvKw5nWk3C93yaRx8/tHRaH0VwGSZWXB3dDbjnwi9NvH1d9419uhd1ojhuU3caUYwB
1swHqJTUM0Hutq4LcGLa16PkO8dO0/UJd32FJVwtQKBepXyPD7z9ieXDmcP2cYFwrX22D59IjVKT
ijlIX98SoCo+mgp0YaXH5nXFzPpozHS2N5nZGSnhelVG82EOJ1F/QJpxgQ6UKTTiFnQqoe9sihmF
Tqm2Idl91G1yaJSgMCqOUA8CtlNbZ3nZL1Sx+aTiSfJlFZfmj86yvUuZHeShy+I/+HvOKmKT5R/3
N38yoLrB+XcIvx+thL+gbIH7FuYuZDmAkXBHKqoAK0YfOdPIYlhdWXHWLU4YHv5buXa1+ZJFFVox
xY8uxu2JGyk2TXb1vXsfIRhDwcg6M/OkFu6owr3oM0mcKY60ON1IOiyWY4cSoqTCQuOIL/SvVOu8
HsdGiDoiUVQRfkozA+bUXp1b+7LauHdR/juT3J0lgfQyy7Ke8G8OIa7jRUpG5cGLn+D4TIFfpF1b
oBDwfNPgYLVQKk8S0TlBGVpudc5JsQleAPmvFqazlliOxXJO14ugpBSttN6sLDSu503X7Wm7F5lT
we+JutqlI936VtlhYbvh0Q2UtaEnM63DoiwtsTUsh+Vgroactuo6VqN6gV7A1Y72lEo+fa26BJN/
YdQOIBcuK0OKTa7fNwFg/w6+GopWaQ5A5tn+mDBDeCpd2HGWXAFqYFyxh33Yn69qmUAB0wld56hn
BQfTF44fk169fFv+H27QguxmVE5O0jATwR/AIwkfLKk93PGKddsLkxOfXmosW5iB88j/VI3VeMdM
iG0oM3en3eA8SBhbWzV6P1pSRRN8x+b/74gAJjxqIy3epXSKjDtMG9wy2Kv4vZt7JQ0hLu3nzKSG
B6iuQRyjcAHRDAy3oI3A71gsxB4HSFxwukexrDr8tai1rMgsDOL2QFyQT/9OoaeRDguvC8e64KVD
Vx08p4WCwU4KtkPGVZTwp7E/IytU8IGbYAow9mBbwfKkQlCmaBaOsPnJkiaGW1GRopHaemqkmV7C
B3rWxNh3aGRSyf7S89fX3abKXn86IHAO6N7rdahT62tRRgu4ukY5SrM0kVqZplHXqjCEae5OJcb+
UZ74WQfsNPfJv37otcaFOPizbxMjdCiYG6OxNLmTIRmvrAFGP/IGEn+YZq/5eEGlVzIk/TbjDvgT
f9ksojLHLe5c5Zmz4MXhTfx1HEyVhge9I9pY3OU+mfUz3dHyBnovcQstWu8cTHnnqhDyuEgBQNLz
RIh8rzOI80e6pQwFoRDFF11RurFzdGtaihufPIwZIfse0SEEFarl9Hcm9TLcpxDOMX9Lh6H3nHwG
TpBNYX8APEZt4HjAICTTtKdfuTpS9gdDNYBaIgiQ77VONiLEZ4L52ejxT7Nf4cwxm1K4DaI/964i
hEWab096ub+XEop87moL4c6PHMxaf1OLATpg2d92quADtZ1PTWupRBHRpNRrnhdDEwfHQAPh/AZV
Wz1/BE7LmuwOktNBG8uPHVbBire62aOQR43wgKp1wEyCTcfkuRphSm1lR/YvvH1mjw4/tDMwRUpL
MBvPbhpL0zjbTrIZJF8/Wh7Vxlr8bEPBld3j2Vs3HjpM04t+/DVAgasY+6ioLCO0MNogxlIY/KOi
iuKbq+0ksL4Hia4488jJV4UemJcmMbA7ZNx3l4RuVks2Pvyuy4Bbz0rEiWx9mTqySPHsgXJL5h5L
dYt4VZ6K7//waBJj//GvEHBCC6t4FjEPhMLzP6AMNFddG1uzCdIlIo7wusHKcqAzGPJpwNBdhkTY
5qUzJOcXI3spe1RVPWjB53NCy1EzjCCLg5TBAvrTUJeTo3f1QQjV15eqFek3ORyC9ITyZ5BX61WJ
+/WrKRheGfU6cYZqUlbhBNLHLkkV8HtxA98lFBKhFiNuiFlhLP4iahrBqV+Oo15Rmz7u1u9C/MWh
mtCAfsKiI0He6d4O5rZ2NK2UkHkE11ltzh9qvrejW67m4NVG9BQRY8NvLYGYjNgN7ywt4UxguFIH
sfaKIGO1b1bS6k1q9RrFQP5U00yHJWvXi8FtR0Y1l5N5oVNBqDYRf00BddhGisHFqT2L3cG1gWpI
GdhFT7ZegKuALlmwT4cSJtuqfWmu4sunTWFo8DHsCkOry7p2OYFy0jXBYB93caboVJJhUOb0km+8
Cu2m8ifBzQfBcssxG1UhmjZ1QF/SmNJVwGQ89PmepTSuFIqWM8ohyAPAYlmTgZl5t3Ipt41+AIHN
j/IB15CdsmNLqUGtHkgWF/oOCI0rPhF5E0Yi3dayWjj4ozSX8TjuYXrylkcTz8BZz0kq2Xvb/LIt
HTOBAzsa3prmJPqzQSjIIhONKvrlDeKVDkJXaB3oqKSA8VvKXrfPu+WjosY0FjX9itKD5F/eXRWP
m5D7nS3F/jzlre0X99jQuvVv6O8IMjYEIa7dpwY6d9CLLHYNBHuSJgur2D07LQ6G9Eo442VJSXnl
yZFDbODndIozcR9BqPST5UpJ3/3tpyTEHrEZNZYzg7sYnBDnWhSPbw23aGBRF7Ldcjb67GhfZ+GT
7kgIsMUkWqddevkf43AnMQLTJs3RjHhs/+2E/f8vpFVF5N+AFsI3LF/2vDaip16Z5dHsR8oH8L6m
ZtauQwF0eXFpgSG97Wy9XUjOa6EDHpZmD0V4YqSBAvM6HTyBONY8F69RQ5jTKxFHciBXG7u+S2V/
hzY8rrQxFG8pWOwcRaGRXES0IEZkrthi1EDIeoEnyGI+F55jW634BJ53hU6dVZOpDdXnOXFlZHA1
zVcqtItk1LcxaR9XHemYv7vwf4I+CDBW8hIJ4vPPqFJGGUMmH0pfk56An23DMeC5XE8sZ586E+mi
JeE9GrWD7EjeNeTrtw+73f4kUwKtBmcxvyEA2V5mOD9VPLqSqr+fdM7q+gfsHYHSH4QCUdu7v/U2
G9/t3YoB6ZEb76qZUfEDmbXXCabSVOhaHJmP4BmhG6eXCgNI9M8yFW8fBbK7PyzYhc0ZK54o/zE9
CRjsQrNdNXBXhhamaUFZWpkyYkNwnhEDRPc6ETgEmVWVZpI5cxYfyz1H9ZKf3g9rsbXQabnRlMlI
LvsjnZRgXxjurn9Nq3PWGucEEV4Grr3Tl/smdbmLjmWWowLRoDVmu5+DMcBktmkF9TUE+eEr38Uc
2K93SyRaexzsO8/gLuupQ2E613dlhE+xAWQA8L6mLEcTsPY7Wrt+oMYkg81WEploKGi2IzmuD+pR
OI6iiirlN9M6zz0XEsHNuSx5tj4/1BYc3qvWxpseOGCO9jpQ2Y7qa73rvFA0oJwb9Z6V8K6wkjqi
nMvauvX5i80f18BtD87GCOU0oF59//7nVw/mMoWIlvT0zrK7kd0p8DQWjs2RvmTMzcfTKaHhj5Io
1EHlv35Tj2jdorek7CSErAlzH4CxTho89sOHtbaZsaBrLO1P4dvWfI+4magpX1Gd3nDhcpbLy1Ut
qq9YGFRL+8opQodo0O1RqSfUpP1Yt1ha0RtzifcsG8z/4jlkdEHeLFyloL/4kQ61QDecDHc8KwtW
Ae7iH1MHr51edDSkg6mSEwDsB84fXQhmV9K7OqgVm0PmA+5vcWNpUMh9J8gb7Wq9t5hqgvxWRDsd
FKfjxx3TyAqQCJAyHYcMPm/BxBf6xKHFxFdNkvCjUd901RReQ1N4nj7yLtbn/QeZMB/3QdrDAtAq
7K3tQk8PVELxz00prZHJar7nqzCht+UVvYXsXfKdrfmfvenKZEWwiGhYHpd5WcJXy5RBiNnV3iPu
dCyxBO0Xl278CKBQAJ6fntWMEOQXqyzbiTSCt0VJRsPwD6zzPFY9sqAYHagvQh3tXw9yb9SP8zpR
sMVMJbbh5wVpM8aeCZZlUzEUd3IEFezeAuYZ4wPCc0hj2x6rEhTeZiFu/CkxhcXQbmXveTrH+O/d
fGlUtP1Yg8HTGC5hI0pON1VnKIhMkjQOt/hgPvisO9aAdiNioxa6XMd1c8hgmNDPY5xZQ5pOdkPG
MrZuBF74WgTzz0aNcd6CjF0tXPU0trECdfMdg4lADU2glywLoTLttroROkFAHGL2Um51dodao9df
rDs8d3CbRjw+xv3GFpOawWqGeEN3md2V9XeBsYtTnsF5Oqr7xsFuv3lN35sL8lZDsynkAiIPBvlD
PpaAswFiINuwT99Y+vo8XLF6GI/wfrFHvhxkvOfkzkCCtWSGoxpTGNIMTx232l8Jg97j3mXmNu7b
LIYvjOSzF1m06Npnxd5cvcxRHBdAl70+QTKWUgFhiPFksaticJH5d9biZHxK0shsSU77hGpRzxXs
0dyD4gsFxj9tPryfUv53Vk1JdBzuppWoeJKUuaWb5gu/Kp+73JgFDFu6hsqcFkE50jaWi6RPRHeX
Mn1qkFfox7+eqaniYwR9DnHzbLdaM+S/EWqljGgi28Ei9ywWkWNTQ04MJ3MfAQiO4zdHBwy0YAdz
cCHg2gut38coKHHB5suEvgTw2jBnGAdBgveIOqXsrfoSuTCcULdbhgtU2E0Tu+/3Rvyili2L1DxX
EYfSV9okRHCxBzsfQxSigizsjREzZyqAgzOeJY1nrMn19KYwVaAEkcURutGuTkBDE4z2KsuIkJqE
xx3ge7kN9NNdflXZcaFfdexbzoJA9QbUX6Nule0xiWmn61J8jVDb/ZIVFEWcv/WG6oypqrjdpC68
NlGagdSSPTAyfgUPU1vaf20TBmQC5QCkIeA+Fy5AV2+W8AlGg4zKRalCNT6yLXbHx4UiQKW9qd25
S2gHW4AgeSgDL8BVCqE7UvM3cnAGo9dXVKFaPyxaFrT7G3IikEpUQ/NUegwcduaeBPc3k5z3ycnf
m4m1hFxFVZcdnxkbucGZWoZkZjDWvJRbh6619NY4T0A54bqqjqr/ONFVIFI6OnC4hLVYwXu3vVKa
M5kfZgo0RhglJczxrLl90ko1f17QeBTpYQj90VqRQtmspCuiWbetF5KL0PiQc2JZ4a2JanUGc++8
u3pquQ+CDC/ldj9RyFn/LANa/9ZgJT0VAsjqlcG3Jsd69gmAg5Vwpo4zNzBgTEWjaANJARqlprpD
0NY/1rqRHIu5BOmReVdkatb0lO6JswggZRgEluboKRL7GVA/1P6gR2gRfFwWb+CeiFN8ERORX8eW
E5LdN+vLNqdsxmbO7GYUhk0bWDgn416bqgTFynHLeXfWc/XiLiVcbeEoGt1MJ/zy74Pkgerv821C
2B6H5V8ld1Zae+rD/JxEnF6vh5LONXp2M5hPc1Aqu54mL/6Sba+MZ6gBCv7mJqnZydVfuPt7bwOh
tqqtKWOVC8nSzO1QfIPWDJ6/YQKK+gU5FAGXuVw9060M4c7xuCAzHdpox38z6Xo67Fxnf0rFGH02
Fcg1ApCPzWbv/Jrl2JYjSb18T4TEfVmgI07UOERWqpWQa7j8zEl3+4r8JdEBd6CaQ7Gx3RbBv6qv
fKFpTtsQTZklMNna1OgYmXATyT5EuyYDUufWENd8ETigmG6MR/RXAP6YakKCsoDpnFN+mIv//ZUO
Iq6oqca4GHrvYHuGPhCdQuRDM3yt2/Oiy7/ZQN2uo0S8M2dZYtyce/AMNkC5YVYm5ci7ehG5G6fa
rdRIDH3kQObviOIpRkfw6hC3hnGaaXSBRa2eI08W7Se9r2OcSPpc0AL2LKOwg8dYBQQf/0ZrJNyJ
4YeXQAWhMfbTT/oWw6tJEOOW+9XWUYO1nyiHGBSCVtP9ur9a+UvhEpUieGS5tpUmZGCBnvwI5bB5
sUl5zZO/sQ0gjPdnTsKGqqz7WaY6oGHwAdwt2UvhOr5ek4EZm8sFMsBFVgHJBhY6oH5mxeOhTBei
csWUwcZYET03HBGwxLr6QHA69uA/uK+eP0vWON4roKlG8iec0+xOCznQsDgWOQoaumiVz3UKyaWx
8+/JUrWx5A5sARqN8NniUP0erYT0bTPMBkLEXDRnH3nzoKj9FxXlKZoXklGsxcIT4ncygzN2mJvQ
yhJi6/Tl/IbL4TzcAVjbWatiE+aeE4xYfWPnHDK6WBsDZxIQLCKuf5dCEsjnj2dwNgebe85GWlhi
PS7ZyHoggI+S12Iti8fEvNyL3S+y/EUrx0Lghc9g5Y0mk2eZZ0RK1q53MioJ1F1r2ifh6+XKYe5d
/T2AWGQq/vtDVFQP4MDdJt7fUEcrgriIIjdDDypKlucPp1IVvRCmyk+yp0IrT1dQj4mDK+kRsHCY
25hV+uVasvgpThDz+gRuOF+a3V83WYSq3y2wztSFSQUUchfSAjEi5SyxyK2/DGWD8g+svXLETldF
tvU0owMbwnrgnPUH5+mS+E7fhjhUHo9T6g+giuVM8KGgnPpMZ0BByz1daWGmJ4V6UzYhAFW5Ct7e
GvAkDBl9yB3cv3cviYguqZzP3/raQg7elApuQRYnJNPjDKiPWjZEcGMMEQhw85ya50h0Y6tfda/v
t//9A2l16DFvGH40dwXKN1FzNOnx6ReYuK7PsejS1h9iG0g3UtFv7bmddsePubP1XzgJ6cPEteed
1M7uin3fj55GN0P2wQ20SBGhWhjkdth7+hqOm9Gp6WilqaYGxfADOcxzdlruAiB7GH3Zvxv+UW1i
l3iq0iMZVI2fraOnNlY/SXmE0LA1ipDmOnncF+nuJ+k/Tm2X5vuxW2Ge409EWvAinhY2fc/ZvpIj
wJBHnoXDNJJfCl876vMYaQo3obyM4MQjinZLdAmFiTNSj0xkzxl597lg6rTpkHqmBtOZacmbj9DQ
zX07L24/kiQJwfdxxBVs//IuiKpSWmoOjY84pFFboUbiy5AGOx0tU4lPvZovtELS3NgnOQGEvD8/
6B8OAV65+zCh4nybe2JH2l82jrsXs57o9S04wm7f82hJXPdfbV78mcXO9vJy57+lBYyMA8FI2ZjB
cXwYKh0XWRwidZQfexfHk6SNqE4jgIiBxklRYJ9k+p/w/l1PXTOmv9A3QZ2PSDB0GB/hjAe6FhCS
E4aLjQk99iNuveY4zivZV55OkaAlgmviWpERup39LoFsTlzEdvI1Aa7X/vyKn2cSb6I+cTuGV59k
t2TFGV/32s0q/uVCZTzfftt84EBQWapEEWDR6I31uf773IR5qYUwMLHeEkEWS2p6YZy1AdJaoCrv
e2m4eQx8sjRrHZMrV66mTmx45uFnjNPlISc9de/wzu23OWypgC9c3waVVdSlq7BdrKAxgeD0z8HU
Hn0+/hp4zYStgc3yoyrK/823h9ZGLw+lvVcWhtM+9o9aeTcNdRUlW28lxfmwMy//yPc//8iaqg0I
9iQVu07C31E63veVxn9SCCOi58ELc4DNeseUaAs0V1q8LTqd/XAr+bEHSKdF9DexGL5GmtD8niZv
z/YcMF/nopYJVAG0JsvSWG6mEiyYvyW3+h3KPUBSHGIg5ihLdYJxQCL+kp5jBgAl1+KlxRvipQ1V
kuWn+0XE65L/NS5hjy3KNGAtBmTxA0WPFc/fQF/A5jp5cpUrZQznbS7o714PxzeT7ZgSUo9CeifR
WVWAvoI0YNGRW1DvmI+4GyOlAaLjUtdC1UKlgfSj6/iGOkdj+tBGIcZKN8GMCgH0wlTQ1QXwLVs7
3wKas+NHU+c6kt9l22EpEMyRDTE7+oBk+5x48brPelPYRQN1RqGj24Zr/e9uOXdM2oquboIf+BNy
GYmk6nCiIrFMXh0GR8t92zteJKrK+aMs9KbbAcEszE0HuOGUnhtq2A7xykfTgb3wX14gVOojWyPI
/XCkYObRgD0sdNls1LrPxrgVtDO0LRSFHa+JfM7PTdDlCqMovDEXD2Il3pBhXcEmhhUsKTKL0gbP
jNWxnrjYcuXIzWn9w1ygEUcD4tKjq/NC6k7XcxCzWhgGwWlvmQ053DhUohX6JwX1fDXcOuksSF6P
PjHVLCv9OOgtcvIpIvh13s0bjTOEzJsaP7IaDRlFwfinoNZEdoCrNK+7mfkSqSYDh6qVCdLSQY4h
JF32ZcbS4amAsbOdRajCdGnff72ZvEj7kChZ2Q249z2x+GYGwDaG25M4FLtAGYz5aa8aovO9xeO+
CK7VO0sEFxJSjGp4EFqbuL4Iuz0wf82DqlzL9MylbuUl1RG0gR5qPezdH9nXE8yRwPkzrLUs4D/+
SLKbv64pAK+IEWGQc/xcWE1kHh4gH0jHGkzhrPDLWzA65pylAdZQza7z3q0bCJD3WWz2fjEoviL6
NX/S/eJmNByGkRhEUqYz6tm8Mo523aCO0Vq0Rhe9GDuwJZXJXK7aevLN8SabNfneKCGoRmV0UCGK
FEKhOh1n+ydvo0VIUAWbEAjKGjejCHqK1DHjgWXmLJwfz4iQCNhUf85vrZRk7r6achz3Kluqi2/W
E1bs2+aHVkLZQ/fRNAVRrv3x0VUVU53uz1lmdPdiFfBJAACFVR5fCN6H61C+OF0H7DeN6vrm7Jgk
OaLKtersED1NrlmXd6JhPV+8L3UxFPCQPcBjRKb8w99168cb8GevLit46DK3Uz5KIZHGKgZzikzJ
Pi5bd020S6kIvFN7CgcC4KiNq88kkidoLUaab+8aPGLlvFb8NWHB1Ceo9GMBpAU+kkxsxusMfWL+
7u1e3WDrptRqcba0vxG05t0B0DBXaKRuPn+owLOJwDMa3eTAoYyXuWeuo2LzfkVs5xVgfbShQQ7+
7rGGgthNWMLVts5cMf5XRCxaBKaFfqzTYH0HOn3gl411JDSscu4d1d19fYNBmUsW7k9rhA/KmPIg
jeR+nzgHt5qaUQS33q038vo8d+TNRCMp719kwQJQq5MbZcYNAwQsugCGC44IeO06CGl48vDlN+7i
a8Ephuypk5OgWoLAb3SY7J6BuYOmfYRWmBIGNN/8LmvKFQ0SQd8eDJzvYKQ7OZn03p63YGWEEmpX
mLQ0eeoQtYGcBCNdys9SGICKZZmL7889l3ljtug4rJilPhJFGoYq7WOEQugxUOwceg1dSEMsxTCG
dxa4WYEUOThMXxndCb15HmsE5n5xh1K7meYPXVTnJoCNzXFIiWlmwKkZeMsnk4KZnByeqEmY+u0N
SWuRAjyhd0/U4UvaYnypma8JQJfK7aO6OAtn//wkh9+PO07jil/YTRc1fcHYUClWIBQEZ1kQnWhK
21gFNlQlHJ4ItJhG8zQy5+eQ8ajrHovLP3v20SBs4MPdAhCpSHP8CAXK3nuHmhWIQvhhjSl+SM/A
LgHNW1cQXHt/WktSBc8WfgPLHOmIDRJs/2nCqamSMgqLGL8JmF5CbN5kWwPERlscn6fCcqX4MEXx
+wM0yv92sHFJ+MDJjFCutLMZJuQ2n+bTmqaDi4yuvC1AO74jF8LmwGZ4juGkWD6FXEA6G2b+adLG
JkiNsyIcIEpJteyGNXRJbdiF1qfHcqcTb/7gDQFg1zwB2v0JlIxuI0snMLfeyaAogKpFAOIFdIR8
soVyCIu1QTUYtqRDssY1Ny2LcCTjcPXP71Uhpc9vio/8k1UQggCFeQ/rnK1gncqGoG1OMXXYPiAo
fq6xnPqeDfPUHnLoK/sOddyDPmT/3MKrIsshoa8jxVMEj6g0wAYxhThZGvoy4Vag2PO0bTqRJVx8
q7LIbpvrwdx5ozoTEbhpSi7JG2PF/OFADPIxOGP44Be2RgFP13lFrxoTotRlLFr5JBvvIHFQhOtQ
fZa7bBGZ3HMdCaosuf3lhte3NCW5ql02sdkUkyPTfnFsNdY6W421AqFO/62sIjdB99PmK9s7KsSU
5nTQFzp8/UrlMn67PbEJP3o7dRlGiw8qFV7EyaRZYBePNN7FpGG/AeQ8JiD+8Q0PqcEHH/d/V1jB
kpBxVywxFu04C1ojxUHLpKOqF7+PMX8pCPvlEBt2uNfL91KgVw98renCrffy+l6alHZut88rItTy
qnCnh+RUCuUrdHXpO36fwkKnuAAI6JsQ7Eab6x6WIzW7IaPZEgf6/doDSAkzS4B1LOKbALWis57e
beiajWBTf1L5YavNFSFHig4xtnWjulw8Oo/0hmiSD49i5rcO8YUnJGBoMT4p/WGZxs51iTBnUlov
+EkXw7w4z9jpGopsxayZECDkX7V1wzcKbUXoSzfugQSkTXjkzIg7rEyA93pHsZ8cxbm6D2A5t4Le
mv+B2PLYxjWGwloIJ32L0I9geQBS5DUceQZNEDLQptqb6q9LxdvfjfvBPV1yxZUFwiA+qgFwoeQB
lMn7ZpVBENdeeJ/imTaMpVJyX+UNAqxLqo+JFknR0hnQujgeH1KFb1XwEKt9pcfMbtv1f6miW9P5
SaFUC16aPa0jXeOAG/8fXkjyoyfOmWFFbdtJDy01jrZo3KLSAD/+0QdFl84F8jlo71CxyeNqLaop
YNDeHKLHP/hwIcAOFW2kI33in/Xcmaem5fsYfAeSNdyS6QEJZo5On2poVaA2vgyeiVcf+tZGSQ6w
KcZ3LQhKYvh5H08/60Pirz35j0DiCGnml8ntXf0VzkoAFywnpkUvKOrs0KE313vigkbeEWgiuIIx
hjbWIRCDV9TAKwm4QnAxm3JJGooqeBlENCxdsnkru9P2CFk3T8ku/tlJASvGbWVNFaNTvy0N21NE
MbbPaoB953ZXE5SYy29HZjI/rFMuu05Ie5qW/E4dZXO6uv1BNKZhOLbdeY6iO5+q4p+04lxy01qq
Ihd5/1gAdkABcWAcKAnV+R9a+NnzZyyaYi/EmorxU9tpm8a5jCBG3eOz0klTYxrl7VbMff7ahPVf
bm5lRS4i3CojxDIHWuv05BDBiTb1893zQBlKRgu5eddekk/SGfjByd9AdXqFAcJSGMLYBlOh6/eD
2A/HLJoadfbOAQeoQc8masrQEgnAkA7GRYo3rflFjL7lff5eU49+0CDRgMQLQMPkR1UfB7iDMMz8
QP4v7acEI3tk6kmyxxesgVaLmZq7bCUDjXPuB7sR2o7dISXXA6MHeVgcCWbl3HbuwJf4UHHXvnHc
xs4fHPF3Y2aVuAgaRPvN87szDMA8MlvUCltvEEmCtA6RvZNpQw8p3eNTo7cBRrskg30SEDxRVZTG
zPVfLm82AzovAArL6/OdBtSYm5pjyznypYs97ZH7aDOXdBTRUTa6llS7gzt1eY6gYJMxZUxycUVd
EoAzZw/06aVvB47304cD6PRCvncDZ2nj+Je5BClsw8QfsHE3GbDonRp8aMBdR+WFDBHpWAqAvhGV
gDgC8Xe+6IyLBctjrgRhB5eMRDcCrtZsj6ewXqScwFuhxY2bZg8ttsJ2fu/kOBITuuzRaUBPQ7mr
UP1NZ+9VI/2q1+9pFmBj1ibT7s7b/DfoYcqdHHCXJsW0LcXtOCQGwYf/SdLQo3ToVzQPXIf6M92a
jnTNJzF8an24kDK1EQAAhjVXEBTlfp5cq3RzcwCK54xgzAjI5vv8ex3sENv5X7MSJqCigrNmk90x
hwkuiW897BM6echQnaRKrHQMYinf8uTbvd9UgnLcZWAHp2WPGZ8muXDXm5omgL3vCMtZaGyqqPAd
PwfriGKyHJLJfx5Z2AWOxwQgYOdm5sYDhEqWczKRpDzptnf5ALUWCqZlCuNk6OWkrQAKSJ7d/gV5
D/h26gfsKW2qU1/7cGITzNw/NyUnuEZUS7gpM84es+WQZjtFKL1AQacw5OIArGOwJjpN13TzjqCt
VpQ7xh4FkFCaueptR79GsnM6LKp6+NYtvUKTnDxfrci7SbD6c3SrPPTzDqY4VsubXe0GObq/bZh5
6I/GY8iWEzfZGH+WnatlwIW/icG+yjj80jEBSkKR80hH9Bv0H8KLmO5DPcdlAqYcQ0v5Gjzu5oyJ
tr6mSH0Hxf+tvjgsQZo1fL6Do3rNuwadgIlGYkqzsbobcs6Ez0PCoYEMHHlaSifkiy36nVtcZIwp
AEaY+/hgPcLpGY0Y7RsI2H+R3jrxN/tg/LqwJm22954agb6K+kAXAQp2iMxuQniNzvnLnrTYdRdu
jgOtL84CCpgTvaai+4etgP61RbhQNnpIhC5atSwEvOUA7VEQ6lqdXfki5mTbQIct+EHdbC5PvSs8
b7em1DJGxPM13OK/buWQ7JticyaIvZSaF3ahR/wNRsAwG78p+y4mAaBTlc9Q9IdqpNspap8yxsUb
6skNIW+VkNSgQ4RwktP0y8CBqfbyNiEuu6/REsT1hfbEV2RyydtzKk79qyrQegUKl5DS7TXIDRwT
UjKflnNCLshToQ5EJh+1A7jBY9UwJcBzT8c1NQ6if/bEJ/2RKLX1CyzMfau57usbodlrgW4Hjdh1
jdN0gOtohEGHmqlIXnjVRQK11igbkesSV3CMXY11Je9Dk7uI7ytOC8oNEJfo9lNISZbf9eGWL5wb
w73ZFpikfrZTs5jLDCjoB8v5cZZQetpgzxCkFNUOBLncHUqhruZFGSxcaoxtu1fbVChB+Idx9bDO
XYfXUrd5bDeTtnucAOuLfxDEXDCnkNcyr3zIbrsnBztPcYMrCBp9u0W4F73uB6KvL0V/Id30KdjJ
TFCGLEjB/rKlvOSJ2dNfnp46d8//LT3NTH6w8xyENcA3+iP7uIq96Bnajj4AsMdMMCiEO5U9/cy4
r8umPfqh0RRfZiSKk1G3YSlT6SvgLsj0DG2iv/mg+CaGG1kWBuKg/P2VPawADCG8qp9U3chjnBhe
DV4fE1u/onkxWtYyhoYIicoG4L+an5X8UEaTaVifiABu9LU8rNtjYIhmKDvRH5fhU2B2P1uFqDPg
6ya/OirLR6lt1bRKV6Z+ueViPHIeGpnDnKLo/SteeDPu8lytdjaEcCqId6VT2iIdWoUP3cgmvX1o
N9lDtzEluRCDH7lLu0WyxLnSHXl4kCJk46EKwxG9LeZWIzJwzpUGGpVplHNcyDaxkBMKAnAHqW3q
nueIjpo8ng4xuhKhsb/zVCzE6AU7mPHNGeff2HIKpG/HN3othJaKOLBgN3DQTM6QqATPzPMDS16K
zyzJ47+MgVjc5Ph5faMwQNv69KnT5KE2M9yo3k4OoaTVkl/9qr7jwcvwJkc5J1nPnRzg1VPVQi0P
uB2D/vAngjve0mABfenP/9PdrKM1X5Cp5c4OsllX1yJ7tV477eO4ecqdAjEV1EB0qILbaohyEEps
ahO+zt9fr4sCx+vHak7iQzBwElSBPPQLM/E4WQgr2w/Rl5LJhXnT8kZiDNX7IWXi3bZC09a9oQn3
mvrP8n/ULqLl5RBgXU8VFrDVKxjENBvNESh75/cmZtKmC5uO5fstWkNj7771XrLv/h/3nAbBmNrD
KyqVJCU/il6qqGBfPkhQAvl5YpCVdHM6EYPJE996B7Z/VQh3nPvsooXoPvh3HtXfihYyiR7Ktd57
uv/0tpvEgdEV0PXKFkR02Sd07yJNvMOicdxzFmi/5IhbC8cXs6udWmwx9FL00u/LSDxzstoxMPCb
L3MvtZ2n3HijAgItLgx6aOT9KfiA4kQZ3ui9tArp+KLRJrcOGjQKYBZEXqjnSli8ZzWrAooutG3K
pXras/w4VAtdcUuyFJuwE76lMhWu0QI2iiN4YlfygAZYRR+Uhe695iXSOVo9XB4d56mydHPqyAQC
eYy2UMaij9LS6a+sC+dranECOOIhH1LP0F8XM72h4aEjtaPbMAM5tda5wrHtsRdJD9N/GCsBmyv1
4cau4jCWZgnbBfXr0qTOWEcfPtHZsYtIpEwG7qyQeqR1hryXp5iCeUQjx5HUMDJMYbvv1EfpyEds
KHhOKS4UlYt+f/x7yHN7ILUFRRpdMYu5AnGihvld9rOpnbCLJWzMAcj4OkaCY+JaPvolB65pU73o
4D6piCVVTt8d0QAJZAVUHE/bOVaMFJaJd30k/3m2DupQlb2FAYoLP6LpWchAhyfQ356vGfRXk6h9
TbVaFmQimpeoLrll02oO9W/8hDennX/nGA7ZISTnDzQ3z8l76JyJpCNL3QcyW0AA2HNb2zaulDm+
3Xoo8gQMIqZzvjH8M3rb8JhHw5lCj9itpPglHbfa377Zf2aCpw8vxt4PcZFEXdsOz4lsI8v719UH
Cw69LWvDoLVPr32FOv3vGbaw58C92Yp53zLrOWf+Ob8Lmu2ZZQIE3mowboN1X14/z6mmrXqqxBxw
gBB3puDiDrKRZ4WdaC8I0xpjMCcVmNwYr3AKSt6Yn/w1nmzTtxdzSVwAAfAL1Y+ARFFEdPGfVlXJ
fYq2NiwbsYqa02LGelvfFPtIvAexYieh+dRUdWTKmru5Iwm5d+vBoRGpXC7Efvfmo/yYv420/qP6
xyU09Ejan66SmmlHml6V/RHQk0gWtWvntIkpESmoyxRx6NAonJqS8BdWamg3IsrQW0GwEIbBhokz
f5P9deVqr3p6/ReZVXL3GAN3JAOywu24tcCs/us4Ea6FKgr4w4sVCEgVlJbCXaifjyEzFGv3hlBv
vegjkF11XmS0EeolqxzyVxdvSx7+HOKxZAcK6VOXlQkFUyydaCnIcYyHrPj1cVGpm3zYlOykb7Py
I3IkgaQPfbHEue8WDXXIrX1rZBlab6pMxXW9BuHOb593MDA+AjT6kkOZkLUbgVijjN3yOXch4GSp
QOolzygTM3ioQ4A1JtY6SIahamUdIQMUKLXztog78zqHO9EBlgYGPNHh6Q08T3rsJ6H133breKfG
9TwF3PgAz49NR485dy4jq7E+9Q7f2NClt3sYxQ1lcsjZ80/rvSfb5PWfHY6UyXnUcZwQORJsmua2
CXiO7mkYihOGtXvHkxv6dRNZIhxzN+7M80Go5mXYRCUBT4I2PUf6TldZ5aEYuC1F0a9O9CPiTDtv
isryQa58L7Y2gfoy02B6RboCgeoUrDJuN3PWYYSokZCE8Ltvy7Q5Wc2FCo4kocQvFQTa8To1njU5
BUHA4YckGSB5MAV7OeOBAQ7kEkmMkT6k5W0mz+tGveOXvx8MsiE+hx+91CnBiXeKDTu/iCcmS6hG
CHRPgNVpeKqXyFN8hb9afcr2ACbuvxlJSwnGWjMfzCDr0Nd8bpeyYsvgEcxGBuBzSGjmes48vTwS
XR+M7pIpL0GUsfZuppoIKJm4us7XtoMbjWeNzSEH8TinbA+iPTt5vTjCBfhd3d7WmG6pVZcUn/Uc
ffmo+1qqvEhqpp+hw2B2v6n0muMqzY1JNWganBCaQBQgPLyJNpBO8E/fA7N1WB2TNZmNVtOp/jUX
IJAIVrrfMaEne83rNNSpS0X3O9E4tgmQxP0zLTIKQIW3445yDYqYl5dGwsHCScjQWG7JI9PjlxqX
ePnaRovAGlIMg2Cvc2qfgJQ490NWEzaoXf23sW7H1UoWVdGCfT6AOz7XyyKAksxjLXMWsekoXfdk
pycYL8xBTl35e4GdtPTmvmUzGDhtDcfLNiNiwBVdjD5rzJwziTCnFfYdwS7Hdkmg9++X0cCJvTyY
DaLqHKo1oJ/8wVDxnOWB6RZN9W415Zj1BBHmRkuUBz0IRtUj47XbVz1liKmJdkoqwWN+m7HGr8ND
wN6zWyVlVXxyp93ZCQyDoIm6VvgJ84wjk3ir+Efkob4UhvIekD+2gGhchlKLGEqWZFMRLtrs+mdu
frSDIKsN1QmJDIWZEh/J76fC/Oo1Z3mbMAABCERg98ankbAPWPp+tXUNmKTB7yqS49Nll9EPz662
TzdvaUX795ET0PzDFsFT+Mk5E/zjinkp+q8PdWjt+w1Gpc+CcwRmbzH4LRNsn19LKQ6+ow628rpE
FIqnI9lZFwCf44RXp6Em0v1ugG3vsqSq1p+FA5ahElnEJeISAmEBjiTOWYu5GgvHyVGRNMCTgmAo
gKR8z8MTCVnZMB5sZ1CXhsBu+7MZZdpTQd6vSba8KOPFOnK04FFzeq7jLpqpIt6AC+ZS2NGa6HIT
cXhmxbuTNUnZBB+iPxxfQaa2llYqdI/jGPx8LENs3b5/s+XGwbS6CPSoPbfHxbDfE9xgTEEspF1U
eyav7+rSoqG8h8yuBpIE7FnlmKhPS2O7wXK90lo7ZLcoUSJHc2iZMDCNuepAe1j0dOTecjpi75SJ
i/rbkH3cc7KHtFZMJAypEwS35er1eGjBHP/wnYcTmL+UAdCOzX/RYPSFT3eWEPKOIC2Z3aIn8BX6
UaE5/V5xYaKU9kdGwlmn2A5qaV84vMvNDcRgEnM+Q6v3SZNd7CYZ+HyG8LJhpq9/qBeSvDx9O0XL
D8ayih2m1nYbmaeK/4PfSO3kQbEUEiliVZLZlX6+L0vdUrNC+7U7VsBxeUPUM8OrT57Q3etcs2xd
zDrmDPA+v+M6VkG/yjQl+S3Db7Ve8jOMSRWhseBe9m5GgzVnfiCGF1mbbYY8ci/UaxhEIPMQQrlu
pNuO21g0D7o0XIbLPp7axko/E3bgSZqlGJhCR9emkFeW2yfVZ8UmMhHTvpItXzBNhDiuxiaV7MPi
WbuPs/D2Qal+hHvSxLye88EvsvhmXdP/oILP8X/dzKG7TwagFYFy6Jczg9cy+uxBVodtbciJtcvw
tQweUFqfspWNdIlxNQDJUlIcq89JM5Ig0fGvQvWuLKkl8uUKR/QqEn1utkHexCFZ2KB0kJqNUL7S
QrfuJ+a0SGlMd53d42MTI7/P8pOgKI/z1VZf2rj8vOFCivX/yOrg0VuYNOdtQglssXtNXBbQDzRb
7z7XBB+KxNbXmuoXsE2ZLCw84l8kH00/oGqr1LP6dOopGjRENSISOqHiEIR8Dr+rEwFBv5QUmTsX
Fzm7KC2xm+1xCKafI9a6lHKeq3s/7obvAPsDFtGjFTAHg7vXtuczriBwGpBY39X180vQ7ETrNDpq
jZhkqdFgDckGSehCf9gaUmzyILnMAtxZJDnYIpLMEc2YFxTRAl/T0JrvAI5PVtxwSaOSYYeHnfWm
xOzcx4YNQw6GwtUNr3pIJhBFilb7qEcybt/UEY5ckYIFyaGjY8Qn+6V/2U7bkMgTCAA05Ytj0XzV
uSsSvaLIUVLE25leRJAgYy7LwyNTF3KzJ8ifjdfQQ2zUjufzeDap4HJ4cms7zDcdFBzjER5MY7SO
sCQd+q3KerZ/GTPCBnKhS/o7f+BDWonB/SE1+JgN67mSVWyVaKFXQachE0YwVdjo5ITwS0Kj7B9j
GJhy3cQik7ntaCvc8qzu0upO8xKmG7XAg0hppihnfEQ0SLwbDsDuLlMToCpD3I1WGttQnsR4jjP4
oRrj/56b0WB+sSLJx4OVtwuVcddXvGuG/m3X9OoDI4fJl/xjKWBffjnNV45kXbWrApONs+J7uGp4
06Qr9NwtWdId37iLUxzJ63cH+BjxC5L7RBZOxfTtNYi0W2R7JY3ut2G8xKiGpisnPphK4X9p700C
dC+xOW+lX9LsqiaFNbrifaR1e6fOejtPls+cn64LjD/1R3FDNm4kI223P5vGt51qB9zMtDKVXSlN
mRtc9efnsULC669cQZUAuEqcFFU04X9zrKrcNAMOKGI+UK80/pEnxpDjPg0RND3nlkizPcMV+m65
UCh3o7YbtuFq8wnsTde7wE7IpbEUC4Ti+m2I1bvnTyN/dGThzUB7yGJ1dkjF8h1MTfU2vp+e5Paq
cQzPU60womPjir8Nku3jvQp0LelnVKuGQO0VU/pKILooI3HhEEWmhM8Hodn7eacG8MeyR7WNnt/O
dxi4uZQKD/Hni/dda2Z2fqpfF1CIfX1RNBnm0kakuAhmVhFQgPI2H5cCM0IRi/ginaE4A1U/8fRb
X/HguKkaBZROcDDH6apw7v92CX+QMmmujbRVTe2Q1RJBCjdszCUmpAxPyFEJ3A4z8GJ3LDOQifcj
VygrdYl1JKJ7nb9lkuPSicB7DC5TvQ3JQTs2PDouQ7wccdEwBE+qVSC2bj/tmyK1JkDm6NxSvaeb
tnfCJu8gJV8+ANE0/sQvOTejTWAlscTJpZ2c4OSIlDSjettgnHD5M3oi/ruUjclEyLd9L7BcABkF
FT9ppZ7aAG8/9B7qRNzUUhifNtGvyMrHVxvsi2N1CXo4NA8p7ARAOb9pFDJXdJwag0wZbhvk9Y/z
CwamH/om22tTgg14G1DTwjId7awa1JA+zEyfjhrCqc6ZJjmr5b8pWX/w6SIJ16wGQFHrZzx4p48T
q7Viduz3BANEeRd2mzzJ15VVNcma6ua0Kou8DBoAYtFKmRlFDUBCPL6X/oxbNB67JhcHbI+0g9Jy
8HpQMAoponPyYuuiLGxzSD6N/bc0kVrn5N6C+St+SMrbHZSvVeW/MsT/FV7T8aCD0WcofeFt7pmy
tP60Mzfg7c8X9xHGpTU/Ahy8iLuF5NLTDEE8fmq9vLaTrVl9GKmji020dLzyN9ORL+p5NoonvQTu
Zx3++N0AFwI1Czi+pU29IZxkYfAzNxd0XE1/FFGocCd2xZPVCRcS88dAhDfL70519c8R81VOkL+K
aX1YlAhEjZ1qztnWlQF0XG6aR3Cx9iiL7kxoPMeNRTtqTXdNZeO5RprnQQVzZyjNH3P8jQ91mdHq
IHTAuU/f2GEmwdUSXWL7Sm4598+DtZGDgctcRoP9+9ejwJBSSDjjvkwyvJMrdigXvaKP817MMW3Q
+KEa+S+tasZl2R72lJiIt549BSbDowgzO12tda5Fa6srcOpgE2N//R2j4ngv45W/NMr6AQKWpe4k
9VinjcMPNPdmfRMkFhEH8Reaa48+7w3wVMGsJpaxhDHqmTPqo4h0mx2nHsGKr8DqsEXj6n0AhUTS
XnPpFMUWK3TCBprBRi1ooK1gftinfeeh0WfFZGUQ5W40w/p4g5l3pliO7wM4lBdxSpagkWEjwfC9
oZgaftUYn2b2iouQ5QsL6jg2HENEJumZo36qhkx/AdOB+5pME/iLi90i1hOfmiNl7FToesltbt1b
wZ9SJDPjrMEjAinjjPIpogInTIQwqJHgTjYe1ErL6iT1GPv2ItdRyP2vHO7UNvza7761nqfV4OjB
LXXPD/bce0LH10QVUHxcSOHW7pSExnhQQeUKpSw7H0l9WAIg26iywB3QPUdPB6w459EwIl9rF4NE
fOeLIO0y0OCXyGIyWXggHTcoR7wQdlbEdF3gmAi1ZXeQm5eaItJcna64R8dCii1IBv/jmJl7XLnr
T4l7jqE9Pv4jPX8udqvTTkiCqkCMZHjB8WE727uET3iwNpSI5zZ6soSr26LGjt4dMC0N73NvwtR8
ZqWvm77X6LDN0VWqcIGWce6ETjyy/xS9KEtN1d8r9/DQesNSiSXh6l/QaIddPmbpoD+NbyRhPCl3
sII6L8DF9lwOkRZPF6jkTg0DGQXaMYUxF9KAs9wvY1tWLXvHdatsbtRDpdG8ORaKzYbN/uBE0K7X
tY01RcojO2UrVNEJwGoNkIKebQex8L948JtI/mkJcRImwABt6QwzzGPkF5hvEJHUuu5pMM6WpG5M
YqhKzqXDUJZ/GyUhBnuwhOTgklfO3mW0QCPxadUZr/2Aw+a1Bi/aTdPc9W15+6hO/9tb4n6yURri
VYGSZ6t9mvOIJa5doD/05kc//KCxNZ4XxfW6nT4TRDnxfUhC3U5vQ+PqBBfLSR2J18iQ0T6mXM9Y
qjXILKB6xx8xlliTa8PA2O0UWj6Rm1Quywob3Uwppw4p+QmWg8whFar2APTModQDlFOqAk9v4tlA
DbBtSu7eBHNhs83l9NqsJ1s+HFlEabJFOjkmGAs6hoOOd/eLGIf1KjymHeJl3ysiEt7tOI+dvaMs
MW3Phf5YKkJdrF8QMjWQmESDwOtkVBk9LmE10bpZ58nGlnFHr9J6hob0/MtOJoqT8WcdbHU3mwgt
NyAygDEYcOtb6tL/fWB3TSg6maha2vva6sGRyKAkNv2c1vq7lIfO+iZ31EG3jmNWy3Jj9rXP8l6x
DrQw8gyyE8+ObDHENYaZTuQcwYIBCgIqkZ0cDVsPejKG7nDd0YU0bC9XmU/bfACZQk4+kxnZJpiK
jqM/FKOpVD1RvQlfke9BXlJ5rKpyePgrqNeUbdnh3cD9CsduxbL8C7hteW6CS+pJzdIQRcS50COl
nV11p+nRDUb84VYNvfqko41m2J5ve/IBn72nvkltg7Qjy/5FKl7cs198AFZFB+mAIyQKMRvAVkw7
9QPAZDRpdm07LdMXJGv38v6A3UTk4zxaumXCf1AIM0xvOw5AcMFsU9Y6klV/Jm9+90EJJ2hgOI0/
pbaFMb9YYzwwWxcKM2i2NeE5UhQQgyOfC0v2UpLbBVDWMltnvoqS+Z7bLkJW/s2N5XniV+93Hj+1
fnEFNsYYOgwihIdaxGsbiAiyPGP3GVY0rRDq+RX2C8zi38zzz6LCkugxxKK58dfrgcTJuUGAjZH1
ODuD8PyQrNyV0xbR2VxzP/I2O84skXxO1vLreagHj5c1Cmc0ySolK3dKccyE52N+n/qdfQ0js5vz
SKqtvlDMN4Z1toUAOI+Q0BnpXD0IKKmFcWbt9JiUa15c/eicwRKUqsS7roSUXKw15dp65A3W7Q6O
kgfg0om2KN9AoqNUkpvIPhU7OK+a4odoIHPx5PLoHDwHDcwKptChCHxRLfngQlsNYWJUItAq4/oK
RNWOXxB8NCRl47JNxWyxOyFen7U3UzmGxGOwKh9ZLj8rxc+wvCBDjqLKjZrMbUpkj9T5hdSBORtk
HUaC2LNi/GjEuJkGTWVAh2tx0bxws84CuAZ+uH0GMrbHaocrmdGLYL30k7SFtZPs3759u3BHvwy/
8eXOEphqfH70w/VJ8BuXN014EIb5YXdPl3h6+P4gMlUZxyG1bhU7lsqMglHcai220i3xsEgL7MjJ
p3aYhXMQ3ga950xH5awxvYuzPaDyjrgKbL/gOaEq68I9nPSTd+hLKx6VWcNQsSiU82dK3a0obC2K
g9fC5QT1FpBnkXxvdnCm7EAgJ7O5jj/pIEHuMUYUwlt8xCEVm3w9zh4L+Yf9AcsPa0iMlXjx72Wl
xIXDKv23wJ7bTg87XYQALuIBolxOQuciHbdal6GRXPc/3VDZVc9Ss20FoWjHp330LLw2IU4rZWbh
dR0kysDhpihkSKw8CkhFgekS4Kvp1BohsS3uN1aHwimXEbm0771+Bry7DO6AGAOxSpY2oTS8GoEO
cTHz7PKsk+3w+79vjh9BBDeSOwgooxvJsp9w0hJWM3S0QAIEfXroD1ixwYc+38XKfA+tgqYupXzh
NyxzeNNp6O81CYZb0tLGwtI25GHjd44I5IdW/cYCtPa/RrSFN+z9A7ePFH+P0+OT8eEb9vp36x0a
9o+4RY/lPRzrHMLbL/8mkolf12/lH+JRkj+P3H8jMKgyid9DpKOlDOzd86sGY7fwlc6CvbMuLF8v
qbLvbkca0EGjGmw9qAcUK5VMQpAte4js6XSfXwOD92qTeIkB6efA1ZKrhviSLxjvDbQSCA2usuuh
FlZ0uf1LUIGUxDYhWiHXcBn3RHGTLsXcTy49q3Sj7OxVXKArUUAWHUoN/bbiaNPQw0gcLZcJiAb9
Q9eGa9XrcV7f6rIFNbXSg/vnGXIoZilPjzW5kRWKJ326fRmkTIq1/FPVXkHpLDCYIcdaKR9xWpj3
GgdROyF886LxrBjY90MVGuMjuUyHURVs6Eiw1o0C0bPthYSQQYRS1ktMGfWWhw1wPTkhsxhfrd0p
XlWd7dJNoDc3PIWeTE/YULmR0Stl19PyxhQqLz7uRnl1Y9XehJLzp8CJTmxmjoFE5YtLtwzJCZuj
KmdcuCE0hHhoa0TiRLKcPGM/K3FycawI1X4GHiB33dkzBq5XtKRldnj3PoeyFPdc1TiitZ4J7Kab
piYaFIyqkued3M6Fa4I8Pnxg2S+kmQlexcpDb0xEedRoBlplaPHIDVD7QvTqJCR0RCenAdT4r6kn
f1cTkSUQoMbfSPSDLIBsnwKTO7R+OpuQu++brlq4He+cnIii33msmX1dLrgK+V5XwL4xEhkmVo6U
A4RL2sdM487JrK+En43ccXJhly2zLp/qSG6JpHbW2iXoc9gDNmEVkhJ2iPEqzs/ogCQfYMY/AVQ3
fBnHXT3zpqwT0pRNuYaaDBogQ0v7mJX4igneTWryg3QyzdpWESeKjpldhsH+elLpxmTri8EvFbO4
yn79wYhK5zrh/RByicdb+SZGMBxP4hLfgoz/Nj/hMb3PaOJldNbQ4y24/erTk+JKEw3v7OhMYpV3
dXUX40gO5e5ccOX9+WC2IFWZijT1LaHaxEUPm9yXcIlwFQqf6k89l6cvjQebrmNeBIejsIBHw3QA
8nOyuCxB7kPFcOlKmo4ZQ1xQKA5LGAFGorXH76a40lnIEhzF2TvuF2lsZc/p8ZXu8ucfy3bt9K+o
8w/usH7TxTc1o99rnSCcwXqZi9cZj6hUIdElaVlB7IolXEcpomnmAl5NFsx9t7fAplyKuCBG0WzK
buRUqnzmiyNy7bXmUPRjv9doUeQHpM8EJXPLBexXGe6bNCVr8NLs5dHggyAEwXbZeZlXnzBmlM0k
HGWpp5bQHj/6S8PlriDvlUKDs70zt3CYBTcRPyyBpP+euhDjtflb7PhBE2w+zBHVwUkhKhcxYpXl
lbo+tQU8NrZNPKgbHfsPm9w1ziq/ymtfbvPptkuB5McOcKnS/guSsCzh2AmvqRc2niH3KffrxR5Y
w3lWIk0jagiCrvm9Jyl1wUt6cGLO1Sfvy8BYeZLRPioPUmpI/HVIqXbQSYC/tz8367CjbsQPeX+w
xwll7UtM2VYeE0kEPYdj2M+L2emy5edea+AJWNTkwz5yCGZEG5yJj5L4JBQuXNllOZKAqlynYwts
aEvh3eHnggUzGUVSAMg8LsrNdjKrJhyH/HFykXgHdMM6ghL3ruINWD1U3pRk8cO/j47jqKQhgGtX
vr6uRG9ioJp35UMpvo95ZRWOxokLCZJEoEA2H10NS1b9Ijnrie8T9ejAuc8PNCkfez7SI00xTmKt
5oe2H/NBRL80YkGAXw6vMwlfSIAsQamqPI8ISt9AMWyp6xq0ftEeoZh6Czpe4xGTmLk1CPh2Ud9l
WEfCBiCrIzBho4tEdFhwGyXyzgjYWufq3/d4iQNO08DXMzlUdOKtOVKJdq6JFgjqoHGCscLxiiJx
YPqiV4dnriJmLlrUZZ1wEOAqtalQth4dcZn4lef2GFNaIab5rJVzBoQX1/7T7wLlaADUDjKESyLG
qyPMGrnYhMWrBEfT057ZS3wP56SlW/IlfTtbc4W+hSDDCRyX/NhZRmDwm536CclS8P3qLp1hZfom
AH5BkGraxUVfLlgRvmKJuWYmuQVnYpR8h223mQzIQfYYaxjtu3p+Oe8wErZCPpvSvVaOG8KWyBYi
j5pC2fJFYGxkVLqqoAvP0GPlYngUPh/TnBYgt18O8kzNLNATuS7WRBVrBeWt03DYldW1eGMgpvhf
WKUVspuPB6zsMOfHV62/ou3nwiGokm2lMtfLW3TCosPEL4yULDqNXZp4q7Ea9hO3rZhF9aLt/Ds2
A0o6NSRkMPWxo2BCE6UyMwSvWrOwwgQ0lioWawui6HXvWsbypJTaPt8lgCTUkkzjlEWDzZjXbK9n
ozqO/BoedWDG7DKVDXrl61mfSsWBVpmYCcjvQMahCNGgMZlcOYsxoIFYzWe8+kF+2vpqrUVO8nRA
AZTNXxZl2tKhn5tex3ylvXjsmnRrSD/e6pWn2l81JTMbkl32ECqn9g2zhCEPRN6WDYzUWan0jvuy
UDgj1yzt/FlVAXZM8SXF2DfVl1OU30ykcWZw66LwAGAH3zDoVKWKsyrafnD1ulKSiwZEAk/X0E8K
qK/r5Ix/niH9jdpHNyGAnlUA4wyMaA/9yXdOva9k6foB0XsS8wTCh2qf7zxWQKfFQSDx8ZHu6TF4
Em3d2Owa/ROJKSDJmnFlXHIAo7BlF9GgNR098V+BLaJx05M1sAs9BR34i4EruvwXcD57P1tJpV31
0fYZOMBzybWlIrnE0hokgOPnJNIoJnLy6M3gtKEbxTvrWFWKEIcr9Gv/GKFkRraMc87DRTJAGpXc
nRIvtteMYBFVETouZM5pdNPgvX6w/kLuw6kfciiK9gglCRw40fs8IDUuKEUtUFVJzqXx9OMfQ3/F
gJ6/+7Tbo5r3EYVJrpwndopRDU/mfWfCKwOWvMUyQ2W/hUa5Fpipvr5S0uMLgUA/435knwkkq7/c
Bgd7MH1/Agh/NZJ1d6SzFxfZoNqIXDfvJ+um396L0rPBENDOMkw/oGiywvvZXikQlwOrrzzqrVwx
FaD+nwEiFSNHKrsN8p8SUm6FOshFgirdOVT4ZcAwrNSJGTihOWtunSGwuvZ15+hAdHzItyiXAzKs
2OUKu1w9ve+m9fhq73OymfYervH/gmT0sUxN8yTR7goMGW3npa6lj+9fryfTCCKBhk1FGP2E9H8+
Y26PNpHwO7PY1vfgCoShiI/1O9Bi6kIwd1IfbdehhSSumq91s4b8ywzvPWV2flVZsZkVl/6FLhe6
0UqsWUKXdfHdSza0IUnh8y4W6oDZD2LQ+Ngi1rHhYsRZ6nWb+LYJYtpP6Ge6oRPtcJ2yxwPcnttK
DiHHrzF8zugwk6kuFH7QAwoo6qs5RfkzE5DfOGvEkESCBkadO3WPe6sVOpPexBYZZiWfKJFAYTQG
8lG00sKw+y3Jgr4BO8xAt4owVfjx//MxQ4Qs5oK2HH5Iq3EQyUhy1ZywYhJZC+siZMN1C0YDT5VN
EvjtMnCQHjojaEJGf+w93DFkZRBENvfxlGC9Xi5aTKXptMGzUlTPpfwVXzGFsPrWpNypVa68ia3B
SEcaq9qJDtIHv4U7EJ2FcbFEi62AlgObNbsRJ+F+8puK7SKTU8CkM32OpipYQTY0R32AntK5gf7D
w3n6bTgWNluEvmynb6rjjyzGvLcRQ6X5iLtmNb4lHAGglAoQiscsc+aT7O+EI8a8sdYGVkmBJMq4
cFKKK26UM0XqDR09GuurQrpX7D2tpCg3Aawhm60a4lHmcQXLis5j0oNA4xYfNVcjMyN9sE5o4Vkl
qggOF6TA+Cz3MEiBSfpWQHtIV+T/RyMPaFF6YB1b9w67afRGhbA+k/i8+tLHUuBhdyTs+TG4uTwr
h/Pog47529deA4klg1WosbMynKBF4AGeId0RqkP7pfT2+QfTyFtgGiQzdCRJ55WcAUOe6Z8mXlyt
uLgwR38XdSnWsHMKrkGVfcZjgNEUEIQv4HKfqRPgghKqy2cggKJa4U51xUogMrYB0nyask4xiZga
GIEniR9OskDYzUJc4J30HFMZOohL372IBdALZZHCTpdVa2kMnIgrYC9K5wOQ1PzdhExFbsKlbrZV
Mz+jh7X76Xf+JnAFICOlY41WGz6ezzKPi5nCfvi2Fh/fTBKNs3QmhRGQp103GGCSSQDheteNULyH
yj73zVZFHgkFc8rWhf5N5kGx3Op0ylgikwvAqSdSsjEwhVZ5fZ8fijk/9Y+/YKoP1KymDO7Z+yCR
rZgGbhnTQwYM+h3atG7HkUp2Tu6dDKlppEUrqiZCPz7/7UBdctX2qkum3OaFXHH6wis3t93xUPpa
X+c0Eh0LtgqaymM+1chY1zI1qAbeNF9ItDiqNGI3RwIUacK2qngGRSCaM/E8a3WC6GEWRqAGRsyf
2kVTRkbhjSM8Zp8gheuYCXzKYn+cSb4VDctXK3jVQfjYwNCF2HtZk77uCS2SyhVPPyiemCwHKamH
s1umz6USUcVzO3q7/U5ZnAk6TQAsA+5l9fC5+9SGe7ESJaP96rGH944HX02dUtTM8h/MzjbmtTH9
//HXFTXxm7PaGZRE+3PNQJLds+bDx0zEZRifoAThOpUmJqnCSuhdRjhV9WWLIeQJQ6HvofqLLUlN
7FKt+uZ+Tv3fmSiSWQx/JN/WjydZruw9JP6nslULIGFZcJjaW2LcneS88q/X4xi1uL89MNNo8XF5
24xfR18gjhoVir2324TiBY5sJO070RWX6uPo9QDylVqkjTuAxvjSmuw++kcBdGeMVFL8uJQSHMX2
9Ki4kqCjRCqHQWcgKsbAMpsiUGvvZN3ikzEZwS+BWJAme0o9iI12+tSYIPHalXEhm4jQTNFdmubp
qtvlNBI8wjf+T9cdnQXT0pYEniKJUEU6XuuhhQ8eZddiCULVOsCVBxP4leBeGs3RnWcouVOuynok
QUzZwLa5cV5Ihq6T8BWhMNZuT5MNYa63bxyJa9BiCag4WXUzAjOmGVFyd/CKt4iJbNobS9pnlI4P
fLrrpnkO4jLtSYVTEvCpu6BSPPq6bR6KhMMfTD2rrcRuITuvIElzdqhf1QNESVX9htYS+6ov05by
i1TwShqOZ7FkpJYa/X2zuwDVCzDs/Wl3M9B16MPYZwZDUXtQO8apYEwWFeeAYbhNXI3MlzydNFXQ
uNxrAi20+DKcnVUpT/l9UT36M2ogPKi/co6m0kI2SQJb+Gq3b7Gcrm8Z8utZoCNGRdNrUyklAFlW
zuoGH7TcdkZkrFBoHFO8IB/bmdZfP+8rinWQHoujmZBDx8qHV32IRwpItO8gHhG/a+TCX0XCMTfR
PipKQSJQJ8U4qaLZq+QR1lSlusb2kEoyVqbbwrjiFqodU0d7q388pKpUl2WEEpkSKi9a7c4djpsw
OsaFDpkF/0e+6/bC7MSzNt7ecPKf+wCaMTyyYZ4W9NyHiBW/GvqIg9Z2W4kqJnlPQcNiVLk7IdPw
ICO946qG2FdogdzRJYTZnZlw1UwrcEuU8MoIA//yIQruvsv3ncDt+DOQkNHug7BtzF4GaL/59xA5
kv1cPLPS8drE4NPzsuacTJx500gCokrhu2Gq5kiK08tLDgMqbJtBjRWJFsMzyeQTrk0G4xsBc8B6
Rjkf7LTBzGs5SKvqpMXXKfbNTqG4/2I+wBHum9Ff4aInI7CQsmPLNKtBD5kDWcmaj21R/gLpywyF
IkEVyVe5kzK9pVkCqBlCeXjXP0a77cSveiu50vbxvKxHLhXGERmytkToW0CXAPoLoL5PveYYtrYB
T+tOPPbN8Hg6VLeg49SNdbLSbfqR953w0Ry/byof9iwYYMfA1rEG4tYZ152bq3J2p+enY7k76js7
nXXiedO+ax98LPZ0ZpEeWmWNdeeyEzBLezp4AzPKlkahuwuu/k+NGm1C672ukJt/uz/e0aHOjrfH
dCeYkP+/2xnbD6Kgk+O7MnDmQaLtUKgx/QPZaB4zmvXL0AW6U6gsPWXjRNdCy+zkFSkP+hH2Fty3
ZpL+ILnjZVHYw80hvNLSpR2j2MVVG/WF+h/UayQY1OygoRajx5pI15Qa/JwjA3cE0ihr6Di3FB7b
029jDaarQGcUZk6vs/zWxGP9Ob7nk5ZqgxKLtkfyAVyAXHOxER9qTrSBSXG78YDYOJwSbxlvDjDi
b69xQrXOxmcPnJxnXv7ih1IgtX8b6zPsz6KV4pG8KFQF+wOjRcFlQVNeS6dJRpAEuB9SOjt6F0jx
5SVDsXdEg2P8yGtmt+utffhEgkM2cHNHUYszND7spWLd4KRFyroko9SPMJC6ZBQz6UBCZi4kNIDg
EpbcxpRXHVJYr/OmYIwt6vQMlcLpLtD2D+/2XgN2tykbSYAc7Nq4kVcRz6xJgBOEk8B1aJIIr7qR
uaXR6ZaAAhH55U6aKIH0xk6yxGuqVT8qDvdMQ1sQQ6JoiORgkKwwLPdGrfutZbWBx3oESzPEFwZG
plVj2WRYLkZ6qAstTcR1SDYeskKYLaxrrjetuOCGOoNUHmIworrVP4lbTCcx4e8SHlK4DxvToe2n
MM+jGFsx9Z0O2sGK4hY3ffSZeglL5ssFDXjlRZk1jFa2H26jHgwH0iU6wjHT2t9DjalHSUDDJ6g0
ugqnc/YKpkV1v7PSDEBPIf/LbxjQuxIzCKx8zIZoa3kmDwnQHuKRsWzg64u8zfrprn4OierhKX1u
ghn5cKdXyFKZtMf+kAEJlsBzgoONcVf2WFBeZVZSqA/7PsBsTTpgx8ok7kz97Gfqypx6ZSUxtqlJ
NjCGtQs9Tfjvm0AnG6hhI+RBQBanq9ZrsCH3b12srUwEooLFApUPzCUoW0wSwVEXP7g9Wy4dG2Wf
80j5Zs/WuUdt41TbMuD90hdJPX0wevDjfz4/oQyJBkNmtsAXHbaydcIZDwxZpvkDaPTq0TebSEwC
BJxluhJZuaQ6cNcz5mFq9M9x2CHQjTzUKDgXUpKRVBhDS7UPFl5uKMcHm36eGaaodQ6pcNXX1Lt5
BTUmCN5HfFfsrqGNNKOei//NnIRtFp2T7VKSoTLrcx1npqRiLTtA1D4esgEYEavxGjUJ//zg2UHP
6IulTJFwvxgbFi7iJcksgTEvNJaApU6893BeTUJ8AuTbNz/9XrqxOeOfjZyCDQJwmjARGLqsyBYg
2G5tNTbBfiDZi9Beg+PNXvIyMJKXFE0S0p+QMyBvts8R9L6WF1TTGEBBYhjuTh4U/SovR1fq0Ite
a+CvJH3B0YrRiDPGT/OMYXa5ym6iSkNZ56M138/Ae+xok5dh8T0vMmlidCmcipgW03dGxwBYLo43
woLuR6lDBFV9da8LlDCGJVaKpy0OD92Stt4C/BmAZgCN6ORkB3RtE4pu+XVBuDCYJkQGvU/HOI7j
G42BVj2aV1PKAM0cDXmcsjlqDgPvfKF+dkF3pXdO/ERN7sGZdI8PXRlX2q33CoDfYAPbf2XZDMJN
fSvTBVI2Bk36GG8Cdox4fi+ABqHnlDF6qGhuTO57/iKvFkoogopgfzWX7Mg72o+yS4gN4QvChKn/
DMxoWD/i+wAx53su2JC71Kz0D11fs9SF2Z6kQEJAvtXMFOUNCxfb6PCzbqGiptwa+ivgw+RMbRqd
hkzFbLAnzVUQNLrRLx3hEoiDTvAUQkotm54qeBfORSzlv0o8CKwyN9HDrqt/Y3s6OrGuEHLTurSg
p6eMAairXVFO1PLBtOE9e9nJmxPltElGsa2p03nIksP+inQjOgZmDDbmLitCgmEpfkpj8Fnoc+IM
2M0vzI8iSvqRu0XFUEO+ft4VMZ+J1Z9P4vPQFKuw+GHRDXK8Dgoj5Ew41+kPdG4egmmLMeELZqxO
ttij7oP2t6cC1c7XdMj+48L07YEn3axaEdt4cwLHBCQyO/CXQKQo9LzsDy3EbPNappa4l7tuWeaj
qgTgcbpMlJQBDOBWLd4I0Lpy8PRTHbh7YMKTbcYVpckBRU08ar4/bBQ5CA4xBY6oe20HsG9/0+aS
/u6apCamhHj0/0hbKWz0iH3WRRKs8fFKm2Iw90YSs3uIWETQIEDVgkyx81oQK7YLJGMHVP+VzXI7
AYVyQ59nopo+Oy2KoSOoPYmCFizu957d5WyIyikr0by/qst7U1te+9F8wwWQiwiS4fpHlTUguCHC
5xE8hImTfcoYhSAQOKpgUnqrE1NmEgI+aWhPKNl2uQxb7/CpP3p4Zhs9CtRGTXadqJ+bpOEUV1yF
0YVri7a6hKhumkRYvUzxs0CHvR7W8gZSRhrcG/eTtuYeeYgANeEL7F3u1uHLKz7XlpVQIGL91H2T
Hj8oVyFsYc+TbTpBufwcyp1JNSE2M6ZPpW9X1JbeDvpdzS/k0qVh2IsSX7kJGhTTZcGQ0Hy2t4h4
8V7w2VqRJaQYuDk3/a7BsJTlvi6lrebBHY9ghyVZoDzm37ayVAIX5gwZpZPBkWgsMIrFUjeJwTMA
dhQtT672AvA6K8PwQPIBsKUJbTsWtkTJHcA8k0gVw/oAoDvFrorDl4a8wFGuCJoITqvEZ2Z/4OvB
IkRKbhKj5U8p9vmt9LrD24u9FKKfROJxy+KmP0srtS/sqRnbEEARGCcgUyYuSU2GfRDKS8zDZ3TO
vgBp1tRBPrSedfDzRf51flmULP+XAHU24UCi1AKzVOD7u5ssI1Hn+QVIUiJJ/DcmCS2NOvJTav36
CMUrgDy7BKhD7BGqkCK5R8Ybzl/XLN88vXwA72EF8ONA7SH+IgVNuKUbROJe3+BHO81+aKWcAp2y
FjpfReJ/uQr5q8hzIGXrEWGbdgcgiyPesE6qvBsaukdfp4QuRtwhSWKjUVIHo3xaMyZsK7JhA1FY
bR0iA6GfsHJa4fIMU7w4XXDtseVCK/7SYpdLh+8tMtaXGiK8IBNTd5akJHaf0JzmjxuMF8FtavHM
b5vLwt8djfzcgwcTWLm7PjnHHDdLbVt2/h52hG0oPvCsyx+u1ZbrItCEAIpN8Od16qbBlHYYTkVa
yJSpkX7GZ8ho33ReNmOp/j6Mk+DF01TLl5R73cx5E0/ZYc93d8+r7yQjx0PWDx+roqSL18izwSq1
QQKYbhSRHQdFzoQyX61okUVE1iAJcVGyUgYb6E8wZcc6ul3TBwlvtag724v4LZRd5TRWxfI8c/0z
zVUF/zsCxWMgnrOvnXWkmhRANCsL3Udeic0kUOoiWRxNfP5VKdKb+r7tC/W+q9lh2rvG1b3F8OAB
d83oMFhrYW7HDgXU5nuOWXJUr1d03DFQMGJqTwda4vrQWO/2k4U3IpRZjDP8YDZ+jBp+Lmx/sMsX
DgZ8+nDZVuJYr5Uu7tUrFKjsFLqWX+VbeRWPBmp8tFnUwa1w/zPyV8GwPNzwpFdqOjz5zAF0++IW
DyAQGU1NK/oDIZqsOLshriEVUG9iJGO1ng29DvHxt1Fh3gnHkT0SXJxGnIexqacs3NFNPz83xtAO
PgVdDw77RguNod/lg5HX4RB/Dsjp6tJcpKkD/fHk8akA+Zn/mdm8V8RDCbJc+t8vf5k7WH7dCTD+
6zKPj0FH8U0aPrGJKpiwUEPt4kbnzBVQ+WcjUmZiID4dtmPpdzq14H0cv0TGmLJMxd+SIq2H4wyz
7Shj+6ZCESBHV8BfVV3sty5gB+bQEAK0COxmGMzGEnB76SSOgaKg3EdtUsaa6+YzfBVQPRPPBjnO
Qdz2r3PbCHep7upWCMeAJ10lci4m7j8klxHmjfJTG+OlYiBMT4naouH3ouvdKfroHdfzPeUJGvj2
4mt434oIijXiDEmY8OG2qSoZ0qaclxnMAitL+1wBGNCHFHfnk8sD9yMVX6g7pswcLJOvF1H1iRJB
qcjqHtgw1L8MnivSdEPkcAYpxquYhRDWxYFjxi9a3iQBqt7V24szTjpMC+LRjBkdDF2NwtEECl5T
W46vXz5Dsg0u4jBNbZJ+gqyQLrBQxd3exDBZmztt4hpV+q1Zvzjv6VwtEQcQVxq5iaahv4riE5YT
odmeK5uuC6SSIHmyuKwEwvOp8M1KJXa0L8qc21HxKe2oRWvdA0as/RuU5JnAsOx2QcxTJF6N7bvu
tVs0eD82l5PgxHEA7Wbljz/ofnwM/CIFpkd4QiYJnmyD0at1cEQfMQwwscQJ7Bz79V9rFNrC668c
oRopbrQtwFFYT/zwV2F9b9yYYVn6tupYwatRFm6DbwWb1aFY4+aXtjPAGg9HwqJnLVOJPsw/x140
KvF9epi8TI3AK/a5ybdciuSVKdq9nbXahol8zYyusuClf7RpF9eiIMUdlJPYNp+fdQbynDAGrSTI
T07F8yJpmw3Vbd/49Q5dId55YwqHY1I0lY3hyh5zWTUZprDbliULMjVX4MMI1Q0fZGEGWYQI9QDZ
LKstulISI22MSLcciGetYHdOF3mIEDG06NI5AcpCL0z71AFlVWPLIvg3hhCWaw3VS22BG6dWeiHE
+0V0M9xNBbjbQIR4sPNObIu6hUtMZ6KrRfNTplR5wjRQXlJIIaKwb1FkTEAHxuyHgucbp6TdKfoQ
RAW4KoIPXHWC3U4NnapFUnXYROSaTR+9nqqSJU1x0syE7Th5br9q8pCnQklZompcld26GFKzDWG1
Iy+5zxHVTBJxl5dZ6YckvPLF6aN1ok8FcIQ1k17+pQAIf5WRiaK1jRNjkQf5cFawV0a9tV1O5zo8
n7xI+9YQkD5vpJZRcA620nH8e0qHGQSPyiXcxSD5Kk6Appi81W2EdPp0EGIQlnohxQpNcQiaDWYS
AqzaCf0xuiPUBF0xbxNQJhXS3PAFqTiTGv6GTlxvIYrEQ9xzX986cxTrASVmMtjsRV9YoBKSCOKA
Vsj5qojbQD2m0Gyb2jxp1cm97EdpowsiwMU0i+Df5RVKf8jigY01acSTkma4Rwr1sm2Zs8QOdwtN
htIuxExawnFWNT0wGZ/OW4RP2nfh0fWhERcf5rD7tDG3oY8m6FTTP/D4a7wey8fyncrpofRpe2tW
QuuWCT8DEpCKHd/6cB1GnTmX51qpm5I1LmQeK4xAMXRJYPi5B92hw637ndIyWyh1Bn2WXwSJhiUI
kLmEEJPARMm1x6ixCRuXAdXWtQESYtXXmE6Zcd5vdaO0JVXeWmxSINTj56kgiMyGe45xw0y9tn/1
7+msDMa+NKkAQeN6rxKFzmafxuRuJlqj3skfUOoxwFzICFld3cSkgonVViKu5XLdRj1NBkFCdfR5
/HLurLtU/GUBwlFlXfLl1Ja3GHTq7HNPggRs5bYuFT/ieVFhyt8oDdwXeJIYV6OuMYaddu4wjGmZ
BESQZPgrxpCM48+ipc3VbKm/How45mqloQhtpfh9wN3/v9hYKHIlmPHVRoXsS1CF03Mx6uVAgRTO
1AeF2pv/jGzZU/ErDjkklaB+NfkhZlwWO287jWDm5yR0AOHIBFKxBZV2ePvx2nUhEFVikwkt4A+p
Q5wDqwtzuVhdoic9N0EiVZLLTHIazR0WlPUsJ/Pl/gAhdyV3uYQ34CVP57el/W0+8tqhkrS1rtRU
QGtsLveXxbjzVjbXGlKySE5fyqaM1dlSZi914yRIfqkwFDZcD4O8tTTsh5aigo8YwfJAjibgUzQe
jYeZG9hYHjtCx/lo1/8pt9TrUCW0eSF2JVQbG3CM6JJgZEUIdfMnrWA4Cijla7ZjPizfWLyBiN9e
cHWGs3SI1+bJLjgnFkATd3bfQYRWtdworcny3uoZnP5XLsc72MwGV4IEEisI/k8XHF7AIXm/bxtj
2pyeoQkZuuxS6UlhMM6CJlI+E+3vUx2ck0GPsVXFhzAqBWa+RkbwCwHKPT0J1cvFBrfFB1PAIG6u
/DzKW+SaRT9a5F0p9653+FHbyu0TKl3jDbUdQT/3pyGC2exiyIGiQKBKYx4BWdt8b5OxGm1VYc0j
JZ5+lUF7GmJFTz52/9zo6g7bpxFUwOZXwUwLb3Aw0uwsGUoy5U5KHKEzZk8dt0HjigthA0e+tbxE
67B6bUfwmLD0gYm6vGAtkiHnS1S8t3S8uOyncsJ0eAkrvuaY1Q/5DzLtsyohJ0yM/WLWq4evFmSD
5hFKCDHybmDpl4SJZ9PAukA53pwOK1nAJeNNIsIZiAAze2pUlpEVOz+Ruc/btw9PJXF+DBqbr7Pq
DuFqAxDKMFEPmUKDi5D9tmSpJdD7Kv0vUTPFHdUnxmbqbkA5EbzQcJyAdF0Cy7FznMO8nJ+NKIon
Gy/gJQrtzmk96SToGKIesdBwy608FQ1h94/hvQxPM6NoxsWSiyhxr7Vlixx0TTHPYwMMfoP7J/S3
9fh4F3H+qDO8PDL9I9dhg8+bMiurEs8mHjW42jwqN9NSD7s/u6+BNvCCqSjY4zZ47GvuGh39gko6
ldq5/i9DNh3lV9e9uUnLESta/ihoXZvMfLQB8s9YBToMySGVk2LDHe5EKGilZcI6MCx1w881bP/Y
UQncQbi3FZRlPcvyQSymsExNrT7vHWT0NzAWjHna4+ID00zu2c+7YxhAxXYkYcSxqFxBdTWgX+Mi
oYREBy6RJnPT30SQRgTn/axzAcLA6wE6O0IjSVcrIflHudxYa5UzxBeJjjhIbSqtjGWlVDq/nxlj
p7qT5L4g3wqkmyUrCuZ8nTbRB7z64jCPN6+UhiB7ZwQ1fjAHxRJiyHm+YotPB1Ctq964sm8pFe0a
qz4x8TwDMwCzKuhOINZ55mJZq1kCovMgzv9R6xNzpdHgD+K2B2pfYx3Wr2u7BXnyDonESnC0ocq7
zR8E1ERWP9Spd9TnCIq4dUDq50wDLMyHDTIaEycUyjDHHad5370vxmsIZ5nHy+fXM81FhuW1C3U2
0snK8FkMMaFhjxKHfQI2rmWrRgRApG5Qd3VOTQOvv4EnI14tIynIdCpBK250ZLp710lfVzUCstI9
wqlvEkyN2hyemYF2xeZkF4VB0fDJinG8vG7USAqqqczhk06HcsKloOIsDPb0qd0J9e24eq8x/hVm
PxV74UYEC8BHzXQqfoJIQl1cN1ngYG+wGw4g4udOZNkZdDFwmd7DqdyI3jgVZw/y7Dvtk6er1GPC
PBJFeSWcAc+E/2aKuEWADQJVeT083V3AE28XXgjl+ENiFNvECkMfAm5nxq9Gqr/htVpUS2IGqD6d
D9NVDG8w3OefDfiXlb186ZwXmmqPzhknnGuGNLvrbUPbhFNVt6efqAjwUT+DsYj8C1Man9L8CGUJ
Nr3PCctQctwlU0u5CudLNzL2tqI8rE3ksTcRKkUHNZc18tBOZDIPRsSouRh4icm2n/dWzk4ZVDFJ
egQ0RERyLadMPYWQ4/ci3n3Q/saq4gVyjO1PVHaDTTG/SG8fkHxVtzLNJs+6LMonVqUlAXXIL/31
Bq/wumfDwgrwcIi15+EqArg9U8AfjuvSKnO23J6+FYmQsr1zQhlkb27wzNd7NxSMipq6d7+nm76L
+Po2c5Zqx73L/858CgufCav5HMenuR/KQZ+19YUWq89jqJ/wkRyIwCpgm6s2RgPOSyKbHWTky4y+
OGwoR89c3tey2BphzO/aQrhwOOPwNilyOgZxO9GP5c/7Rxi/EoWNUbf1K+2Std7BANXwMRHwRoKV
6CnUUCxT9TTNnBVbMEmVHsQ5QsojhhpKxzI9DIHLZSz8HMD1KDpxvTR3EpE/46Sw7RG5iS/7uEtm
PgqeGTtPl5SHDd7umrIQa3HoLS7VxDZKm3/JTrw8mVMSAV0RisJueQEZItRdJ1JAlutFnAuIMxEw
GT7HcQsKJPnqs2N+ZFBtILK7Q0MlUi7InvjMgoM+e+h3OvSGvtHncslskZHzNPMH2mevJw1Z8Hy8
aNYHO1Z3QK+9f+Xg7nNFk2LXs/BIbLlpBvcqelCvIZKFFwvg7Z0k+LW8OZOWr0Z8D6ly3Eeaq43X
9p0LJE7ayDoTIAJmoY+JrP6Frl8unzbPg5xKMlFsZh8RSsa8/cpwV6zGArHnvM4ae5/W+D0Mf4LC
yQIjRbsSZ54HBgRulpF4O1NI9F/5n3homJyi1NhzD8FzSCs+CnZ20rqyDS6+/TmEJ7XenQJo/jiD
Ua1ICbVY8SgKjMmZUvMyaj8eUZ0hJNgSk3VMNV8cBEVoLHJQKVMJAcrrvUta7/3X8XXgGKnq9hCb
k48QCtKcWO/cFqPXk8+jOJzn7gnzKwDA5hXuV+q0x6BQn3x/xBwFQl+PJyk2iXZ7NqQONlgraJ8y
vWCzFrn1jzLavFsjXRRC40uyQajwtHYLwEChCeKdArEJmrB/wSf4Gn0gYSCTWTzNp9mLVzaZRi/X
LUjEMCZ93h8N0NJKEOa658nMPRJjf+z2JzCY8izgut0pEDwNwmJMbPEy5ffH8yOYOHgty/jKk1Ea
q7CUwjnDgTn2UVHrSHCKw3zfkYgPfcoQvcAodT15lZsFkEqb3Ix9Ym9TG+Qw1Ox84ZAWV+ARj7Q5
5g9Ve+7tcwNPEp2+gEHWOWrsjA6yHjTiWDolagobZiD/eQ02EvbRNN6lsdmMg0fE2Q3DqxIpyqs8
o7pFyUk5QdONXKUyDLUVI/zHfzv9i1u8/lM+6KGag7LpTsB4TXyv5gFQFBh1qZMGUe7h8cH9FHjf
Jm59keZaHS4Fit1P9UQsxcYDFgg8g2FFDwg3XQImk+tMYlNhft2A3Sjq56AlaSyqkzJDeHTXIjFV
Sn3zoqD4FkC3OqTVIB/e9YYyRLkQJS8M5Q0P4U6uROpq+/XWr/IUd0CxEWEr57knU7iSjrg29k6w
E8ZATGU5etnuNVD2OdRG21uUUdhFhnxKJSAxqaimg1fzxr8qY2bjtGgQcWRXnJ1/0YojFBswldDY
T4q9LMUxRdSnmyiCvES1/NCdI6i+6llb1drRkANhKsLS09iJIJpN4HP7XiO0qrXcZbukF3NXHdGG
B37p2hQ8Re473ccQY5aG2oVxJcKqYH/vK6dNPshSYxb36jqnoatozDaeb6sxxF9NxJaw4QbnQBfm
4HPbBoia4fBJJ4fbPgaHXCsawt7kBw/bAFiTRjRg5pPX9N2GBwtSVlzDQ1Iso/79YAuKQc7zNB/J
R2t0aSHP5FbmLvAXYoPqITbhr6q4YZ106c3vvbRf5zSlEg1PW5pTJruzlA+O4hLMxTj2Ab1DSQd0
JbzZ+r2Xf1kcaenYz6LBNDIQbIbI928g7OPsxmn2hN0nk+JlqaGxuvMrvIUPSrbWdWdAtyXdNGCH
MGIih7xZbUWEjW+1ag4vb5NiFatZx5ueqQbJokPh6eBkQJVAHrJ7ggtsADgL5Ba1+fuWE0pYTjyu
andGJf+Lnn+IdfLU82Il5ND3AwQebVuP1TlucZg1tY0S2iQVm1ZrKRxNEr7WoOeZ8UWvHlXmuX+q
3Z4LCg1TqZphTO1erkEMfB/4NOcQDmen8cLvV6mNE3PGblbcfA0MkHSFzP2PesoGZShxk1zt7yIa
E2dOQyLnNlyWBWQCpANAmaAR1y1VHlNOfoUAAXkV10uvo4z/fnNs3GdYFckj8Bxmuiszu+g8XKYc
l6rLfq1uXRluKli+gUwGt+pwtkAOidCRUSOSnhar1XK3ojqc3W+cE8vVFpDtxclsgPxeIRGfQmIJ
YVUhL/Cs0ZO/4dcf0bSRFnEz4Gphi3IPW7q9ADy2TSdBM71q4zYrQg7XAHmbLwyO6/pqwyJFNwoQ
+rSXWi0c1DifTLF+8NWfW7fUiruUy7TaGQm6hBrBx4MhbNSDJFcwJNzZ6k3G357WCIzQxpo1PlSC
nED36UmpboSQWPMYkzjSlgofYGyD5Gg6oHz+L5Qz5/b02aPeQy3V+wquERCzLYWExE/uG3quA/Yz
Re/4khbeWeffnAkf1fCaRIzLs0rUHZyvu4aAsE4DFbQjt7dyJqvMDhtRdjMYdSCkCdz+4wwrq6ec
IAmNuwXYo9cZTzgfXmq21D+sFT05gVdbRNvB/LO7jkCvgxqHokDdKMbKK0GsplX8d4tLaC9zpuJx
szMDmK5Nb94r6qacrdJsYTcB27EgOq+7SuKk6j5lj4416O9wvVvAF6LUetbbQta1lHVtBATrVqr2
aJyAQuP8NkRmCtldzFKGjuL6fAS1FcML6wjpWjhCAWtTtvSpDYaKOkH1FO/8mziIMuBqEphSmK9V
eCAlfktavgk9YmtkcyShWBMSXQRetVzs+i+a30TPs8YCyEGMUIpmfnGWjSC4jNfKEX09hW8P3JpP
g1ow54dYojlJ8dBJ3XaEPfb5fJyBKNqWK44uMlLQRKzb+iRkMlF/iDIfhavpsB78YfCJzKZxl+B7
ic/eYlCCNUM945vBcX9OYeA6CreisW7BJfNfVhq5hfn2t0uG39cIQI2k9lOfCMDQhFbXUDE25wPq
kZCnYIj23zsYkhutPp2Y1WoJWytbXK/Im79BNwcG2JHG5ILZrRFuMTHuCEj5WnQzjiJHzYjZGApB
+wul9K4Zo6dVmjMXKEPyZ6rnH6AQRsvDlDZ4x3QioRjJlztTY3LT13FV8U7YUnDidt7PhQgFHn6z
tOpbpkByCnFGYKM8sOU4W9yWp9OLr18oJegDluLyYJycQ9aIlSExdILGL6tFdOCyZFlVnH/iJGSp
VBIiwpaQjMd/UuHbPMYF9o4ALt613Owgm4izWEHTXfpu/4e1iZ5iNUodKb2L/aSn7xpXWCLhRtH1
S9y+QE4s3oVAUz5U60Amk6UMBjpozfl5gEZnilH2epLTKk4J0Y+til0mjDJQwQ6GFQ1JPK97EewK
ftf8Q0XOQT2DHc3abbPdZpCkDVSBS4MuLBSJxB026gGeSnQZbEeimx20Rsfd0WoqV3iLqJhN9ijX
Axc5fe3niPFomE6F4j0vsDHWm1x+u+ORSqjN4m7pKMXIUmhrRwG+u86FzLp1ZHNS4Hy30xVM+z+e
PPBttpt3Pn602mg8QlmrbJnDFCCQXGm0YHvqSBuVdnWrm8xpv2d/eheNcSltCRtRE8awAma/fzlq
41MFFcOgvmWRe5njDtUKRJvoVUbzpry5aU9ZHatY31Iz4AZxjwe5gdjjvcwZHoEL7Puv7TgUF5vQ
dO0JTV5iF15Qqq/SaSgjguz6XeCjEuRdr+qtoIdDmNrnHDzcIGX1CDXUcVcsBaZNTBnRoYWXDAZF
pdwxB5wEpoXb7yU29s3kHVCnTD7iAJTScKPdaZAKBRzTmewL/hD7v5RVSbv1LEWYytfDbHTYf+cJ
XkSKhGV2oNcnBfJiL9ubd9uSMuy9tncZhzRzBg1UEyasCEiFQUZZzeCAJke23q/2FVqQTO0UjEAh
cMqbq8u3PZcZXD0JkD21M848vFQ5teoHLG2tGu5ugeOAvYVREJ9Fj7iPFGOdyHfAFsBQM2VbVuzO
jBKwcjNMT/2hIzjV0Ngzu0wy5p/S4ZcgZb573Vx0/X/LT/n8F/8rM3ux04UJ1NIf4T94mL+QEuaK
+ePwYBV4lhlGIS8PUN/BWGeX4JtePfwOAKuXeLjHBvR19BTgqvlAuuHWiPSjmHZfwhjmfTK9naB0
SGnQtfAklvtHk74i0fAqedE6ttQmRtmEaNHvHA8z5JnZSNlRPWXyhZBfquYBviJ5142/smLB519l
VwSZ0smkltDDJ1HqmgjqB2HAhunY5ShWjuOgyLdrPZ41vjSZTxnElNf4vi1rfEYh6Vk9thF8ZK8X
iTgOy3dBZnX8Lwg5aG2jbP/WZs/lhRKmH1DAngiBWx6xMCVjx/nfrsHgXbst7effOZ6YS6CaGVMy
I5r9mlexH0Y1tr+qo6PjwUkoGt0q1XH84f/rj/GKkSYDhzFBsCExByTUnJTPZ18yriayis397LgC
wma/a4eRF9vCMDWX2qkVrGNry9rRi2QJwZa8m3jjnLd/Qe36A2FfFrLlJjSutG6QUE1O9SpjQ3VA
qZJKdgYbasVSAj6BPqCp9Q254XtTJz67qtxud20ltr42c0my+Te14OyzeA5EWK05X+6N074Kv2X0
ZITL8rFiYOVWwA7IFP8VukFs9gFgun25N1OCmMo7Q4++2tyQSyTnLWr1rI2pagoLp8e2vLnD7GKr
oI07JGafbgGXV6IQeh56zpeEGocsg3ZN4bJzuC9RjXVqRxoAuzhPQkwTptai2ppyDUEXU+5dPVp2
P7WdjZojGQu0qILZXKiq98+bygbRcYIbcHY0JpKY/DHteYr6tgk0UUKNQJRXeKFog0Zx8Zb/ESKy
A7tW5OB9BSh2UhlT6xlqiyZGWshZC/JjWnu59cl/7VL5PMZobdn1lawCvEKhijMEHT1jcGE62dUU
mjq7S/GviVUK7L5RxKING6L4jhQuISTpCKdicwFXs2SX4s0XHMLgLKIfE4kkm2NiIxc87O8+DdEN
WBx9w9DRUKkm9jwXZ6uhuA9khQRpMsHavie1/vkSt8hSON/Zt9Wc15wG9HVGRPWjstCLqV4Mhp5k
DHvzKsohEFh2M9y69YnPL1vQJX4RTBpkqjtU4/XRH+tB6FxADt2obbYsrYWxrLH04yaq+X+McMiF
bQopN8OwidW4GnV5Am2anglem4Mc3KV2a4RjlIRutVVvE8DrTkmtdIlwdK+EpdE2vtoWmWsF4iQm
ALfSfhDLG5BvPIlSAts5hJWi9SwznvX23sacBECc//J89+zK6oyWi8fYvmriY1mt+ybf31wocj1H
nDZhMBmSFBTmjwtnllcuWpBEG9IXC5G95D76p+gyoloyZ/u+3a4GhedzRNL0jkmXkaIkTxfT7lz0
T6vxfk0TQ+9hKvYJuCquSve+0Ajbe7lyqFcnhozkvxNm+5lbcC9dTdtSq/6jJO+LBJiUP1Ws6njj
S6Bmxpa2WuPgYU4aG7/YLYl5xtjxYERSU+k8MroQGT7UJW6Wmf0zvlw0PxHM5s1xgN1rB7L9S56e
F06dQxNof4OAUfZ8g/fUXNnEQK+7H3nEVuqH1PYnCtsLH+AwXPGEKl+Rqaq4nkqKvUgGyE006uLT
34g3MtWNuIkntX3RMsv9DKb7zzNj0zTG6IV3wJk9L/jzj6yYxDOLYtYL4FAegkvqiieLMZ9pdojk
eIujkOQMohZ0u4NvegGX1f/jkcjLQi2zBVjy5yGqTxKL+5vsWtWVOGo1OFSvLzq4zgNGtw+SX5Tc
B3hBivAC5NSRAL8nP60yjnYkQI11hmJ12cVrGhO2vOfWn3Jo0TEP8M783u+JCzrwW2mt7izcs81s
LUc+bgaEl1c15iSTuDOy0p3L+BYY6xv4Z3pkJNVsX0bWCyB0eyh/nXJqxBEstUXAjN/t/mlqZXy6
1nSoPCYEj+8KZh+2wzikKQPo2BAkeJuibsIK9Ww1QK9iHNdJJpPxZBBXuybBk+rW/XZIsOFl2vja
aARAbJ2s3/5WUrmYhy0+R5xY5qGwjvQpkeF9vVGtvKsDkv+avo6TZXHEWWZWVUeyAgSqk71XXPsJ
P8msOHX85GmGSQM+jZQOou6blSnHsrHGqDYpO6fW9s08BNX0PR88smdw3kDW5YGBeRMg2vGJ73mW
JBx2sMlXTBVpY2fNeTdFtAebw7+SKN6xZQmqMp+V9scjAPi5mrB1+Ac9hcIqu6HwRhbrMcldZCwr
HLkmGfH3OhJbrmJKa438ehSnS8B2S0kL5r9HGWYct4+TzUiVYEV4jCxM/W/uBCXdqwkbP6iDokRZ
FtEJJaxJ0K/ravwOSo+Z/LjNl27Kxcx/YfQpfqDoiV97g28gLTErjFfmWngDXul70YKZ9OKoY4X3
G3iprhQDq6I2DPRHszTFbbG+O6Ooa5pJe2VlcT9/RhV57WTjs7XhVJMJhUDHZxeskNeLUIhP4oYm
1XwIYvX3NsgPLgfjQBWUD9FPBYemPEaUAldfh+TRW90JPNk1UnBjzLJ2l+XFhTqRMvUan8kRqA5O
2Po3cH4XmTkNK11oTjcGPyE1stluLjlDmpZIUxi9cWz2OSlCx4QuVxayte6l85Qn+0s4CJ5E/GL0
vOw2KKCsb29k2ODGuA0hJ4Wmc8FQmEZi4bnNkjKEdKnpiC0AV6MEufFYWJjMr/QGPNnO2HCoL2F0
59srUf0XhrftbRhDA5WMlB83s9BQPLkl+TTYkW4YrnoN9ejz53R2JP8Dh/kozPdlxNu+Hq6KRqlW
pGt6Wn1OfzEmJzjY4DJJpuddsIMp3gy0n04rRJ31/gGtaCwBeJx4gy/zjgYIGYUxyU+/0Oyy1aRg
dXTYDaHsI5EeDcjGkNnDsrsCF98fE/i5Tsb0mllF2IIeHaj9WgYWIGQG9Q38y9jkoouA3SSxMZ2H
5MgxUl9OawrnHyPvW+ZlUYlLUnzSM0FyXQCrhufXC6WlP4nLFND8xPy3LSJ9Q81mOKMqHTML6dBx
tETPeT0Oze3Z+fHDdDTJxjQbGx2MKlhiD+bIxPu4Ni06PgPQeJVqMY4dmTrSgPYGu3Qm93cCOFXw
iG7uYCawLmI8s4zazhzxqdJTZmPU4tBEMg8k9JrUar/1dwe1Ob9CKkBb1xyuIAOn3FZjIOykjXqx
bY4ooQ/2Oc0r8MhgcWvYYbI9QV2gesn5BSr6KapJ5tD11HaDwul9X2YBZP46rsQKNYq6RmMAZdaY
0Q2umP+KJuXZJzewkY1R9aMg/40jk2mhqpUhr2oX9/Zgxe8GJigffs33pTlDwLO2Vsw/or7zj13R
KbQrhFXVK+PVhB5a6ILQqqym4CE7AT2ceV8IUeqeVrhwouiJX87u45ZWStTW2qr8EKUk6i1yXTze
qpjHnQWE0Q0+vAVies53z1PKuZqqQZ24UnrQ0B2ztZjPIN0QaLIADEfKzH0g4jQO4abwuxyj/Zav
zt6CaSXFVt0Uked8K4+NmjWuOwXLcNVK2l7JnkmNJ/Xdb2De+v7cR4weJb/rQnJC0Wh7qA2aq65P
CShfZgAdYTIkh9hy3fptyLNHWlRqakEOtEFV1noNnaFriS2G+aOikWMBQwnGR0Y7VTKKaXsqABXD
gS9D74KrWetAHgYJHdrqvbZlYrXweMgvvSGcaC1xv+qu27Y10fc3ngBMIKgpZierUh2e/Tlgi2Zp
9eO62iIG/g6Aem0UWYKZ4yu2bZBm3WJP8vcADlL0/7JU1cYdapv0y0OYxsWByAWm9y2ml+15eM8M
U7tmWCgLrUH8Adw5JVhlZ2RHhkYbYYLhUOjyxdXOS9tiqqBYZbRH+vlF/caNg5Qok2/IZDa8S53W
dhbCbpmozyWzQoevrQOkDQ9QJ5yMFuRqJsJRVmYC40R+hNjsW4qbvfb1irSCIrbzWL5EEbp9EYcI
BgRPCShD8geB+bL7rD9zn5vZv/Bgw3h1+NWDENGtfSKNdcGymYrCpo7sq8HL5EQRpsSmjNN4kaFv
LFAK2OJyJA6eDY43sYpi/YvPTcFWxC3KK1bLJ2NCEP6BCmm2UKcih8rH5ZxoK20Fkb7DjZ5o7d9R
SYuYjJt7S+YWZNbo0HCPWM9sdgt5QjPkn+YXocyqKLZ0iooGPuoYzxjIzmT632+qjjQYrgEWiXog
MunPovnGLG4DgyGOPdIwqNcUF0cnukkGIQBXts7i2h3wfQAbCFTaq/iOoMHtYya52IeA+AQCYP9C
P6c4QCgcNHxo1uKsmGKo8apYkCB2N4e6Sk1Y1j8ZavRenCtPkGWvvUFQjR5R1WsmMcvnHJRmWBqz
PQ8XZo/NlOC0R0K3CvVOSua+lx03aktO4vDS5wGoICvka1Fupxoo7VaN5tQM3Lu2MapnbP3Jltrg
XKp7DX5hUeqyG/yA7E2NFe8h8zzb1eoRsaWm9yPOfUJcLn8U2jVBGgcSgPvYzEIQ7UJ+DbEWSn5E
Qry2UBYtLEi2fIFFcs/V00yEZwfnPbCUwfuG+JOQyeg3X1mhS3vv3QcJ8yptiUxU7+06t4Sl0Et5
lh3u22XkcUP59xcv8AL7ulMUEVjQr2/WVOnyNU0QTmawAfZA4reZf12r9Gy2rAE2o0QdY6IbQthp
RbrCBXYlw4mpk5eC3JfO3DMsL6wfmt195KFsxjEZ9NB/+U7jIfmgcTl7FsnJtHHjst2oChuzmqb9
ScUFaV35dX3czIUN0WiouYk3ynV+WgIj9p6qsrUQq9aA3/FB24ovGvAw+9XEujdVbpS5bAZRHhJS
c36veUfRGC+DwzTEP7dgVoXwuXbQPpBVjg5GtqM+uVUaafygBJAStn5ukYKh84//rvob0st79iJx
U1E9EfNhTfE2dk4e+1NVbeK2ULB03vwEYhQDtmdfp/d5D6SqpgLhnvqTiD4Ml6Frt9Rq8ibj/T0g
+Uxrn4Hb8EvkqjP8d6iRJv3AP9rFWcFgvPyuSPOc73cmfVjRSCPjcUJFKEtLpt4eHP4nG5P2igK9
m7lZyElxve1/8Mfos9epN27NMKCoYX1fTvWKGV20TfCTrOOS8MqsgxESvNONUjQbMvt2j4nYjvZF
FwganQ4nsMt04/lHK09R1J8fH61HgTaqXIfnZNLOjjYlIzetOPmqTHcBGZxg7W3jH38gynaX5bmE
IV9oM5LLAOX4I3sydpDLXEFMJbT+e/QPqqbHUHGueD0WJj38bkf2YjWD4qbrMv4RWeEl6PGD4DGc
+thUTuqFQs1KuvjoreKgatDxg5VvNw3AJGmkh82vdulYN9LApFtSGeFEWTX5NcJLbqpnJnnA8VG6
Q/Kj0P+YhBBn1cn3Iv/im1REccDvLqESNgLRMKlylnBt4yIUq7LVXyBdTv7AZk66yqpuwDayfkGL
lAl4wOKRYyOt/mpobXdNbuhBoRJLxMlwXZmYmqkglNotOTJ/p5Aq+w8L+vTUwBNR+cq5NgD+Dm1Y
Sa6SVuZrtbxhbR8KpJjs+FUGiu+6FIpkkfdMkouSZid1ThhNBoV4aa38N/j08Rks99zrzXow//Ku
ZyMnPimWJPqYq35jgCNSNE2XXB0LWSvZxNZQISs0VyxtoCq1HnmSyMrzcsU/fY8+51vlDAzbq9qT
QUW361JzBi6/zFRK2H0x6vYWPaFt+lTRvtjrWkB/9NmriaAvMOc1FaMiaHIsb4GJf4QY1rGM6y2I
0SpHfyCm17XWCyjYvv/+e9SEm49n48xd1zsIGSR0YCDq7EhwL7zzbSD2s6Mja/KKvv3sowfD+YFU
n3346prT1pihJVt1cMRHWmGVFnRsDQbClvjZenTmmIGIpTGUvnCG1c7lp3nTiIJCBjyfl9naFOyD
Yu2NJiX+6mbcM6/y8u7BGKtZ61bp1OjOXPUf3ICY1zdrPLPLSgdr59UxmSd0NZBfWh7VLUUzoEF2
sX06JjfukjXXnUmyE7V1Gbl+7TEnP6Qs/dMyzvYeoehRdiIfSQtzIqfMut2AvoBvHNhXhhhthXxI
c3LGy1G7i+IHjm/pCBiyn/9vVJ1WdGm14sj8hFrxuREA9VylooGN8wpGgjDkEknD9k9VS6tK/bOO
DvGCRLUE6aeQeHZvSC896BV/Nw/nn93XigQui+NMuBvlFAJ9fNTMq2R2S9cqt+TcAK9S1jefq48C
CHqLqhOY4wpkY3ZKlqYDSNqsNIGdX67UMYQarXVd7ATEtR4NsysvxWa8OD3rwkgFVTW2weHXLS8l
jh6yvNMgrgYMOvpsh0zxp0ZrbfaEgZ8UKOt4x/cDg+I1s+XA0OEshSp0o7Pemy9hi37IJ6TAAofz
j/kgq0JeXauEp0Yv4OrhONjiK74HTf5FKfQYiS98WJD//5VTcLVU0EdkoQd2N2Uv5aFbqZdJoeT1
c+xKh8ntwe2lyCwkbYtZHO1xnABQP3Mz4jmxrF7jyq1/QxK4ypwErID7hSLxj51HsrFeP9UUa0LI
T4gIr2MpfzRWhxGcl2o3KwmGdW+3F10m0bZ+rn6bUUYW4E8j/hDNx9MFSrUGDj+2HQeOpRMuZt8m
lmk/KfbPCk9onnqCzLHr2VNKyG9/4S+c9oX7mGxGOk7EZdbDa4td7XfH8LQbr7UPuldsXr8KV8Ds
er3DjlK4TkX0D5EZv9O8oBnJR/W3Ry99giqcfgatyhItvTav4nSTscRdwOFi8A+6Dcv++hhgdIhG
pbcRlBO5Y4lRo0vme7BbV+85A5XiVap1ykoEmTw6dAVLt14Iy2iWtOWAYsTpDK4puksAmdFc4VqM
G3cn3jt54cDmWE6FU1dD576IpD7UhbCA4S4NdXMdW6+vv9o87ELdk/kpei3yzaNd0ErXc4TOc3F+
hb0p/ZexkVrDF5cZK7AMdbweEvVKXMQ3R+DcjvGNgiOhfa2FOU9T6ZuLkwPPzo7XaP1Fpdh6eLzz
E+96+mhpsuIoOn5fWhR3ggfcRHE+akIgRSa9pZYjjKrnFxLLl4KPzue+WHaBV6QuRt5VVmfBuS3y
DRRTOKQC10JyWLUO8uDNmfHYDoD/ud12VL8roQnbRzTEch2RX0aaZli7iC8vsbdQIm3U1TlsOFKH
O4CuG1VWEkRa74Wa0vETFJv5RIm72WKaAasC/zOkl+sBKq3j9U3adsat84Aev4xKeMwztHNm9l2p
lcv22aTk6Zh086y2BXASqBxmhCIVBXapaWFOVCRy6kGmD2MwOMPpR7vmWXnGUVbJh00C/T9ZNIkl
34l7l3v0zTz2p7ZA00zA5vKUzdGxGZsQf2kv/P//biODnU8KH4auVI8H4GfGERT1ryC6mKX98AKS
0eCn6FtfmDJR0VHWmYukterZg/KrR637E8x2gNFWiDOhKanKnQbC22/f8G84kv0eRMuskd1mDWD2
qXn0D1Oet6FssvaM7bMbQTVRnGgQVUj5ZhROA0WmSg+jmQIAeKb/PLfeTmeRZwGdlVYhs/pVmSCI
BG+aaDF8G/1l9vwCi60vxdQj7yY9yNzFdFRrnvgiEFYzNeFIY6nWquDF6mOtORdhK9U0Z4G96qko
SXYbtEdjlQ5QdRK72A++fpa3kqZLEd+D0kJUiDGUymr/7AcNuBIiESwCTkWiUcwycI10UY5n0tLS
JfiQXlIwF8pGMD0hnvOchVGp5v4+4ISruiVnb6KLWEeMzOPppiVJ8qTGJL2R6YlA5gZ2hRLypgcW
kRCb+KV9vRimR7W/isOkybX6TuYGq63bMDisAm1KunVaiLhh/pCtBe9tWEPUlLLw+TWLhL5tkoJ9
9qleR1+Zh6V/3v38XddjToTfngU9leDSajsdtUOelf8doU8KtUiryZq2ANOkbutZ2YvuzonAVath
mH03eaWP+AB872n8q/7WRRr2lghCvfeAZ2ITkh6gzmPVdO0+ZAVuhFfPrNKfWqJPyzlsx89EL/bC
HiGJimFflH6j3kd7NSQkPd4E0HnAoJWs3txW/CO5fTh49iO2PXiiHwJtHquXaZn/UiRCQk2kqs60
zpZUwl8B4eyETkGVyG9Ui/0SPNCuuNQHHZ5wdvO1vstdxo5ksfMxeC1uNG6bAs4WJX5ZPD0zYLkU
kQ3fmpEEcJOhx+AFmZv8LrROduAhw4PlmWR07yvpWsfmF/Uuvl5//CBkoqePnr1Gc2+5Kl4R+LLT
9TfrqcCAAGR74DpNcqclvfPDRJ4HXezv8y7WeUL9EAWHmdxB3rT9K5BuwkIDSeJXOmbW6KIXSsEc
E6hV/cmZtuRftpfcryT1/2zqiCiHLPQux212Qtz/E3VHgalO/RNth207lM1nXpr3eeks0vgnoSmw
5aammgmEOmK17uYvc/OO7+CLChIpmc72MO9D4V8CDeXMDdP2Wgh3LHSOmWZ0//FY6CKJf2RvCTtz
OpFL3g3kJxj1+F+fDbMt7nAtnGhFYTb5fSTiV1ilYCFccAMDyVxPVv7ZVi41qixoXw99ocfAgjXL
ZuOc9mk5zso+iS4gHlqfRYK+YGuxneJAwTxWiJVda9abgRrTR1VRw1QIlNZqhcOP90HmZlSnJTdP
w7HkmPKefLo07TsVGvuv72C2kfDouWVtw7SyqlVbQr3PldhJLEBPRxAg+IrUd0lMPvFMdcWJ8j+V
4tRrW/xHy6P2wR5e5AHcM3CuaQsKl3VJqQexl9jQnYdYhrEJHp/HmzTop54Dabp+zJvilGOaW6Kk
MnnfUvcRQ9ttI9+sAeJs/nJ79bLuowOGTS7M/hO5b2Zy8P6T/jcmDqBUmtx/OMFTSrZMDhtKD+L8
EXIIkmuG4gzva0MhL8WwAlvR8NRQ18SsICZQ1e68RWBNFaWhxTgDx/PV74WdfAWHB4/Ega9VmsOq
WCbSIZBswgpwxIyHR7zK/ucRkTwFxLEsQ8Aa6RZRYo7pqUqFbIHm8uLat4bX8W1zH4CZjcv8z/2d
UvuHiIwlkqKcchvulRUz8yD134CWItRfDgo5CgkJLgdDQ/YAQi+WHKO12hCJrMFmyuWYl5JYKQg8
oq/I0meZ1ssNG1yjBFNHq7NuRkJeH37BylSwV6ABfiekREsXvEwsnEbRzZRO73NWXuc8dUHzoizt
MHyUYFdOj6K5I2vNKN9sNTL2THCYUZx4nlr+sB96XD5PiJk4M6vdANp60CAy2J4ktx20ugjBx+qV
MqYu/NxfeQzpStPfYjqjO2b1O6QNeknriCeHoOOO/FD+sJDLw+F4UdnvO+q/h+Be2u80NcTTL0JD
T6E3LtvWwT76Qs7My8WxKTQa29AnAWF3dwsV+GeZnWzkAlDfLaK97yOOhPLjX71d+0NrcOug4Ivw
Q773hKrsPe+npS7FAl4MS/kMMFB6EcOXdoyPGk727G1GdpMupLmWQZWYDSxodTed0tEPlq7Ws74s
lidUN+Tpxn0fMJRnf+YBqqciPwdHNXXZpdUbkN9xlNAbZiHKwAzqQGMUDmriF92dGVLSFVnS8r8+
NtQ+B0dshJfjKVRPbuCcjNGEy3XX4WNBZ4GOlhAHW2GIpev7ZrhkKr4NayftDZN1dYltOfqLlfuo
ZbPPI3HhXaswZWb85Pc3GvwtJnkQcMwanx5r6uUl12OUVWgv1hU/ghXLXMHyJzgieZXRBhimxDtr
JvzYO5OmdVS+obtmpQdKo/4xiXQdNyyi234gPPztovsWFcb1AU5gba6gxiHFRMcdS47K4/3XAHoC
IBPio4N6r1tlwTFjxRhpDZ2YEnEJd/jBAbasLPq1mlbBh5ItL4sjRF2iisn0OQFWoU0RFyFE37io
ijQ7uonJKh5kRLv5axTpsiR/Ebn2tXHappiEhdHL5FqxbtW1DsR8IjbxY3AydRQKCVOOlJNX1Jm9
+ZXFOt3R0CYBzVfcxSHivNPQZ4GKPGRmnW7m+/20l2m6KvHR7XSPvJbBPdxOjYsvzrhPbrOl9Tz3
ZovKXVFORQIMdRB7pb0PCoRNiazWDKxS/rhPY9g/d2pXa82zQc7JHJxRCK++IIDmnI0ejVjWMWnj
TXxvPa13Dw9+yJzEl/XIMrPYlzch4O6Kxz78+US/kucuzwWRKcWPSS5jSfWYlD+QbOCS8wKWg7Jd
o57ICFAyEKIz1U5pvj8i6VLE3ewxErW3DGHmNnxO1msaUBI8W1pFtsUZEr4ClPugtImvXHlMXJqC
9JHhUUqHZLKGS+w/ckUeVj39HZsBk+1fOhBkoOa87jSufzAQLV6ph26wrHK/ZEFRVKjvRJ/P3/NJ
ajB8GnV1DPFRhN2gGBGT2Na+2EZ8dOmxGLn54Kl/vmSGDosIE0MZmMF1KxBqqkKEqiFoIStbUf/6
5Q1UxcaGsMoaIATRfL8XBpM9tT98TWeysYmZCc8TJT+29aXSe+KBlDZxCMsDoVXCV6XyYAjB3X4A
HFg6KoqUU4rGvOzUMjNCwzJ2tPEokSMI2HGQaKxDIUiUJMbmAsLSHJevNcERqFq5trMp0/6RG56T
cidE0J2oCFZaR/dg6mbQiCApBYTIgrHwqL3pHPkTy389w19xtJfxviTZDxHhEhpiKR9/ts9cSCcw
PoG6gL5q1/tw3U4Ijm6Swscce/Pzj7miYE7Pa7/7AbgZJiGnqjXJciAehjJwYpjHeaEQ9ULj32CL
d0MfkcogILq67K25VSzZw7EtGDmYjCml1i2cCUtHU3bh007nrfQbhuGeFOl7i2yDYCsm7TjVR14N
vkudsixzA2OeoQAGrchSjnkDNX2C+XPY8Kc6DEIuACw1ccnq148MCXrZq6g0Om4FRqA/uXJJSBR7
rBTsQkykkITlKhu+H8avTQzu2PT/0U2av6VoSQdQvugNYht6twhFltXGSV5gNDnr2rHMaxw+ka4D
q1Oh3lDHJ+w/QEZCdOeFWMz1SZGbJF+l6XMjunyfZeRzdUKCi9sALNhhDxwiRu4kPMtIb4n8b/to
TEGZQEYmDI5WXVTxqjUw9cDFHihSxo/XWarrSekVP10d6kbG36hvW9LUlH5+GHmJWZ8Caen1nuaB
cseJPrAPm1vsAmgZi3GWOmOh+tCMxBrisX5ccZVl2jiQ7ADzIhRKfnVtRVTDEjUXbIoKkZE/9i10
CxECo4X17jd/PWyYyuRtURjXjJf3NKh4NWT3TVYtpNmngKiOI1TNuC0TsRwoQ23xqQMOKaCIZWRt
hIeL6W8H1tUiWDPb1rmCjZzA5IFmXvrbyD9Y0/C8Zvu1uZP9sXw/OA+YIU4xKNLeVNhwrMKOaBWk
bFvnURRZIx0XWQKB1c8AgHcqQqTz+lr72H09B9q/r7WbI9RUFnrAUueV2WFebDfMGV5yxU5Z8M4/
x6phhqO/RFKVaZ5a8SOs54BXq8oggW+K9nbm3leoBp+7oAW0rNh5aXVfnJ5sCF6DymOvQb6Fomxp
U9TgK2Q0JeMJlUza4SMEGsVDMjiQA+E8VorBj+vJnavlxTa2ow9zpTyPKFJILNDreC0Q1owzufjm
pf8Ldnshy63yOQ+ye841cof+9eH5lkS+jYsAbNU3f68zhfn10+AUZOzKcYnrPtZJUpug4qVzH0z9
fR/a+U6LlhUlXMbDz835UnCSSauqy8ZP8lGJfPr36CIaCl6/bjMkWiekzIDMS6E7mVM8jw9C8Sl+
EmHyuH1H9JfnQJWAbwxpfJ7/HRx0mRpHqr+8F8a+Ix8bjAflboVtgwTiO/26tmw32b3FC8OMVNr2
JfBfAt1T9SpgqaL2EXErV5ZweZPNafPf0uE334r67/ZaFiu3poVHpssZBzp6ZzET/spMNTYocuXM
9Zr+EirIaswcYTi3Q4ML3+KvFAUUzEN/LwATyXAAizzI5LjQv2xAkqndzyT0CkhmEdfOQBsgy+pU
gIaYmw2KCGs++eBoLkMaeS7it7ZCY04o64EVRfa63o3hQwWYd7tY5v7pJIxk4nV/N0dfBQODPfr3
RDLDmLHKIErGZugzAuspG5vQnXNDrv6A3QcttCvEZ4p7oqvScux+jRctE+QoxpR9fyb6vQGEJ/1m
M4yDIn88H2XI6+Os2X+ulJRJt2WQkKGIlIItWyuZOjnHasEHk6pV1UnyDig7QN13JApWrjWdpFPv
g2+JCgYn/EVVVLuerjYqNSNatTVA5YjBlBq410EBQzJFYCc4kPvoJQrGj9pmwCSkyDGcNzTV0hD5
gv69hs4No28iG0pdodLEPRr3Fh3oLsFw8my/26ExF2jr38lH5/Jy0QljSfk2VnYLjTmVlHLMjNxK
s/lYFuOIpNgkVM8/Zx6zT7bSyo0zgAid0alhuNnwO/votKoiknKs2EW1SSbK8uhDppzYO2j+Ui/b
mcxZANCzkh1UVpGkvouwv9pLGkH0K4V0T1F7J7KNMhbOQEo3l0Y6uYSzNzeUydTOnfIU7QnDBT8A
IzCvpuOBQYR5X6maEhfdk3MM181odB8+jLlcBGgG/Wk5wustcw44ZHp6YPsvXxb1luTVfqZAvpY+
LgSpThKujG5y2ylNmyuRIM8DA12TgYn6Qbhdz1fPmLxJuL8gJjLeVUStU6UBjk1RwHCpUYa8vuaO
DYdUhSFSSIBqy5u6cOqskqFJzKTnF4DZyhBAiq689Ei0QaaZFr1QqU5wHfKTCH9ZjmJ9wRvaQdyP
GUG8Ms76kTIkOcqJbSVSgspuAdyl8yh8/g4YI1qtylGNze9zkBb3xE+QXpwwzH6fOObyHnbhD1AR
BZ0uDhoIZ9GseMJDjxlW+Nrlyd9nXl6eeZj9SVAPlkQ1h68hxBqC8Gw4blUEj/7u8x3ZTw/k9fD8
cRu21VwK/miEekADRy3vOGYnzViYbH0Fh6wVqoK5Y58ilIkVo2onw3VYSZzDWlqVof5XpZqYJj7r
n9mjs104rwlNHIOY3rNSE11RvSKKLHb2k/h7XjaRSDsOIcqa+lZ3EiMhqNMzzOYQO50DOa57kHRL
glayAz/SmDmQ7duhwzLqPhNqUepQ1OdkXOk3RqSiT+MdllqAMBI2JjE5JF8I7Xwre1GubiNL4sy/
KTphuIAglbVtSfSj0T2EPavPy3GLL35cQP2023rQvTsl78onOoZWzom6TLcBUTQ/7OoAW3oLTXdV
QI69M5D8OEt9SL4rsRjvcUtNOim/FE/o21zFt8AaC/FIwV0nsHEuU+wUTXFo7qNEA3m5ayAFyj7u
XRFTF+YJPT0bQeTDk/zPQotcvPWd7s62/eVbO7ek24tjkgbWYeEsSdKggPUaI60w609crTzqmed6
iFKNhyGrRMBpgBywjZbH4FsiaRwj95to3+aVkbN+p2+Ef+JOzWMWuZ3Y2Ym3n6qcuSk50F3LK30e
+k0tdq7PtS5uIW8hO44Zv92+G83ESGWkGj5xwkDUSXBBkWArEadj5g10wQUjM9oX+eXGOBkgJQLF
HfMCjdO3+QuoEs+N1ZVGakYN1e32rn/EIvuUD7KYLo3T3uakCVrWKq/fhwCb2MWVvAqKonXBbvrI
KLkNC4gNFAXwQ/ygXP/MKV2ThuFyHvGfeiNGDQ3GihgZbeGANdFE9Wnhm7ccGNE/eckX4kEtnckZ
vXw4mp2vyGXmEZwhnJO7jUwvqiqNgfaZ7EYaFXRbwPzMhdtm0UFYr2YDGX3jIFSnqokXzf0tzirX
vJQqopsI0k58EpGxtepzIhJQA182x7MU4daSnNGxqfGAR27S6i6yIkyDrh+LPZrMrt+0bTcBTSQv
b3pQewbLvkFOlMG4hrAuYisMYkcZDBxpgh1VwsYq+5sPiYRt/OdGYkNY7f6BGjJgmthmrTVf8dHZ
ZwhxV16Q4W0BVzn4vdJgZgmsWikEA1MlWIZ7wkQESDt5coTeckvwFKZKI9g9TS6Ug+CYlyuvVq1u
cuRrTk8JrNLYvFhWGnwKSCH+o6vnJAi4P4K0FaCMi+wz+LeiScZ6+ZA10m+q0gaW5U9VIDZ86OGu
VGqKG6m1LcspKNIv4neBmVnrGaOOUvFgvA98YMNA2qvgBfz+2qpcBrEIVnmOHjzEtTtHoXWHrB3T
zskA/hRdRD2gRaK9QfWo4Sodb8P1fEP3MkoXYY4td28mJjsdn/NX+ZuQK5sRoigPM2Am/MrmCRQ7
TimORjGViZ3+8vHJ2hZnYbgUXDX/TI9w+/DhDXB6OuOT+i6Uj8mAfr/i7lBC/VdffUq+zjkaUJCW
hCUjZzAqVxSM3ZpoGJz5YqZaYHfPLxa1HSFRZ518+e44azm7DRhpN9i6YmMLe/OpQb777duUe5uu
GY/Cdyau/XXbzk3wvJNVa+GsAB3njl3cMlghMoiy7h1t0T6qmLP7W+khK55ItesAC4UUQ8RAdFWw
oo0kasEjTg56MH4HbQQy4KwGbwDqropxFG7V4MGNNC68ygXnz0qeHwRXBUbY4RSrm4bv2LI0CkIZ
BRM8mxUh2AT8N/Ueqgydumg+6/m0xbOcW3pxUmUQzpHXJbTGLlB5cXpKIa0vEgZc8ADp6NsQUT/P
ThBhvNvWP6jY+CgRb0EaBTVBf1SJGNppcDkwAv0QiRTdLyYTX4NdUg1sGlB/JM4TQI/YX4bb89/m
ShtOjmKxJnJqPeWzdesCLH7IEVjxAegFZi5nRoW8N+uZHj5TEo7DnAhC6QJ74zzQCL6Yn5NDJ+rz
Dhc7mekqMGHP1L+Pfu02YKJkbXsrOrMwWQFi2ItJpqgIcfj+sKSWHYBG0Rh2xiFNpv17hnO4Agxt
MvMTMBM1Q1N+RGwQtTu8n7pgGQkqasAUsTpgMNrzglq+aTX0i5sHVW36HMnH/KfsiVJayPfky7nY
SMD96Wzo44lHOszLPU0jkNgeTerbQdSqG5Tm9V1Pv4aSreIrbzutJPRvtPKgio24GaDe29fAkxUo
2U6HreAqVlgsvaCZ3xwhOSZso0mKvjPfvhZaRd5HIr4f0fu14rmnrxm0bTEa17QrPj09S5YXWyPF
bPwEBnCdNNQVMT11UWClkrmqD8xC10HZiIc189M9uyUG0dndo51xT3YkImpXkoXC0m+ihmA0ns3V
NFPenADDQ/fFizChzbeP7uGdHeS5T0PcFyL2y3yKhRnsqym4H6IxR0rQlFX1TQWXz8eqcx35rtzh
8DnjTTMxH9Bck+ayoZg0VOW3ELwofbv8urJH4vqQ7M3vtRfWJCiheTd1J41AVCs4bsYR7oW5Wv9u
G0dIi0E4B5xITzv6c5TL3iLkN5B44Uh1raEfGbdbGaew0Tu+N2Gl1ZcA0TzH4115tgIeSheD4r+g
i2Q6OAefH+RGRTduutdtD6JH74qAsmcjk2Q2IKw9An9U+AWqIoUY4DuqXi8MBXvIMKe9To0i6jQA
nXe6BS3ITm24+TL7wqNwRqy5biPQSs1H+hZwqTsuyhmIxpKYH/hn0O6mMlci2cTeTquhdIRbdfxW
/eC0Hk+7gawgf1LHgTGGvBurd1CzFIBJ1QwgTt/XDDm9ox9dLwspzFcyR0Z3w1xv4bdKqyK/eHaX
FeUOcjKiBMRIounPI3IPTsQzEIoVAHc40oNFddpX4zs7aBFZCmk94nTpLVRth8bo/R4rwQoi2toH
LtknNX/RwGKzIDQVQaiMa2ZBGJp3fJWN55uaCvMrrQ79B6P/wuSRU767OtVyVcewPYiZKGZfaPp6
TZdEraJq2ivNqT5IND6bheAxJNtocw7uC8xXLSj24o44l9t8RnAnJmh6hrjjJgAzM904TLYBnZ7n
s+7UrGHU+dEnd1FrTBnFBRp9HTzCTI0MeMNLgiLfpemuuycPVFveEFjDju2z2M1XwJ0mIJ4iYbWX
9m1dtbRVe88ToVNgQEngheIIR8i+LGsJ9h1i1R2h6JI1DcvsxWLzMYNhMU+2zDyq8BqdiGn6qBQI
Q1bSt00Jv74V59xLDoCvQCge6mgOV3gNCZVNEqyiPUCO2ERnQjoBTR3XITtInCmxB6UE0YysctG3
O2BCw6XZ0ZB5cE7wWp47qmk5nA6MtnllLGwv8gsO0LFHEJV/nM0qvfG/T/yVK/D6bVGXbUbk5Bsy
No19UkQ9CksU/Jcjon8/6xfIIWDo8VJ2P0XRWJ5sEhhwR42D4KnOMA9SKm4DEJFGBaLl6gZpjd8Y
CHL8mboBVHr0xHoPWOHhtx1HiNzZZ04/DXgerqwXceAJw8l9vTwPl9XGwP23Qmif68ueSeR8UezL
xM2VX/AF6cuavykpkFx8BESRsWgr31R9GqSnskvGp9yGNx7cKK3ZE1tiWjcbmuYnw4bX3N4gVUuC
+9ATL0Z9zgGz2rfQs3VFEQWOlqdlM4tjjceGOs+hBayzE7cKwcWjsQe0lsaRI417Pdjcoh861LT/
6JwCzC6wBZsT5rKQzBfk5npmK2TV0fHXV+LxXyhlnhuF1Y09d634GZMBE133W9z8MPa7+u1/LQvQ
uKYyDOeeaXE09tJnestpDf+DBL9bg2uremLx9pxT2oqMDWViXjL1dXLosc2SZ6ZMAS0nBLnOzDhL
qfB/EdMD5J7kx/KyuZjVx5OcBeiQJVy6kK0JFBwZLlKd0FAexsA100CW5ACUpilMm+QjF5Ob3Knq
KnXyYTgzJ75/FpNIMeeWDUu9X7ne1PcWk0esHHaRl1LzqsWfPnDCtlkGZaq9jsKdcnZhYfw+KNC/
JVuEMe5J/XRERpNdPA0BJsC7pF8s6/9x6pX3ecm8BJRxfibTFz/NsV7Kw4/TWT+DIcWbBqSkI65y
j535xkVjltqzoa9mZ1L3N+oOxMNUYnO1Md2YvR1I6L+fcF3U/c7SSngd1Pa8gsawyx6Fm67Eb6h7
6EmZy982r0eHbEyFVoqH8lcq4mK1Q0zLavudXjLVkD3LEaVZ0UfDxpn5tLUM3572fJSIBc2LMDFn
f21swOY03vKn/BNzeV3D6jKFaVHqWTUUB1UqMwMxQK4TRGaFWvqOk1M45etqsZoLY7RBEvEMri+V
oNmszm8Um2NkPkQCzKGrqSs2DQmNwsL4OfbG3M8//NQLjSHi4pwEEngqWFpQuvGE9vaBrnsYQz24
6X9m2si8iNxF29+VqCRFG1P1jglLP86pM14Zvm9A6QhKrz6WUgZ14WIYvQITNCT6NaGm3AOELDgG
NwU75P23IRiu/0KtpkHHt4Bhsi8iHrzGcJzre/+ov7KURf7BAotP+Y6tYUXVOPAPEp3VuJS+B0c9
unsG0LcxlQJkqo7St/Rd6kg8itc48pXHWhHJC8w8dlcmvb/hTC9abSqAT6qyRtQyLUl4EJqX1qQf
pfOH1QRgpHnhgmq6/QILOEhoQInxY/xiSuEMTbUiYJLy3o9kPK1cI4sH7xnTxx45TdG/8KDlF3wc
T2siCQm1v+8n2cPV/RIBpUOPy8UnnOE3A+CO8/+okhlDsCJBiiw0cUm97+bj1RlbgFBA7KVypBgs
0MRyGyz5HAWuSY4PByuY2zPWxz8O3mnCAltw50uTgRHWQdWGgLG9aqg2nuNtxpwF19CplcnGOOUA
CZi77kuCKzUT8dIePH6INXVJcLxOj0/9Lxek9YfhzxnsMgWUXxNTIKwq1cQ6JvI2xygOW4I8vg3M
2WaI0x0Q2bXKBB3pQyphp3WlnsDotD960kW7kkgh7rVVOZuA8JbUFvz+FVNkZkVjUeuYyp+n0Ueo
p+DuiVC1YpafR94SgxH+sVsgfuUYVI58ndadU0n12Lz2jDf5hoJ+T+JrA1MwRAmn49AtqLgFgTwC
iScsrSet1VtMcsdUVSvZbe7v92yqv1I0gWTyl3V/jswT6pb1/mkPQywUyY3cmWdSdl5h3zTIphx5
toBhY+AmQPXzQW231GTqFVO2BmBPzs1qufilZapE4mJWEcZ2KOr2Py/duEy8mvg8Q8OzVUYYpJnB
RlniN0tNyF3HD2XDO31xBe9Why6u2x21MC1YAJt/ZeQNVQgJPUNl9qPOROuvvZTKZ62Q/rvFWz7a
DpJ6fvB13O0Be43yJhoIWTzlGgjlXfsLdN1VftcodTN3Fii6MvFd4RbbU5WYov3ecqx8VRMVMhds
F3UpxWkv4uHXouMvPJYotNDbP8dc7z47YwFwptHRxoF2rkXqPkyt8utf8cK7suqtK75k0jTHZtDX
s9i60fu7PtvBFkJmZvQSAh8CkOSJotnLHiq+Z4frMz0vMFqxD4ZLH+4PUeWD6m8iO2UEiAEf6jhu
Z5+w+E++kIq2AkNdvtDD2c+DCF5Uj0tNZTh7IPYH3UKYiImnNzYhr9GtZ0kaHl3czPls5Pm/Po9d
XCJ1Q5o8Fnvxk5j9WtbHZqwkMHvwceAsZ2Ta2EGv2rZ1XShlOS1jos6Ali3ae5XTK1M1dlSlYYBe
a2jD/hOL0zcicgBE9At65iHn/H7uA2m0K+RQDzi70Qbdbk6CFwbkCu9C21yoymJp4Nq0BU7N5JpT
lWQ6Lt4F3r7UB6X9m7kAxEJhuXcRyqZw3I+bH6R/b30gPsLy5N6AI0aoW8VgCNe2L3u7w0rs4YYh
FvSNEk2ij5cjn+fQFQD1Khfoh88h3yI51tgEfgJCJ2DhVEhD6ZGU4Z69O5lCDxUat9g5AdN2mkm+
3MlsfC177rk5PTmfWiegeo5w/xNYvbJIjSlFtdpl5NebIqwk8OTgCjjcgciXoHgSrv0UVk+toNGh
RRvvmhi1Xf4o563vY8dXcxcHLErx60e+g171jUk4EL2I/epOal99R+c5/CRRNyMxfy6wswYDICoU
zB0RcNHVuipKHq3+hODANTnOLPvIvDHGHlt+w98l8wOTiY2DCliKwgz+u2oqHrR8TQz5cqgxND/i
Sye5HfsJb2WJ4QlbzUt/wr+YiZlHlOREUrN9vBLNQJM+urzZCfOxhoNk1SZnU0sQ7fd2LhlnKb/L
T4xh2XUYsAdCFUrR0UwqbhW8/uJiSO++ovfuxklDOjaMzFKBpGoAlNweBHO4gwmDgIj0YUlA01b1
n3C7UY3Gc15tdZwYBHsNEyzBvo5szBJ6AxlfP7jMC88rop1ctIRNSuO6PZdBOrqaWqfzgZNgx9qV
yt8807dBtFO8yoL0eig927Pu3n+nr93lFWBmUlMcDl8syqgMbHqPvH+6KONzCGZONjJEdq96uNbU
KTCApK7491kuJ0qo9Zvw3+OZHdAruQk/hBTETnWf/mcIzfY+VAAubL9EnyfLaXwyaqb2gGhADeEy
MNPv7qY15hGCDhxdW6syrTgKHOW3WaqVArDLe02W8aDJJZiFrGbN67piJkXkd8jVx+zAm3gpYYuq
LEcexEoyD2W07R8JLH/t4WqeIRlgJngcJwO5yOBf1CuMn6k+G9UtCR28F0aC44pEgXGeX0NdrVVj
2AJUtFZTQdsZnLFEKGwPCgHTqmY9/j3G15/Y9aGTgT516jgxgynk34HFJhpwxX2WJRNBaKchwD5C
t9kPFTQM91O+G0RgCg6Aqx9NM288XFmecPIZR1e5vZZxKWugvuJYK/XP6w5UQq7cGKQ9z2fqFm6S
S3WOQBXpWUIyF/56AcuYExGirjD+CAlOTKiOiIMtGC1DASJ5ACJJfFlETzJajbo/7HeNRPJNGmS1
Pa1DBFjzbt5/5T2P/KF1aaycQjjyiubtqLQ8hXZd2YPobMiAyA22rIcdGivomgX66nv+ckGwoWRu
Sbb1M4hBf3ruTGwjLinoH5oK9Ep91KCm08BXVZPHbltWpD8npHP+czP/NI2Q849WZezCLtIomNC0
wKgJVG9NINf0ly6Mt2lLlBn2x3AzejYLqwpzlreksOpqziog8c6Uf/ZbUtEf8bFtgh3OuUW1xjHb
fC13bwd2uef5ocW1CVlXuKTHC7txP6bS6rQGyTrmYxme/oN8Kz0RF3r3MjxzLbgy6guR4B95PHzW
L1R6BF/NZJNC1sJAyyrupEoJMWNcEAdpSQ7vZUKL+SpMsLp7rHwVcqKY3njeHzIbPROmFKzwDfJG
+H21El+Vzh8tlCXkgZRCkd/J6F/FLf/1a2fvtkYohtghrNP+0HruwgDPxZvBck8S+t1djmPdxr3Y
yeKpUbBO1Uw9HHh6h2tde/vwnU980/GDpz3p/SiaJBgXSe0PYkj0JEZqbcc9EP9C4f2UTMeKvu6D
qr6P8dCLT0ugZ+Sd/pwuWY36z+WbLPutXKOnu70rO/QvzdiXUjSnlX8lakRCMtTUAEXirgMQmM0E
z7to5qp6paINWVL0DQm244z6x/9sPGUllzHf5z/ys+FBCBCKlz26R0Bssi4BFkcAlzrtMzr2MC9a
+Ur0ctKbhR8bMxHxdZ4SSH6KZqE92r0bJOn5XfmFadJb+lm3UGEd4ds+evFNVKnfhdK0r1yhEDzc
2BIHJKSjkLZJInwcVq6fGpMMfnrWr5W/90mSEHdBel6RBC8iOGl+E18CI+JYYMzn/91S+K1P3ApP
zFQ2BppVbgSUQR30kUTrxMGDV3pSeDF/P6L9q5RMUA/Xhq/OqLp9BE5pwdB6KtfDgJjp5Y6XcDHs
TBMm6gElswNViql5yyvwUZeWkhWM/rkNdus/OcxUDuptnNVodZdlhjLGrUt7kKwSKCyW8EiGCOFC
hnxeIYmWwSHs8D3HZswnJjeqOSKaiHQKJ2gQUWCew3cTA1fPlcRcW2DNGjE9BTmlTddpOoaE4VYH
d9tv+TAh0a14h0I/vk6zu5BxoY+gsAZSQoS6XH6qaWWEFA+4bK1Wm2+o6U1j4jUkJhuA1j8jli3Q
VR1RXIKOtAwK7/O/kOfU8eLeeANGmC216mHjIuTcy7o3odzmRNZn/33H+SyILYXEOgcFU8neoX51
ycbAp9m/003WVGius0giBSOBxmvOu/YrRwy1IAn0ouLPitzd/NN3yBOWrH1ZQd5f9GIh4cUwQOe1
wMZe4uzWbnyWPimUQON0wHluF7ij90YJx+cblu/uFWmBAEHDfkcsurY9kxwdjopXuLMcDi+v6TRw
45pO59FyrL+nFND24vxncllL3lwMm8dstVHcPakLpYgkZHUHZeqmBPzgk5dQtO9N0MoBn+4RsjPv
Yg6+VPtf8FPmWJx21DcaiEjauaPzVtOm6uzfxwrlb+1r3Ql2dxnZJuzSP0dCLsW1zJJcwlFJnYHv
P2g28s6KCZ+15W/h7RW3yScuQP/J9GNYvxAkFJn+FMCdxrn2O3vXy9HcpRIDqNdMqxFTXz4MQ3t1
VxRqxxESoUwzY3S0SKHXqa1EHJj2fH8P5ZlqkZUYPQRNLIB0MAVTG4w47+eOPe05TpVugzV+iCPo
+rivbkhNnPhuNIrcGJIf5VTbHUuuCaT3kTDWBQSGX/rtH50FFg+lhoNbfkJo1wLIwd8nhuPzJGiD
DWuxp28NG1g6/4KjFLw86RiQ/gm6HBJMYO3IqG2skw4JWjaihPo3NZnhXOejLnveZRa8VkyLGzRl
u7xYRSZfZcPYJFBfQQBM6htxrxL7acBSd1F87q+6qGl1ixC+14ei2MPevApk2MjCLRSoqpZjGDe8
58cX1Y+fH/W9Trztc/EJ2uiDtYYd8OzOZjv3zj3ODW7wYxrBYz59elZxQk3PvB7HbcY2gwXbW5tJ
9JRbKZJlWrRMVsWwJOk77zH2cpdLHXXnBNVe/o6d21+kxiO/FLciSgTfmUGFy73+cECEHUrQiY3P
B2+59+WqgV9yzLBJltpVvRUaLj+OFzZTkG4eGZIURDPjdARFV4A9+IxD2mWb8kfqOvn56VjzfgFh
DGkI1BqMuzdY6wfhAjjqnDUL7TcBNBmw3Y1YrlDzsPo6Qe96rgLY3XxzSM/0y6JkpLzFKJ3vZ5XT
Nnt/u8R5UpH4koJkd+JA+Sz5dmqe7M5a5U9R85s2Ql66rOz5wm6/GZZfR/3fJu54qURiyDyMkzNu
3wslL1sM40V9XpMJU+wmgscdlb935UNoVROOYYbhnI83cea5vjLLP45ahSQabRIEVx1WIK0glolP
uYz2nAUzAYBvrzAU3PgpVqchuS46Wi/EZ6LRAgno86qhQ4dSXjdQvkkOSZsXBRVQ3z8Q2G066AEJ
x8pLlXjrZDVmo3FYJWvfhoSRqBvO1CUTRMFiIfB7kqnjEFcwUE8W0fvgDPmkJw37ANhyj+2T/ffh
y/6Py49432cifYm1BkZnYLFXOV6Z1bEqImRkYTQZAa4CieMI+QP3zUp0OqgDtzT42esX4rPqnrWd
ZwJI4JVCy/QLXqmRnoYbWDL07h5qOunsXtYT4J/T/McUqHFbW1JVHinRjEMLMs3un8J2Qab4f1v9
TmwTNRwOfzgazvS/vA+9va79ggAL5tZRC2hpaH5ZmJsxouMSU1WNWdJvtTIp12lI8kfR7XChQyFy
s5xTEWS5mheqnYB2EkgEL6OO1E+phRDFA5saNLGNFGieP7bTpGQHdDymRv1TlgjQzssT5UJTc8T2
ganujIpQYe4oA1/oc4UJUR16aYqtYFksMwI2QRfHKEg9BdhhQ1zk3uyqPG3MFC8F2K4rs8mwp/nu
gFF7v9+q4EEhbHLy6KO0Flymxf5x7iZd4VwYgXnIMwD03vCKD/aFj9EVaJ9xEB/4BUalspT12wNT
3W1lXx7BzzJ3DPf8zLgE5WMAwtN+Ibx65oLSs/mOm3AoPHeYHU4pwfYVjIqOk+xQY8bUfvyI+4W7
shkAG1rBGE1I7NljkpH+GlaHW33nCEe6/ZSUaoLS3amVoDIppcsz5mLMohr3knwfc3R7v6iqD/va
ZI6lOmUc6KV6UTTMBV0flDJnf8qMJUg9m5Ic247OLuhbcHbogu2QsDzJPG6iiC5JobVO8nnWP0Sj
L0Mx6IlCVFX/nJRPOuBjxRnhuYL0YPlTP2bkcpb29YBd6gMKURaMPITg8Dki2Rvv31ohBuSlHJMq
oh/G/8KNwAoM8Dl5b+f7b0oaIjvL02vgB0t5415YCazgpg2eiPkJZL9cpoo8XS+srGQV+0qDlsXB
0NAqwOS7KgvJ8uEtBXm6LUR37RSdFYGImw7WktBsrr70n8xAHvYXW84TrEN3ChUy15O4IRcKecX5
1Qu/RIajeBW967LkX9aSn4ZFojX7oB2oHJG2J6h9VuMKVacM3U6cbQCHK12N/uZEm0AFl/31eaDP
upXXCotARb8FlNkrIGXQwgVN7LpSwP0FXSL82ThROu5h/L8AzSbnbuNpeVk0zLDiGaGnYJ33OtKa
f8d81ciwWY6XFS3vf7DlWJTnfSawisk7NXCimDqYicIT2AnM2TE+NNGLL7taZqBnXiV9gw1FUTtr
p6FchxaVeuDa17LBSszXCjNF4koGsIYujfADQeb2I5lgdXxoBFac3rXg1hgxwPnI3tH9JD/fyLcw
LAv6ZuQsN7XZhpxs8+X4uEwm5jXKzQ6np5Eru+Qy3n6ThqlMjleEZL+PEuo7k4j7FVrkphMOMumE
SKTcgF0kytxZ2gxl6Xv/InR+GDqbGSa1e9oEmg7o5ptUxgzO/YxpP+YP2bB2Ll/k4/kwnD0gHIUM
ZfpcFGt8OM35qanXb3FlyujLWNRbFFZG27KrWLFJsQuk/e5j3QC1U9r4sUCesUQLyjbzGvFJ8Kfm
9GABBiZanLFhm2pRSBdZwGNUP3DIrv9tVGV0Ehkci9Be795cuioO6EbblnGok5CB8zPaTR48IkIJ
IFsemQFQmUWlR+eNToDkXi5G6yaaGfvPUEoGNHdxK0JdxPH29vWRVZ0rGaOjpR+RE3fFz6etu+/M
pYAacd3o/5vMOiU8eeVRNBOBNt5tVYP/Y+oBqREYclBCfS3kJXMNK17a5jI98ya1b3MXuWR3afSu
c5nUUSyPfACHJ6VBTd7G+obZjHJebz48MfKp4zTSv2TZ3+0ATazuXQeOjvd0m39DtkC9Qeo1kev8
DDQ1hMgK68ovqXUKZM5fgfZ2ZG5VNe3rk2IQbs4bzbwGHl0cz4hvmxAl7JKwe8GoHLN6OzAcLHGv
5YA5s0w+t5wdMJhEsXAUeF3I7FDIKcPs59wh9aWzZSfgSbpNSIEILuLNJlDd4nu5eZOAXKT+x/NB
Ny6K2fOTlz/TSSeKB4sXQf/gBBA/CyoVhvx7XQ+Pq1lJ3cfTwaLMsyEefYy8q2M69mH1rKKK9ygr
/AqPMWtmG5TwHGkx09PY9GTTBvKIKvGHWm81h/PlnKG7l5FdBZ9XCXRy9Ygg6HXvwVrNVRKWqpEs
IydlDemqDkM4QLxidv9BICVugmZz5K6QErWeU0feUkHXoWX1oUEeiRynPJvk6ehyObZgePYZN59R
iotrzcjkjZenz7aD0VvvW4VN6vKownN4wDJYSolfIKg++w7zHrFgFuoS5Sbk/CtNWfBY1Y9AXnDp
I1DlJ0oYgwLgXVmnMBx/E8ghzOP2Q1YCrcEYJoGOva2Ly0z56Yg9huzQRdiiR05O+G6nglN7h5G0
StqRXXRASTe5mlS6qUX10L91c/XDcO8ZFOW09Pwj8uSLUMMjXnd+ODlbpW538AbDheyInMYbQBen
krxfYOCkIWlKVZ/2Czn33NVBZZCL10sUBm60wRKt68ndsZA7MCKqWHMBoREhueLrYF1qrtxKEbcV
++58kjmAYfkCUZBYO7B2WL2qFjJK2NcrSAug9RKI1C+3UB8M5AXc61ltrUe7W2sFC463mN+t/ZLY
GV79DjHNLoOLG1mdC6sMZQXSMCOfY+8JwB6RvBFLKa/lbxTFzHXzViWZbmJYsgPynnxtTZf0tiMq
GIAmtD2WljEaVWIQIjuttGea+RcHYgQDIogk+zLf3KwfXQ7ymmVJWnp9oHQB0NNkwTPr0xiIAUZ3
96HCxREEaDBkLLLZ8YNlYeZ8uRlmlSnZ1ldwat3g/GuFXh6uA2hiQqZ5UBwTY2H6Jc6PVLMIRkPY
CQyGi03xx8R66FahOQ8gnGPrTpx6ildzIFo3s596Ma5azuhXkPIEDA5OyHCn+qejPuE63aV0F7SQ
cnDxidzie6v8MnVm+ppuP8amNer+xFgpktqq+40J5bOypwe54ggE45qs6MN8WsG12kZyun6pgu5G
Nc2Idoqprt8FPTzZqlwdFLznLSeqZ43g1D7u4Il54mOd1iVOo6mzPyxG7Xy8Yi7x70o7hjjnKTab
ubw6hAASgLXjUVrICMy+B94pkh4AdwgPgaEvDvILMEjMphQa9xI9q9g8hZyIIKQLkV0i+/1aa5Tg
9M46gxfPfbYIVDLpbcRzJ7ZMyuBbEMLCx16KYplpRjQgU0cO/QyhmGbllJDs6+FlTGXEMEZ1AZ6Y
ZOOI2az81DctrXNARgaX8MDAhwZpSEw18ecIuF72sKqE6SuignFC5YqIpw4rT+YT7hqFcTGveJuY
tDdqWxVWNT+53gR2gJE5v9e88V5yuTJK0eFq7uZfNluKpTWLecO+qT+Fj2/p/8QO+c2oEflP+m6f
D19kXUSdDx7myX4K5os2m8al9KK02VNRO/ayYN6idH1WVXGViFrc4LSaX0oCs/RmLAVRB5H5llPv
UGUkH17XpDEZajrvjkf0YwARV9t5gcNwv+KgKEDcbjGy6WSjRCIHjwwJdxns5YspkUt5G7HnU1jN
o8xUM5uAjxWNNkn3aNRCdpRk0VGIfKj70powtk/POQKqrSQ7cTaljeQfRFab0uias2hx5k9JQLHi
pthj3c369UvGIifJxGJArZhrV2Vu6v9IshAQv+ProRKXw0P0+QQR1qrcHChVX6wb/RsZa8t4NoTr
TK9UdRKMRtiBAsfgTRJ8pVrcsqwLWPmIbyNkRNvZHNLcbJikybE4E0ci2uBYWQPYsgE6oOdxlZ4S
6DajenIjNZM/aZFnlvup3hSy3RHpsuRRuCz781xKvL+qvdnxTcbk+qvCuyE9L6uQ8jPv6c3OAyob
N9DdqXnynpA8AYDQ4pKE6/b+Pyls5ug+hrCrCTfg4pOpeWqmr3BQo6u/4/mRFizb/gfEewujjEQs
36Ygf/puTLXMslf3/VpP99ogXjDfQlBx2IRmKN4KWhuqF5vmAgJvFyMtpGF7Qe7wxaMi4HC5qlp+
tIgbxo2pkD+7sDXRLhPAPSH3zjscecMZ7xwmlwWLn5DNZgRBSqfKepQ9WIhrTqSg1EZRjGu/P1ke
ZgqV3mTXU8DNNCtjeT725I2Bz6zrya24COgVRGWwuqLrVwgNwy6eTVh/887vaE8hSCM31oWjq9Wg
nCNnLGwdccuumSEzFAumQ4DOcL/xlu/udAWV1A2EvC1rU87jC4zHpt5TYH/Y66SLmtX7oxSewp34
+dgPG97to3uYr5LJiZUaN9cINFOVmVVR3HpXmSVP/VXBssWWFrZViG+lyJK0DowIFbr4fzWSJN46
DXcaIDQQfSnMP/cnSQDZ0qXQhgWx+fqYtan0jY3ARTJmk2lRVDAhHtlsbrx0VpmHSubIS9LzDjQx
wX0UkzjU+qVH8nisYEcstx1MLE9R8rheG4bQVb8Oyx4xVd0JtlNm4MpVHBxo08H/6nEPpdirheZJ
/PvjzPfuCE1vRqzrXTmZC8lrBWfyRd/n+6qAnGNY6I6Fi4p4cWN3L0StSto2aZHaxRKlB0+waigv
/LIpzphjDVqPQDftUkcxgFMm0fVi8ev9NyolC/MYh7xak3v8IxRwTV36YphLidnfGGrdX7HAu5KA
k8XYWTzAnZnNV8X6nHd7TEYPtTfNoKJ7R2bo7Mm58IaohAuYCJ1/RrOxikiRlP0EWZtg1sBfbHSj
7T4VrsvPX1CygXAc5xXM4DRJ32NHke0bdcFTxnVAikKey3r2Z4k9vqhGAaw32lOOfnyeZbvcyKdu
tsQiJVVdHFFdKRXbicbAP9XQEGIADrFU+em1QSD+Y97+GMvqVQzipwi/MdwDTh3A+A5js5qtsbeQ
eWJ7U6a7ICqOzZLaBBNgQ9MO/VeHI78IMixJrPDbX1w/9ZI48dUO0mJAjObp7aBPqawrxeAleZGO
nkWm6lU0nhFuGvBn07E/DqonHNX+ZS4KINEjpIkttXVhqwcQCsZggjAN8ISVHc7CuoMDT9An9Q14
EPU79aKJN7KieO3XmiGj9FsqTlaisB1HWaAfR+oGwoEHnZ2mBgUzxoIPkWO/i35oWvKvR2bEbHqg
+FfzjUnJuQeS4VC7R4/aoGijNI1Wkbea4gOscCthf7wkD+c+0wD0cBpu+J1gDWjgO4iE09ElcySn
u8U2pXynSrbmIsVSHQaTvS0sDJ9+HYwL8xnN51mWAa+bpqR34jIe1LftSMkGmMS9kCj5cucCBxjx
VLWro9lN7JOGeZPJmUmUzMKbADVyZGBK1MZRR/UVYTkcmuAKZePG4I2eYu/lGCe0f1gFaEWOtrrL
cTyUm9qVAaglmNxDEt9OUsnMSPP25IU6C1k66UXTC4gYy0IMHCm+RkdBdm/SieqccHeMM9/tjd0G
0XkTAa9jsO8rWcWFBWPk1wqhnUiR1EpisYGMCD31PmpPcA6vSOb+LxNzMTDgHoMgM4gliaJeJrJh
YCUJ1ILJOp4vYx1ob4TMB9MgGb+3xcS3LUV5wJbAzUFvvkZtu+tMy1sbJ/f5SiflwkaLPQDY9WKN
AJGVQkZQR/4RHd2naTa3N6os9nyE9tqQ6ILrXyajpRQdwFdub1ZiJP7DBpsHjeuUnJ2fGC0R103w
zHf+VfyoP01Af1WhXDsXK6Z7WCBSvHkzueX52kA7L+fsDFt07hNJBaxmOdAp7CJWHLOIymwsIoPc
VbUtDWZ6meIZVST3dmMkv31CAbFyzWNRyhCIkOI91kyLMVLcxow+FKqVRLsdhFJK/+ibf0tnnNv7
yubf+ReWCLHcuD7vg+Gxowu0tPWXCp5RxoinJ5HMJEqXrk7YKXxn4TSTY26Vuc7PMz9FAI2Ycsn7
UdY6fYSa5PzcieYUHsgiKc6LCg7MtfNuJ9O+B9kWeE/tQfUnvCFIqAdH+od56aTnVGxhaMWgAbJZ
fvshQKdwTAbRj1wm5kcpfI+8SvBhZuKV0Fh2wI2iFSejnCi1IZB42aMSkY0ZHu6PugoKztwhoBMm
coBPoa5XMsrvQfSXNUM+yy4i2fmyYnTCYXIg22k4BgkZjClFqa2XXcXMhEuYrY/cgrunO9Uim91f
jql3zU5CsJBsfEZLVCoUw0O3cw9qkJStJXYbS9SrAtctWUjIeBU5quncL4AhwEuxdHupZN4vEgyU
jZJi50HkJDXHW6kS+JNjt0w3KG6NydLmbEMFLgZwkBLpmhaWPddbpFn72jxZdDt2tTYCxv/rVOiw
KtDgFOlLWk+mLDZbhGD6gPOjionOuNqDQHFmNMffI0utUwDmQpcVsRxNB9nA4uz6fL52gvubYRbh
JoRlYTGuz3NryKtKx+2aKWsfx42HDNopiHm8337GRq6s4BTZwxyPRvp9tsLdGBgnenPSl2HWC6Yl
jsvYPqPiotSY31DWbSeyJB54BPjuDDiU06FaMK5bI1RVaXTB0doKaMwYrY65zsUIalXBoWG8o+82
TQuoUPYBYp2Fr6crywSg3oDW9uziytZWINyEvz8qAlky+qLVRxiu/x1Lug3GF4L9FAkJGmBfg72d
jmGRJXUJb2v1Y1de5gMdCWta1KPDX6Q200AgWt1+62q6TFHIo6vNpT+T969o0jHw0wZlgZcHJ+d9
mzjv3zB6bHKd+Z2UqHsJMVHxfSKPXLERGFhzvjkZO+twGB+Ou8Vio1eX8u3K7OzbpLX+CLJBkkWG
QwGKPDV4zyd7Jrupw8slQtC9/3vTPyJ1d/8xrWaCfkr9AmzpQPTh2qYDVMYJUj2Q5sFnO0Cmsz2J
MhtC2ZQsjx5IVBDofGeUoxCUgvvbGlUEmT8nmjNN/YxmwKeCZzl+c2MlMP2OzXweLoK2JWWNCIwD
l5cM3vB7XVPDKYYUt2eLrXZ3u6pdM7GP33fHbS0ay5i0FPlVsxlDLjgvMWKU8ujl8yAIIEhEfRsI
VqtLze1sY1jJg9BzWr/WGnsXv0QTdjypKS0H4cIK+GVlrJ7QaThsDeI/tDc1JfdrbJMtekfQ2gai
rLUhNcyKuLSzm0UbvfS/ZzaJWc+WvZXsvtS/QA4Y4OHFKX6NFesidxcvzH64n0Xfb++ReXhMtQoP
aopFqVz1SG/DyOSA1GBMP4jLWt1dYBtwXZ0xQDpuVyNdT+VAs16Fx9d8Ok2tfs4hHyKeshx54E5g
g7KCu6gv0WUtBivREWj1znDk8dtVdQNUG6vsXc4RDjE5tMv1Uz8JPfp3XgROZPzp4GCMPUFBtiym
pZrDwcmoRfFOGot9Kn8XbMlHBn3eRAljpQyV9muckggspMNi2HyvaaY/SuTB/siyKdDwNRnAW0JI
Aa2c8qPUqDBPZPB8hyui9Z7pYkVJV6rJgJuj6scUeSoAS9nY9O8KVkgoXzTlCJ4nBmuV6PzIBRdJ
Cf00Jc/67nqM6UA4I6qvaGq2jdIocvO1XfXQAcfCmFKIY9b9zv7zztaoJlk7w7klrW15POuMKbmq
8SQ6+GV0Burb78S6l+f2gaxm9iN3/uIy/qIzIz62xfMg17ibLHAAh9mUL9M8V7zhDNigsCHCBooi
DXIc4XyWbxdYPePoU84Fjwhxd6qUbSn6H5iTNyAVAkPmKkbGdEIFB+TlD3HNa2TxgWLgnOhugsG1
ZubGlmPsS/9w+FzCmyG3CM8M73/4pzluefjhX1B7KKSiJDfKGxNeILlaqyGVRteFgzSODa3/6hxF
xKLe5nwYdeVhMKhZpRedosv1bDX/EbMyPpp4PfEZquTKK0uNRMZzVVLlC/RHx6f2ghFpIwwkQwzR
A3VX/upiX3NMzctq2oSl6YseToD1vW4HgB8HDuJZXYmTYNCsVqSNEV5wCyB6uVb0LI0uNICeCvUA
hicihyyo/cMStkJoiTi35LPdj56PZiSPXpnqRoJGqRi2MfIiMgqEG2q2dqe/LNHiquBbO8BoAuAw
A76P6rEFSbEPEzdcZY/D02e2GQr1DIHaGTgQFFH0xSfVVQgRsNzOVt/J/VxhcYk+pm7QQcqd4evR
I/Fw1yj9bDTfSynVq0W7X8o3CvPihAcjm5U9bWojI0Tx6jKmQyE7Xee2aKTL2+OMFgq7c/WF33e+
LvALm+9NWS7lHDEisX2+NayrrMJuntMkhy4i3BwJz8WKBGMWO12guNRki2aitypx/2H7nCEnHxO1
IQLd0XCjPA5dDUWDwqt2l2lLIokqh3yz5f/Qhp095eNHTFE/9BUG4uVJsAmfH8BuESIExMNQpfAm
bO/LYQ9zbWMP0BN63bSpoVp9chUPzHKgD5IGA6Wo5PuGJvju+Oes1iY0FESnyczXaTKkJ4JyAIua
QA5yJW1cmH2K7E8eUCir0wHrqQIPLIEu5sICfTL0JONPH/dNf4t+uibwYEzS7v84OH9Ud+Up4Owa
GSdGr622LW3ekAOSvL0J9xStZ9Ht0soblTQ5zYnBVO1F2MDIaGDtUHFZsSk6MrrjewoLFDUDHoba
PtkSxUoEK8+DZEhPcJvOZv0GxpyvNrK4IzSST9KleGSxvti1kGH99aUkeRTLiBRTzbCDIo/uXgW+
BkCUjihtbFXBEqL7Wlb4z2/gy4d1PeVdA38/mjg3hiMi2ejNAu+jYykgBnH42L800P7QVPcY2+jt
G7V/XeHWg3Mu+Y/lKFyJYNds8XouWUUrfB29AAX+oC8Ec8f6jzxepv3zI/xD/hcTgGuAx9YxB0Np
OIQrUW2E+nHy5zhxJPdJAQsdE58d7WoA6Vk19IVT3MG0nhvIRTFCavpyS9DXowqsiqcGE7+U0hhl
SPJEAI0KUNc467b0RH+rhjU4YDTdd4cSGE0lPqfWiX0Ui5dwDo4dAGJrYhsZ+5iBs+RkRx4vq9Vl
9pAuBLbSzDJbwMswK6opV5a9qINrtbTI/Hb90EqX/YXE6FTPuJ5NvrADcfYSzZmQs00l8AaPnwg8
4g+IC+ZyoEOiM0Wr1z3uYtcfhAoOMt904tKv8+CbPy4g83u5wQoCHshF69Zq/VxDsXi/PRrw3u2M
cB17NRu1HQaHcWDaOpod3wsNu+Y22c/MsYiTu43ABRxr0cKMzMaTvvT8Kwr1gCwE3cFHGgrZJsIR
E89oUJ6QawFqBRC1xuGaHjl5QTfb3wYtoP3O/9bSGme243bQNOUCll3A1+tCq9wpVORmNHauOHp/
ce6j6C7jAIqweMp456NOpuO7c9d2KuUl5Zmsy2eThUFOSM9VkzJ6WyybQDGFEuAxR+VFuV4PAKML
qQcendFqzM1K/Gs3IgzD0jPNh0IxahvnGBCLt5UIWK+Y8r8odpdzUwNa2sjPXtHIXfkY1TeRqnqY
XHOrrUUQU3xi+0uToGYg180N5XqUG8k2UBEdiDheO3Ulw3gMaRkbs/FTrrx2z4d7af5QyU17yOI1
lk62riCpVQo/2PqW0c6GwgnsfPgD/TcN8H4Dv8F6aaevFvdr4IkWtM9XEoeqAYpWWnJ4MyhnKZZq
Ii7C3Sez7lj+I74vSoIMA8Dyds/Is1f4tMWzzO0Ie6hHrqJIf16dLA1bCMxI1n5IfrGdFcw4An3N
HR1s0Q5gD02h2dbILwygcGeY6/ZMgRA9tQlYhNvDjTWO+AHmExSz0idHtlOgSV8D0E9KWt7jbII1
Jeamojc1olrnc3YVViKTictWNabVsTRWbQ4ebym6aQgIvpr6yKl1R1T+quRmzGAU5/8EShbmtLHa
LedXEWVe+7ow/tl6L3whFo6bHZClaOaIwZe5Yq4vzkf8fQM4Ctjx9APZOBKYloDqK6DwZsN3erqO
p7y3gSlmfeTJVSz2JV7vtofd1JRfkAZmOxjNZ4iS5Y/UkaZDTvx4BFf612Dbbf9ae+VVzsFr2NjN
U3IsRolMej+0mjSZYu2FiUa5rSAtBADtgIZ4Gs+IuGGw5o99243/srGELxUTNQ3Hf2IgMMSwLm0t
5wm8j7taeJ8PVS5tjU6r6XpqLh0tKiXRpcrrQKHrBh7E3e2KZnootPIO9qG6bR2ogYz9/IG+ivkB
1wwPnaFIN7wMLJ/EyV3bA3h+jiW7IBNnEaKnFb8OyR77VWnQYm2im4FQgBIRhCxpfiiu8JH0CVC2
HjEhF3svKG16+U+SP1uOcfBP5yS742rPf5wj4lRssbGDQbRAGBmycwDkMZQYWGqY78Bq2A+gwD9x
vkmMysVFzq8ChC3YHf/Mt0RYJS9OwXVqGIO447CvTyQi9JNo7bueERbxcLEkJ14w3V85ZH0XCkix
xwhrXJ7C8dKsDBdH+MO1WcPkvh4o1CczQ7Pk5/lCtSKSls2uK9BxM7erGZQ7BADa+fvObVtwXX3x
TFN2eCpOi6u75Nrq7t9AEJ/hZyGYH40xsgkwcoWIcQnFJbYjNw9o8qarBsyndfYVo1/5WkZOLnDK
rG7SpGtJFQWueyBJGrApMo386PdH8vr+mF0FA7eZidLtvGkLzQjjEIqPAyG/NDdxaA/29o/fVQ44
FRklh+jclpr2g83Gq/7M6OiN/4olIuuKrrGH0CXvwBDjO5aS295ltfskBOdRmtwu3l7b3mKN7fdT
J34hybhvpwvzS/BY2v1dv9BUSxgc/y/lK2y8Okg7M8CHc4N9Y+6FbM4WYxSKSnSwPORX8WI5ZX2G
B7BoGbgGuuCBQnQCc5anMqDdq3A+GQj2IfV6PEJFIsTGhTkS6Sd8nkZZsbcWAIsCQUe4YDXIYWfF
357uNeXhJ11KgC+ex2v+MJr0Lo0DvaLZuQ+6FypG05/QZ0O4/GtvcwvUtWEdSWJGf0yIJ4WT3Y5D
P4Sf3EzZoU1mhPuKBwS3Vp311LFfc6BHj2TBzO4s37rPWZXmmqGGKUxCsh3TVcp9wbD8XozxbfPB
r50t2G4iu6rCTFPZtZUG7L31Q6Ssf02GxPqSvO9nOL6musXdCiiN31P/3OBRPL6dnFXOLm084Stm
oEbxhO+Y8WG7GJz+EhNfTkh2zkGsAkpPqNOZ9IcMu/LNu8G8YUmoSRL9DZFRlM09BOyX3/LhbLCs
VqNIF3lqPxaC72MMGQ4HKBqOcdD8/1vUfFfbEzsKTjexbHndp8PJs9W9tqQV1+syDJq9Yw9UVY3i
2uhxPbLjmqaNYAYwgqpKfwZBupuS43wfuzyDxv97lnEDdu1Th9mbfgWZPMESQIQE6sNhlS2pIUfP
nBs2YTHDBYuxGQoHL5DECtwwd2Wjk9tsdLRxQifKo0HDeEQKtGbxJU4cILhXe2HZL05gvY2bTdFm
pUCct6k92q68bqWsSe1T3sMOL7lrOEOPM3UuN25U7gFu6vHSaGuBHvxCu/6YOI7sCGk07yIU8Khp
WpJX5yHFf4RGPfo/g8wQAViyMSozUkuc+g4DvCjjMeBD90GTqGW7l+OraDEhkoWXB1IZb1+nDvBr
mPF+54wJNHWGq8M5n9nz0SQzgEToseWPkh1w9I7+Hv7GiZndwFOBcKEPCT1vOM1TmnnDfwowjcmD
KEBV2PmekL7xmtMP54Bf17rAVKbRiJoT9gOii+z2sxnjlJFtv3PhN9Rd8/5JgFpxG1vFMtGhuVTl
wj040mtXTgMMhY6F8+JD6zBi8Jn+pCl7I6VP1h5Ch0j27aDAkV05TXXElBiPBlZuhi0e6WRPjocK
MxoUqm3U3OIpQmMCQovAWw4ibgfKQfjv+8V76HrVntQj9ssa6tFR6S7mdYiRgKozjAONxBrs3ryn
1a/vsa4JvyQSYaaHX1IjUeRiG7znHjgH+kH8UexnruUnTdvRUctbvEDkBlvaFSOlnnZLuiiQYPLl
m+Hdppfz0imat3yZuBzR87skaEG3/UUhNtcWgj3Uo+pLdv2OnU7WNrcFEbbO6gJ3pkKrSBQtW3DF
MtV0gF0d//9m0uR+VLV56K9DQ8zXRjCWZWGN8Exg8EsSMgpr2jfu+03DgcJgpqJRauSpvSIEcTSm
IuXjMtwSXXkTliCqyo64dXCIfTSmVo8jmdSngudhfJ+vWLfaJMBSm9w2XB6au/y45bCW1rf3O5KV
JWCVLfc611mdfAelQoYPAdfcp6Kdt2yGsXR7YUyBINODjDK8fqguwM3soCba8xybI+vTIhocLUEr
I5I2dq7LeCcXsMpPbPiXOTd/eWaMIZr/CbuotwxuzzZMNEc9ZDtZELQiP3BJ6i2Ky63xrt1GrMIt
yUcQ0yBDYI1i0Y9QigVdPCL0Ggwpseewy1foSfDtOCRITjy3kefmiR5J1eDzWwLDWGW6jwsT2RxE
IHiUAjTqpUlFB3w14A7gYE+axmWVlcnYoEcFrMtZBLN2ITCXvmfmY02QRZTdaXuwpS1C8LrTg6ZI
AFeYGQp6hoEht8+6vlGSn3Y2DZSAhL21zhKnDUF5ocympdu7j9PIpXC6W1U7GF3Nw99KhyMm9Ulc
tgA+1i8cX2lXtpPUu65n66SevUgz6e1H8+k76znQSu5Uhh3lnkkjw2bIgECk+s7fT7+N11ynxFAb
OCVhF1bgfdufHrqmoo7HSdoHiLV8xKIDQ05Egc6QbJE2gBMS4gP1xOwNqIJg5/sN/VoPh6ZIfu+Y
HItwvQrZAnt2o/L1AxUWym0Rk5quChBeGy2tJdzgkBCgKZsrRIbI7nqOfWIWbM1R0e3LSabO9PBo
RiVhHOhgP1lBrxrWGUfZAaDEMLEVl2FfiEq+S8qXlKWzDItAbp422cotg96otOsRoPZ7ZZUpdOTW
TW5HSWMYpfjXj1iRE7gbYIZoe2+QNsmrJSzA8Fp/rrncEcJ67vZvEBuXPMGYGviVMPUX8QbNP67m
rewu8ZQlYwqks9SEYzrPR/HXB+YQNDWTO3OA3tggJtATJFU1e+xUt47vcjXU9PH5+g537oRUCRtX
Hbia14kstLmuzsgo4gfHo6beGFt/2ZW0H3RoqL9vMKQA0Y5xaOGwU+NeUq6hkLmIi2W1JXmnqLHR
SfJGAs6sBuLPMlb6uymbNvZqnddFWb8I3YU8TtoEKI3RlEZMltTQP3rhHF8YWCjwmdphsNvHA75V
3byaQXE7q+UjD7TIOjeTC1T4PkLy9jy1fqBi/jQ8yJNP7osxMKQ6ULfd3ThoRzZygSmg8sIp9pv4
HZn8bKuCsBia21r9+FmY1Ld3UyTpqUvbq9jYKYVp0PUcVbJGSyeloXXbWJ6BEP3UW/kE9HGNme2Y
zQz8WMmS/53E1ANJn3t6RMzTlxMYf2/D0/raWiwiT3LW8/jr4oLcC5SaEHyxyrP8b++DFRzfOelf
yDJbI9wEcEIm1B6mk9mX0O9FPggrNZDIw6uQmFjb98z8pxd70Cs7TjlQjrtLUbw+IOeCpbjqKcwd
1Z2C2pyBtt6S2Fcc4cQXcNbMjZ3ra8HcH6swUkvGTXBft3ey8WY3bEnuBQ4xzyVTzQEO2QN94FnL
ZzGO3Pc5oJkzx/vTdpnz0uDxPm6g0pjfxg0wdmDZKv6YzSXyJBaO7f95GWBzWHxxdupzqGb0+WgY
ZUPWefABMC37x5Sa98fdItfWGjYdxBexeJ5BwaQobUfh82JKvqQdpLEvCWRvkN2quy7Tn4LK6K62
QDX5Ki5JbuavS+4IHYqt4nPnsiuXqxVTCYk1gyzpvU8ydtMkNKi0yXPhb0OnhsSo+Pwrkeq0hWJs
osx7S6cTZLbyT7L6qVTAiww2NZXsTYpPj86ha0BUTSDpMQVwRJDY0CCpKgkHRZxwfmeIvN4s1Myt
25Ckkx+0KsEz/hJ+SnIWQNpGEs9Omtght2NxngBPEtEwKOK6JM6flK4f4MeZM1AsP3NOhFUE0U0i
vVhUj+YvtM334cBpCRDfVwW7eKnVgAd4i9NG305ugSNX4QsQkxbtPti36HkX9ak8FWqZxIDdvAXa
K3kUjUT3+FRMT67iX4NTAmW/NyXyPQ9lck2jyFAqOjtU770HOQuYRhtqO0V+b5xcW0JigVAFud83
ZmZBXZ93ikjONDZc8JPEx4ECHuIDWBuBRqu2pvmNMQfKtQRwCoyGiF+n4+IAVKmv20jLcKXI2JoS
nnSMjzk2LGRGyyoqAneqCeCn94u6dyiA8caxVW/Mrg1bC/VOdrXYM4X1jtvz3IAtKYaQIDbq+Sjh
D+l9aScaAqPvXHbjwM0oDacvei/bLtB7boNK+sWN9m5h5HGqctcWZSmGjWjMjP3+xIEfV42ZcAyN
oRe9L5oLldWFP840Ow57NdaZFg7NxoEoaxeDxhm2ygPSdSYy1vkfrE3Gc9wUUhMMDHdZ75wcylsx
pf6qSdOEtXeHKy1qNe6k54Kw8c0DOdHAGdAC4vJn9vSNXgF4dgDlILk4KTV76qO3V4lE9gWT6CaF
aQ5tCbM3h/nATNnpF7jwdUEGTY/f0Dkf4z2v9PBuY3MPth5+y34vInINU5CbvNpscCEBhw/TwL1y
Qc+KawtRG9+hJGU/h147x57uWIuJxFhcu+XNn1+OF+NXcO39a8SV0zspu75QBm51mjwvfxaaV7oY
AfS4LCW+mUGJdHAHUvBGcxAS+ufWeRlXW+UcgAxUfoQBzlCMoXnGDGsP1F6IbklMrMLZ0tMw+owf
51iJ4uhHUOfXL6eYUOjvm9S1Es0qef+L1n+jks/TsyztHd9XmYSz1v4bzIZN1jtCGxvekTtMw37V
TidIYeNbfZYWq0wDjR06MtFDzoApXXpCd/ndEA2tt9FYMmK2It17f93gyiDIz89jJc6SKfeGJ9g9
gbQyHOXAlvQ9SOuk8gdqiDVs4kXArbp44jF4QS2ViGsYHE9EIBaHoKVNtM8hBwwSF9YyGRF3GEcs
JYoPPiy+vI+AhiWPJDbhZQT3dXMO72+OFhajVf9acGOYQ25kuVjjPyuCqaLiaHgauN9Y6I1FKQCp
qNH0tEZFyiL5m/NQdtrpVXcW661sC1tz6IcZYZpkSBye+nuRixvczrnxh1BcpLlJi1tnZM4TpRnR
dnEed76PUZbTeuJhVEXsDMguE1day4FSBAJ0b7wvVuqOrL7HMMubFVP7kQzyTWfGH+Ox96QCBYqC
xw5Rbk0YXi5GkuSL7ttB64wqeCKf8qfXVvaYqEqOo9H7QSSRbjmHRYEpRUMz3S0MBSWPK4KfaPs9
DI1lBpFdKd3PZcy08yGeJZk7QSWODWvq3Z9Q58ebuOMmPzaqIgHwLYGvt3CafjV6WQ8Ela2368ci
aBWs2U/2wZpqmApyWNUmnmc9Tret+n1OJx99E4a1fvN53Fj8ggY0mr6uJtyWFwLohCdH+sbg97yh
xY0Y3eAtPon+cI56IdLj8SQzzPqlF48ADJXLLzL2/pd2VTF1x6GYt8URQ+SGlB3hJu4dqk2qMTDq
TkCuRPEy7dx7SVEe3PonXTR0r54r6kxARfSTcs7sEL1HeFOrHHueip340NtQbCU12Rkatmb02iRb
UTrenhZsewDn5e1yOPzuDhOTcIvKm/m581GjPt1iEPOw/CK2pXbswAKlfd68zUICiHpMr3nnhX7D
KMwVdi1pJru4Wb7OtXN1PU9A1LGCy0rWp7yfP/eXbnyh+e+A2si8rkdWlF3fF7MImUGZB/5by8Er
xvcyA/jYjfKZD+yB6dREwK3uFgXugwDvBc+YTgD4VG+mtc9Wx68gaaOkqiahczh2tbYb0MxmwJip
U4Tpe+dP7sGQTmkvFW5rLEan+2NG62b9qtYxMEr8EeHokMBz2hJ9kb76c7bhb6ZKOt6JdCAuA8It
D9Vs7VdNdrro81uXuTS02oOHvCc9/c4gLejuvEmiMcVEHbct9tDh6Bz0KRwUzTp8h8ZixDimLC0Q
ApJMI7RtuXZaMxJ/72VP+huyVNTXCu3IPB8zNbuCtb3JQQHUgvAPlaOni/j/LTJ8hG/8bbd5B9lR
7ig99DTM9amahV7NaJ229gl5wZei9XweN8UkCyd6Z3jGeblwt8Y056HoRONCk7UIdJPMnzA07oyd
FUWBuGwIBD9Yh2WjbKslwYe9tGvnrSRin/Qc8kdALqESySmlBWwDnYKkhT1GV/5Ppb1oESQwhpDU
frUJuVulADLRaROEoQ2wi2+OjGdzppzrKcZ0bnwyOQqRzK8ucRPb5yPoe2ZLpfb/aGN+4idlhhbf
ISTn0/MNSnqM+arlrW/cLXa5gcB7LeFFkz/S7HaRiJaz6PYzpPWa2uOJ02IVKDkA7LQQXyHHiHJU
dPTc2p4kojl/SWNxx2nI0wDf0XmLni6F430ormax6NnFWQ3CY+qSBiGLuAaSqo5dYi03KxWpcHKU
MgoxM10GuOxydQLBLIDyauWMuTihI6MSSI3mzgi7CAuI8vUeLKO4+jye/cWCx13tmDLVOCc8mhOT
1o/ldwE3KyWmkkbUb1Lu197Xqx67oHzWMuuvi2RFHi12MMgjzRww2uzfXV1LEjx2eCwHK93MxU/O
SkFBkx/3vlassTN1rVziZGyWbWLnvmZ4BevQDovWtwoCVfSSY6iK/7ugM+IETyPbNU/CaMJtdBQ/
cqIkw/xwng6WRriGENXm03Bl8p55dSc57RTlDxR7Dgh1zeWUTgYq4O/CwPSEe00tUSX+N3bFK0Zj
S1SnpMVOVMSfuKPSXMCec2x2+hl4it8jnoJxsEv9xMMG+xbIYOZkux1IlxqmQsWRYojNNxuSn5Jj
k1H/Z4jr+2xvU/sktwAEtjoBdn0Hcewdef4HjGipMLat7GUk3YKpQ9EfALaE5fxPalFjTZPC2Bou
yg0mrQvIyHJsblCTlfFSPIqFkG+gsyXqDJXrIkUUjevtuV+9n0rmN0Kt3pHQ6PO3F+96r1P2DjeD
RhC/UL/UmX09sVJCBFmj/Mg4DY19gorQlqrXyyMO/G9gJox7sTe7dK3sjcak8oXlpPtkKZVB8X7w
f7zkRBSfvKvlpX2iD2bxaRY+x9whbocyx/uUUWUTF9P3oOI0/s5VrrtLU2nhEe3EmiOuS302H0yL
4xodVb/PWAco4JrOk3vCeaojO/cUHKJh8otIM6s/YLNPymq/VIH9KmunuhjqdgqLcAPlw1M83Tpr
qaorTIucUejytMTTFifx7ZnLXdkW554j0sT6dn2oNaDR88eShpaYvuOcl2Q+A6SRjMTTI3S173kx
74d+Iq/rzMRjltuREsHND0eA6YLoX/0H6FO9LnVxMf4RzZFicwFYELJaQirZMmZIXmMY/eltmspH
lxMl29lE7uluJ3WQMF0Zqjam5C3IBKa5OPW2KC71MJykUWEHb8MQPIdpAH9GHziE5b6sfPt40Ynn
TGSzY/oCsSEXw9nRCVVRivExMt2TFJuReZJ4g52Y8WssRjdJPFWsDODwnUjXymqZORdFuQSN5Jvy
TSgQDtK0aezMZmqavvHL3zRv10301RS+UH6BkVNyOeTJcdJbFgXk68800az48n9ItImiA/eMniSZ
2yDKFo/t/inr4+PidCiKKT83gxn1AyQIT+okkDi1rBfKB2booCAj52JR7bLEyGrpC1e01foBXMvQ
qGMzCN2hZ1ZFEjPSlT6YVIx5cehShD3LzpUZNMh7OmPzhjGfubPuCOdkNbCv+Ez/7oVxEPaK8MOm
kWisOZ+87XcpndFhFYS2Us0/bNWkvcT/sbJEClp4PIkwpn7SL50kJehBMhOlmRXcMR0RW2dD+WOq
Lc/gqWENjpHHT9qiPm2iUkAbxm/kg74xf729K/Vlqap+8VRvk7tqzuv6HacTk2l/hox5Xk3gJdGx
JekuCA/GoyPz6DaP/14ndALQa0jeX+72aa3HmFl6PenVz2DpH8llMuMySyynJvay78gCQTfiwhXv
EMMtWTWutIJwCSmpnZGzvp4/5NICkEZSQcvlwQABxYC9Sp7eEkAYJI80BoZAD5xQqu0FUnfahYe4
hXMD4Eq4F+iP/40uj05qdsEvU6mEPR1cjh5GjgtQm+BLY/5vBSmK4spJW4hXUgQwIRJpxQ4Y5qvk
Hlex53Ux2o2Sw25kG4YAsGC6JqbDNhSauQ21OsToYKVSf20gBk4/EoEAJbiQzVlIQ0SXcQN6IEhy
nnUzwSLccppzcHyvRDnx7nVuVJ+8ZIlI0xUVr8ovig4AURkB8MW3H5WguXmUgl/hngi+lWn9jfo8
Vk4GetgBwIx/tUFptCGBZfSt1MMrJIb+uuW4/IYSwO9Q61PG00ll4lgwBwEfNCjP01sTceXObROm
k7mXRyZncIZDQDZA0OPPRYXgPwmWwIwlABDGFJQrs8j54PkYjJLIBbeO9HEl+DPekFAzqEPnG/Rk
fhzALiLQFcmROdmIHFlSU0Es85ulpXnVaVS8MvvQY2OFCG427vyISm5s1KyTouXTacXISrk1J6em
RPpj4Upygt9G/26gdOtELYtp+zJHjP7Zk3LrPBSkqX4IVhPBNOCq0OcLbztvaBkUa8ZjxzgrGdTm
qU6OIU/CAJUsJSs9NnQPP0b74ZXfl+FtfYB9/hXfmNtW/cUJz71m/mxZieu/rDNx2Zki+SKz7dEi
kIa6hynpB0nRHLlHloJFCeB9VZkAGz50X+h0evAJFm48jQivue2xZVLorEyNGtKe8h1bepdoNk2x
+jElCglzve0xZz64v7UYPTkJJLWueje07UD0RcxhswZm7xHStLAHkc0E0ZABgbS4JHYcSMAuBCLA
Fatc6WMxx6GhmYw7kq4/HN3FVcGlEUbvelW25QIAx3bqE7yl1fToxV+9dPU4KWuBAOKtefA+oReg
vZWTu9Y0ViWr9XNrGtJzSijcD+RtxB6N1VyQUx3CLNV8ZZ3piPE+1SWVMP3B7RaMWpVODhwrJTXN
Gbt14hrGyU0O0UYdmf39OurSULLlxpi832C75+0f5uL5jqiRavkwZDii13tdPokUgzpUUO87nC/d
LBt8XmdxXWZQYC32OQMKoNlW/StAHou2F4IvbUsWIiIb1CFRWkKCxZqOog+3w0i5ECs4iH/a4e55
6x2UwcbzAwCtBg/O5V7MI0X6c0wTaN19R1SNveMxQ37J6FgyY5MzPafpN4AF52je2Y56QrVP1U1o
+pLtJ5GTNNd6wZFnhohiQ8hwaX9kyEwGvpfBODShyxMj4MPZqKqGFGUGSLa3i3ETdnTd1GwZCfaJ
k+eLOkX4o/bf3/5oLrGrES4MoN+f5yEtor/FWN60D5xc3+pU3kxkRQ2OQ0ysu1CaFm3PxnqySnnr
yQuJ3VDgDycP0Z6WallpmsJv4OWr2mB1asqEMbtKWQqerZBPjY7MXavNsYwPYBfo7+ijhcAatTUw
wBYqlhtP1YamhgKuHLHhjaUSAWXneRqF8VfnR70ZyTbIfSiwvDCIaXCxZPrUMeUYIn6vDbyJINbx
I/nSmr9lx6EpGa8BP8oS2Oh2c+J7BeoG6K22wrBGw5TdIFFjVqISrlK9zYqQaBE724EoeBd0ZqtG
oqi4bXmCaQfE9thhuQUypmMWgQUKVjJ3htbJi2L4bX49T+BwJZMlTLLBGBbrvrHdToktGiFlYM1Y
dzGgyW45TZlMDEzg0f7//K+CMxo/tGN4qxIz4E3ogjQFdZ3oHaDzz21b6Iy5FJYYz/9bswMF0dOv
5PFIct91ybfv/ddBvmcAJgIxvFugbwIQnxBbSHxZSrz2Ro1oMCI3VXL7QRhu6SMPMjjNzYAgvP6q
qMvcylHLYxgX+LcOcdJLTyxYFtZntBp8N0BUMqgq9Qedns+Eigb8X6xsP6Ra6HVoaGsbb9KEFUAr
8j1cvsHW1MDOGcwvRS9YfduL75acfjfVbzh6R5+VDUdhjvSSSRnv4QwcWoRfOGR83yrmFU9K6LMy
lN18toWzXq7rFjANQEIN0RRN6x63tOIjwJ+p8RXDd1kWI3eehV3YTgo/1Gy8M69NHmdzMGOfg2WK
uXGxVAundsnEA8mRNSveofYyujONlYw4ju+bmUE9zXk5to1SQe2dY7Vc1avPi5o/zOfnQ99bic6z
F1NHtqzWIHeoH2S7mSvVZFVLweW5vxHsc8qWePpZ3283JWcnrZUOlXB+O60V6Q22F427yfHabKdA
vcuu/Nds1jsks2TuVjNjq4pZrtdm02TqGYWb7gEG5ixlBaizV2Uy+c4H89UvjtHeSN5La512Kr4L
e4dEYGPDHXk3XqoPazGNyB9hkqioRkrPDxqcGA7ffd3yqtzIT4nHNzPzJlcgZlOPgPOI+B5Yo2gN
I7chDv2u+iuyvNkXyrBXVvWagOw9QQz75qrNCFNfsGHTf+cZLSqg2Iq4eU99R19SEKXKao3A+H6K
FYtK7f5eV67cOOLamVyoJ0Pnv4D9w7VswbFTXeDOG4mp6H1bXlY0bN3b26eaE2l6dQzcaiiBVnvs
oTvOs6E+idYCNjRtnZOE2dd1CKN6aXqpJHP5Om0Fwq2H58Gd+sGdVGNIlrhRtT6OfltRYr1k6kk0
cV2ue7inVUUkj5fpN7FZo5qE4ImgGvjI86DXmYWKROi3U97nV8q+pJ4ZvZMQDbNxu7eirdjpDdte
fED1uOgrzsw4USZbNuGBgBRXXwjB0rmksD/h8220YGHex9U/RV97MNVF8MXeZK90p0BcPgtKWR6f
VMDVrh9pZ79oRf7kEbqsLE9aZ7RJDwdXDMP8ekJSMSoRQUudTw4IqdKUv+aLXj4bDJqPib6PUhs3
3negnTcFMWm7/b3tUIiUuqFyiAodAeH8Gi3hYUg+CH7yDdTLgGcq6trjXZSgkKR8DmWt030eoRTr
3Nzcg+zNp4I5uWhuiTk3AqmpIDhsLOXc4K91RjXKnxQWpcr9UIcs8tZUpA61kVa+TkjU1b/gqDtb
JFppGsH9YwD9A4aq+nNr+WAtQdQk6S6k6DOxZ3TJcnFppI9YNFq8mQk4HM8AIO8wz6Z1KHZqCOkc
2CbC7V8AoLiakg89EyA3r3xUSCc6FLvK2tU4G2krwYfsUjhkaFIOkWN/fuOcfD0HlMINA56/dLsL
+nmZso0GmHxi+qmK2Fr4oqx57A2HJq/h0xBqtTwz4JuO/HV1YNuXrdeQ1Wqk+rMWODpLnKyVfbbo
87q9ismbzoOStxB78fhZuc+q31C0bv61WMb/mcqH1ODn3dWuNa5DuMk7l6jobGs8klWLDXaTTsk5
CQSzTnqKi1Mz9EvLecFKZ0toYPmBSE3pmqxK6rqOs67AuLau939FlwAJ9YJtRJofZxvxzogkq0W2
Qd1bbHn4ymXKh0Hv3uwe1YqJOM5W0KavGuuG4CKnD9TEot0Mmhhgr2ABETzlIiAEr5mKx9dB9Rfy
yE6DlSVo9TJcjQP3qb1YU6WkxQeu3YfvnYT1khypclyXhx0VF4SKEEcg/7phrp49mrKEYU2kKjzi
Z60HR4rmIQzWoMlkLpVdW0ifE33sm4u3CgCRzAbY2JZzahvcigJmETri+w+/938w6DP0BZSoSfgf
TizyGh30z1vcTBquB8BsS4Pw9IRwN0rseedb2omVAVorJb+bO+qyaXNLWgWnTQNeICFJWUg0fm9I
u6eMoNddk+R/Rr9/iif3d/xzwRj8N39SAmzsGuavTYI6FtlrE/URJmDByc324mjvR42u/BYFegmq
N4/jHu7K6j/Y63TlB+zwk8CAhPdW8X6dbk3U4D2Vri+DHKc9Auk5EuTmxk3oRUbW9GtihGN8KlY7
GNghRx6BwrfHltL5D8tgcspI3msfhPYeQSoCRrrlr9iCRtEWy51aamFxRzmv5wexSgIEqHcYI8si
oHxuCzvr+PtH4+tjKVjW1NqCVUNsfy+P1pGJ+K07eGoIF9i43kcxxb99B7aUhzv36VJbjkA2ANzf
mEaCyOyOFBVln7xoqsZOMafnehuPSSJL3zNLWtDljJZOl3/fDUUZpeyY5E98ncYVGYvXO++3mJHN
2xWqTMsZ/fyzm3MMUQrUic5ZiUUpo+W7cGNQtCXm6ha8AyMmfFmBQ8vA8EgApFIonxxyZMxdB7ip
ouldXHDgBKpSRVRRu1pAWLHDRpcQ59X7WSoS+3uHi6s0rIoh2iw43/k49otyMhtkiYKV68g1wJFV
eyV7z/D7GHOXp8PyzKSb6lPl1Fn6BhCtJa0HewPkKdGWKEqPVk8YzUXcMDwKQxiBAo6M2rKioUvO
swSqkEEAKw1XzZqUNv6hc7SpRd+iErdKGlTANFYYsxgIgi6kxU4esYmV3pRDBUGsLZjMA7jnGJWv
fSjGQxL1gmhSAIm3HLLCTNEwKQtuOrySfxe+jjelyx55rcUyoOLMB+aJCPqho3hL+IxMw8KXGoWs
cuuUvREXoGA0ZDgLHBLUJHx8ytJTdhrsfFqArub1OCa9FvbLUZZvjc20hIh4M0xIfVHeruH0Iq6w
K/O4GuqT9QTKqzcdx/gU7laxo+m1P7Z26sezImSkpn1qrgWZwVh+Rg3QxcQxST3BSTElwFbRu31T
9hGm1YEsmv6kgT0Euno61R8tTaLf1EYV/4kWN5rBKZQBUFyQArvlwTfleo9H4IczrWL+A+6XFzlg
8k3e7xgc7y4ZG1tde5hxgj5tFib0Qd/VYQJdigUaQGxG8rOwKfqcl1JmSSi62zKqphXatBDhGPz+
/T6EVmAUVnnqCzzZyqJzPNtBKc/t04FGEIWNAx9KGgrWuvaPPLoePUNka28vlApXHxmWOCVNzCMb
PWUdd36CHVfFLdrnS8wN1ye8GW6iIL/70ctmsPKKxHa9IIDpP8sWdwrGH9QOJm1vAZACqD7h/3sk
YuyzCRevCMqLR1s8CPWYo6N1v2wADF0SDH3kS8QJ6fYc6/BZKgyyV6XkTKAZLWTJ1wWMDS0UECGg
7ibblRAZG0DFEE7WwTgjZCzGMAp8sCPfDdMp2nUDpsDrLxDEkPXqFGeWyCjRFjbnIbET2FudHmRy
AxqJ1BU+IY0ra++ielZX/4s/X7pbRM28UzuEhMrbNLfx9uob+nPBXMaVn49/M/dazd6anDxRWFlD
S5eIxDQjz3zIZ1fmQtNTSveWgTW5Dd3HoL3IAsYJpdKzC/t2f9fu9eIG6HRibslbt4vNIWEktU2Z
VXQjqXYGgKMCMFtJ2+3W1OAeSnkM/RChwSYKsANmOm2IBtvmrXfPkuobOmbtT3HJctbYOHr7cbor
As12R6Ct8eYTvjJCND2uZNn/MVWAjF6+cDF4GWCoWmryW4bfiD7zVZZIvqtIgyCJQnwaaIQApnnn
d8IgqWLNJ0qjPfY1jPSH1YzOjNeyP/f+wBb5vzmPOr1VyYJ9gHZnsPaHq6/+S1+8E5+JVOwpn3q2
Us2IOPBkh4CzyvuQsTBuanHaDyII/5B5T2P6Zk5cdCYgdLSjnEUCODTgAyN4ceQ/LRnTF4mBl31q
8K87gz930nRk746I0jmp2VKUKAkFVyq8/paaDiszXcRxlZ2FjSik1WKwrDEQH62mD6YMop7uvsIK
VWriQSavFCpZKOUqeztigTXnaC0mhFF5fyoLqxEIgwx4/G4SwIdLRoLEYZHp8v7eGXRlMZbLwG1b
VhNplCGW2B4F7Aj/P3WyUoJ+e+pmWI3dbb6pd9ulgYO3h/cvsbTLR7hNk+attWAX++zyVAU973+y
+4i/+nkCu024IfK4pDD7IL4ST9piqxISTyeMcXRv+o7jId52b+44EYK8xbBkydZdT2HMAesFweFQ
T9lUybNMTIUTtFTT3sXE4gKckg3nAtjNGzP/fvl+J7RTjZIBfZzvxQ0cfUXi2hqZGYoWJmdfzbQL
XWSskoZskJQEYS09rYaaM1l3KE+SZb4ZkrsCOzE9X3m97npNQGxBcPkTrCiT3SXzSt0uJirHc3ED
dR5U2hBZD5OXHLuoZNr+mTA6tZyoI2eSMsIp9NBlUoQOHkmtfcTxCiappEZsaTEDxt8R9K8J3SDa
DDm/e70C5QN9mMe48cUXQwU2glxdXwgEtkdQEtJFDwursn2echieqiYzHmMSzjF7UjImYhVO47CX
1SV7m/hSG05cHtR+gGqWpMKbFMcytmRHzfdJzli5yfvpJxilNa3c/ROLgZS7/TBjM7oVTCVurusB
SLETX7KTYR5lfjHi5wwcXToZbQqnB/X0xwgbAUVOpCuI0F8Rxbx/b29Bf5Xbai06wunKavB9E8O4
PxvA8J2rr//++KXFPLKJA6X+CxyRyw9F/emZAgPxXZ/g5q3w22kjJoyptc9Lygu9diFK+VO0sPqq
qXPZGuB5bwDDuRjgnq1TPNruUXNZMM1/z6x3gGDX4xR8RFeqs9CFhnE9Sesmu87F642t06a1pIkB
5gvlxwa41hLVw3MKibTU2GC+wkjQ6Aoeki/sWi2phHMEnkoNK/EcV8fWNhiPJ8rxaMnVLjs9knpr
FWO+dUvR8228CnG02QcZZFkfqRITOxqH7kTV56LrwHHjh+s0vquKn/FyOo7TfHcmpqRD7+J7yzBu
uGRNiQ9pwU6lygb7aLQIrzI1MMl9jY37IKOKiKYeZru/efLLhS+TGZw0aOuiDjwrwp5airUUUh6m
ddt2xlUKhYcVhBqsmwRwSTc9AkjvY/Spk8OIGgN0IdrafeSiU8MOSFVrpyhuzZKcQD8+DZZAuaUa
3fpcft3P/QmxBWSL9VnpiHA8c/f9biRhflD33XTsBOIiJQCj0wuNU4Wd/B6jMkm5GlzpsxPbHNUc
csJ6MuX8H+QnspKdOAdSexoEojODISLic2jf2OylI466h3vHgl5WSnm+ngOieXFbTHu01pbSwMle
uXB+rnibXixmpW7WfQqd0o5eNWnuR9ruANnmliGI1zHssCiLBGa1TdQew5fa0XvJLMB8sG/fTAqh
HkcBvQPAEPqQ1Hr8nOY8gc+N5CsiMwEE5o7l/JwqhuRbMgyVFt6O9H+kzpMtd6itIXDKQwZ8ylxd
N3rXLp5OOkfgN0C6YmPbkfBYWWjhsniL2Hif8S5XUgh8BfJdQItWfxHWCHhm+YyMpgeDqNInkFpV
GNyd0bmqMlh+tAE44DldtBhL6+kqcjfxkj0Rb5MWp8fXhi0Kgl5Tiz/gNV5pUobtLgQ4kqAPHrri
8tYTeXs1D5UUsMsK2shTLGWGiqoxAxAXKMlMoTsb1Bd+Z9v8F0LNZBjF8rp+tmNNgUTI9UzfW9HL
LnN4zbS6uHOmh2mxqJ63FvsMPfV45iVGD9rMkH/+59rIbY8JI9YtxWMRDSUVmaqGvOklzdPednGJ
Tha6Lq1wRk8B2P7npjyRCRhDFN31f9q3ghlIlcucZlFLcUiH8YSgYCdNPpEtK32YecdNeXGTKhS3
seih0HiPGrcDMvGKX54cAx/7NDxAfmWpW9Wh2sIffPIpN15dHiK3RhU4V0klAmE/YupSLraBTdF4
9bufpdeMzaYyLsswa8qgcrR4Jl34mVsODLl7TIV0KqrvYbYa3b1uP8hEfhyy8CswH/tqdj2ken+t
CeU9Gx3WqMS8YfJolSKmVGznGlAleIENjzrT1FsM9pPLEYomM+yx8R1l45i3XbBORlpqGaCu99WJ
b99yJIDGmN53PYquCE7KyNvtf/RD3oFp9+IaIFZUXCyQMLg+9/c4u8yd1dNpEwCC46avFFjGQooW
b7aRY9IflaegBvJ47einZAQvyM4+qaYKyr1yEplfGtjo31xvxR5OZFVIARvxOfnVRSYh7sfSThRt
EAVOPVRC9lymdZOOg0jLYv6jU+Hu55kZBtCT5+/i7eDhND6jh0EqihHriVVhQrx56yfMl+S/t3lm
x9UXIEvanIx3yxIffdzomkVFA0VAhCPMJeYMZ8Q5uWi4jikrHoRgcpFOib7pwgZ5x2Ie2lp94joi
GBgzw4chv2QW2zXC24uUigs6wywVvJqiJd8hsSKwz7ZmxsNagsSiA+B6NRJf94dS7uvOH8+j/u/a
49dnHX+tG5VLX7jYURHTmTjCAxVdXyEDoYTkR2wTD3ACRFNialOl8lBPCI1Yu9KCUEvPs5SAcz7p
EZRoRAYA5QqO+4+fzn/yeeCVTEWv5xcu/8hzxe6eCfkkDdXjnS6U7qkm5gtrfH8IxFk/ZB9CFHBd
aWk2x2ob7E7r8okY/EI8OKS0vnF5o3adLNxY7iZnbO1e8DfZyhc4HmYBfEey0ts3mUhpU4Gsv5dv
WBAe0J3KJBxwGSqO0JPIX8XBcv1TyrGDi6BGcm9+L6bwVPRiVY3yGmC36Rqls8Y7e2kd25U9RcDz
WHa6lyqwhYbl/dPyNdE5rWR8LFS3/EaikixNcAGFV4MONDopwMy/DbDjGnB++CEW/Zv9d8nGmepr
voJ1uAvtbfm93dG0P+RUCqpN2UENqu/R4I9cRrjxun/A6zvJ64fPyOf4LyOOzsefkIWi+ebbqiJ/
oDrPjLCoW50FVUvBqVxq5fm6FiYBZcCRVB/m/pdfjKg9FnCxiSsb6vScT1CU40I9pOpT/9SCR03k
q0rN8g1UVxX7sPesW9F44nBoxGh3V0Jb9WasfOD2i6OfdpGw9/hdB+jVI1xk2liX/UUU4N7LYbyG
ncJIU7g+46wKaZpdVk1oKYHNOMbg+U+VqCudWGqaf7ZwQgyYLXrMnct1exgT8WTSrwA3wKsoF6rI
1hZE05573kRisEz3T39R+8nc/LG2ycg9G9E+etRsw5KDgDCnUcumbYUrzhVDVK3I/GYlLFhSbKMY
2XNrek0ATG5gs+IXnKw5uynS/f+qZarN//FOsi9857l/siDnMqY7++BSEUIRqppO9t2tSLYTOzAs
JnSGqLDQ/Y2TI7OdxqMhWEYhhEW7eTcqJyTOUc5At+HzozxitZk1mllvwo56zdkjffgWY2n6PSa/
SusGztrMg7l4cm/4F/9dXgn3UPP1bc42Yh6vd3Lu3R1vMYRYcZrSAEYb3u06xi/rPO7Fx8i07tmh
X9dX6UtMS0NE0fv1Kg/anSYugdScIYBUaXCnjzASZrhlxsHpc0eqjngYSu0p97JuEZ5JRJoa9mgW
rU9EkMAk89aiuj3JGyDZwdmaiwlaLxwn4SlEsAnRK1i+RpXJy6DVFziJnm2wXaEHKT1E9abrv5nn
VHNvPADLbTCdqBSS9/T3S3I526rc2mJ75pVTkAsmI+lVEpOwVEqUUjmwohfu0xWvR36Wv9WYCXC4
VxYXuPL5fY1bkgApHuH7x8KdSfZCzgLaxbUEUa/nHb1BOy6cXtKwZ8h2oXGKBPH5fyvTpCfhxEr8
L/I7fMCb6zL1VkdElzJY2pbqczJ0lpN5wSHID5oUTglZYA2ymaKwlYEj9W1Au7I9e8aRiIQDs3qn
O5Y/BgkBW0K5eqXiPLZTfjeMIrsa4doXWsU6QDhCv6JL0J/aWy8JEx7krHn/f4DxR0Y1hifoNhxE
dY2q7X3Q6PnVY+zFgENHrYQc8u564PZxGgS/+SFUJacV+/APFGDeUDBV/gy0aaXcy3mKVLkAVMeV
LnItn5eeRMk3tP8VU2jDljNaglG5VUGSboyf25hvGVzXL2Htl6kMRnZqGljgxt/AE17JstiRoG+Y
vMQIKajSckcft+0CfLQ5aVmJWQYKS8iKvd5C6uQ/wYj4LhKPoLa9TjtvM4sgcx2OnI0xNPcVqw0n
SGuG0I4aQOYSW0q046JZ5ayvJEtcJYiXuLR3QElYEdK4oYaX/AVJiVO8O4Z+46BO+MAejqxzBf+y
ZGJzc0OJSmT1YKXdA+1YWqgN3KXPxD7H47sSZJlEOh9t9LyJRhiDmyv8jthrqSlqJTsZbSSXC3X7
oRN429umD2HHbCJZ1WVuvkCeiGBbRIyRUV7uhMRjypiBK1HqZ73/cWaIn0Fe8a0zwbF2nQdvsxxI
p1Fg3VCAsmcMJYnD1spvpnb3vKNsx76xmxxIfLallESW1XBRLcaNt8GWHRqW06zfsgP0DOxhHiwg
20UN0y+ZuEFInYYZ0yb5WE5Rmo/ua99t/QlIC1Oe91sTTHK4Cj8BZoXkz/XLNQc+uuywJuAeUExG
AU2rPp9EptZ3tVtSBXGliSJCJrdkGL/ErdoRcbQpAR+T/jPw/nH/guNwQkw7SercHAFRY2bmVVQq
5FxE6TOyOI+7vWu9YZEK65iW1nWRT483+T/hEDrLxOcp9X+N2iNkSwKw5unOSaoNJjZ7EHO1CM39
aIE36Wk+fAlI23GCG7xxFvU4HxnFOLaIokypTt56t1NH76OYoijB+mJznnfEXdzFUDoHAyg8xk0M
EF/Tf6gQxuG2ZMUaAfAFDCvUvSQ5VJjd6KsV+nFFS7M1/j2JyedU11XomBvUEEYGKlYNRDgjWUKG
3UutUzJjnkhMxCSZH+wy8UaE+D25JC16Z5Lt4Q1jucTjYCS5mt0lKMY05BkgTy/fXqhEn7RjB9b9
uyASHYU21bHCELdLn3a3xGBg0SHX9Gnhc7qYyQq7GrKoGj5sYmzZiVm+jNY1kjsIssFoHgtBwW5H
tlT//Pwlf3EIJqZex/MGSSH1tIuCFP8sKz2dfZy4CuFpfOxzxW+AUyk76EcJtWUFGZHlCvMdt9co
eJdtnmSKhDP70rEF0ZYBYSFV5uxnJYBUbwjGLNsAEWcaJAlgJylvDQPRyv+JNLzgO5EzoFwzjKYr
DbVhnKmwh4EOAKefgsgCYUfDOPwNaJwPk6Xvct2q5FjugEVheQ5z1BTlmajBLGA6P2rcUhUE+Zf6
FUXwbexIADRPJ6HpVi8oZqL4FQwg0bgSvH/ENOLckfLJ5fJdr4pBkF1SwmWCxchL7M9Tq2F+IAjc
/L/A1dhBNIS2k4PyBLfHd8mXLioS2TZB+MLTr2QcKc+/LcceKxBhvSGKOT/yD3f/7A1OBy4vstib
SF5ulchlQ4JxEC+wQnUEd1tijMNpZ0xcW0WAcvv8IEqRiePCrMBe4cxWLSB8pA0Km7xB5ypMdize
uWfX8PMlR66CyLJYPaALQxPJXhzEWOezMXrK6sGVNiDDKyZxNzuVU1WZVHYf/kCROO8JxyONQkZz
U4vw0qICnOI4blaR/+ZZEBcj43OwwoHd+qYeAyoSxUWBwvgw93+WE855GMdBrjVRU1n/S5wAyUa4
vaArGTYhjgQn90RksRRquTly9Hn5qVecBZdw0T91DB7aFhdbhvalVg2Rzw8p+IrUEO+jnrMROesb
iegfFv/2v43myhOy7tGr7k57R86HMiOHWsBhljiAXekxvCzSHAqPKYnw6feaTOOuNUDjzPzAkVQw
Ch78q1feDocqZEqfnHgbTu3fofM/vOEbZm7AQoAt2L2l0BYw9VukPJmYEFz9GldzZ53p+x+oRPH/
NYJzncbde4Fig0O3vj7BfNkiTBEBhCA3ShU7Lpi+majBARDc0CLe5EWH1crcLyu8vd0jEa3URIew
MZG87ZFtxPXEK1VcJbcnNUhovGGj0BNuO6P7+ZgF3Rgq9TgQO8/+NK8hxU99h2dxtP07MnKyZu7q
9Ud379AILZH4CGyhc3tJbwGKlMu6wOrTLoZFuCNoGZ2K0gJC76BpZna7HDtP1hiFFwt3brOjz35K
YrpwU0SrQ3IP2P9Ui9I43QDoV6IeVxZZaKOM54gLPclhnsVEi5L+ACS+9iY+y122m+VBa0qYJxMx
L0msU8utYIOfvzUTEh5Uu2c6zqKPX9x7ng6U/K0X7UjMKJHIDe6r/IRxVNE/LDyCoURGx606tqv6
0aeLodKDXU4V1k9+ahKtBWBVpgGChxbwX0uMKuE6Kuuy6v/c5ruE+sHSBs/RkAszEHB3LmgwE1AT
qvJEAxNCv005CIvp3oj4xYbCpX9CEeYCNgQSkVxamK6aBEIqn5qQTtTZbA+5RTJ6KVpktSowyrDt
tdjSwEtpChxcSIdIFP81/71J+h8SWv3GOAoekj6hCVbiTMK8v6FefX5OZzI5B2utKHqJyQewAig4
ARmU8FhzbOW1gEzU36juU0SrtnESyAXUnaYO/qldjjgq2YL9TGIxJb8CUdq4ElAn9+pPL87gIAd5
mZT9JPwO46v4T6TvqBtn4vHjMLqmlFMvFRea4wB41slkqbbotN4lpiRUb3PSJfIkuINqrI40wRMR
4JsM2jTSreQyLOAL1q8gIxrh6abh5Cm9ISA+nG8qba6yWQQUfU5gv/06aBd4/7Tzbv1YOlDef+FJ
eQfcyi3weEX/IGvYg64NJmE0rkwPKXmBQVCcH7LhOP2aoInntqUnAcXKYv41JQzjTOnpBIaHIn66
GpRTqeUZRCD0W8afEzUYX0ov2kMnoX2u8pc+9oF7pNcbGmCSPKRqhQwDGonhnilOBcv4OkYi6+Dw
Wl2p5XoVPqLcjOIyQ53nNGvlnG+oqX721KKPGOJ0mrtOqquasPdTE9mUrJIDrcsWOIytTVFG+XjE
5T2VmnOjUCbRFea3S7ouRmmetn6cSa22OGAxJthWRKiRBpO2KO0Kbj1aC3go+PnS4CVjEwg4AVFq
qF/B6CHNGv2Mkfscjr2NBYvKlVixyd3Pgaz5SsLTK4jvwd1XAxa09CPYefoayL5t6tmUWWIZ8q8X
I9i8KB0XjkNTyS0ibmvL6gSFLLy83H5zGTnuaFAsGhEroruKm8VDGOkBK68g3HeWpzZQ81TKM1Eq
y1Yt0AanMaTR/Je+LfYy2r+0VvTxLpZMMRLFkkmXwFTykKhXPWM2VmIcws5OFkUNYWz4PH3hGcog
qIxtqO9rsre8wM9h9mqSeQkNkw9BY3Y5sksla0srfBy3ZxF+0i3Vpg4+a6Hp1y1vZZ+yP2UF2Q4b
+tNzlKrfr36RvHBnnQzMlffk+iWr2SGEssA63o6U0YK56qWIR5qcSruBaRP+wlZ8zlCYbA2rwhVX
RWcqksGA8SOR0nzhzt+ztocwSAff+vkyxzeeqyhDyIg8RoJzDQCao/J5Y8zFmqK21CpzsACwLQxB
9ujYM8PvKjnYWFNh0J06Cyw/G8D1L2VWevJdUBBgOTN9gXUdZgQpqooCeltNf30fJaQiNsw5tfQu
9jKonD1VITGHUbFx1DnHpuhi1We/cORmTE///8a4kQ6UcVE0PvMFdwr+fcibcjg6myn/cirYmC7F
SsI0ufJVn5V+gvSayDrRrCJqGKocBczO69oq1PNYFQ6KEiKbQApSErprWpLoIHGGou/auHIcEqML
OycB1vQCx5IDgIsweepJQsSF5IEX29aoILjHlaNPdDUxIStgIbNQMehzMEpbILVa5t1G+2SW3Vkj
YdXSU+CzMExBRA54pRhEPrFTe0wI1yEX5Goz8u+I/Q0FtxNkCqgRxkDQttCWzO/cdtZ3v8jW5Vwb
gnyZpsR4EGnM7ysMS9UClMVCddFEc+ySIX6xMXN67YmWvnsSK+r2fttZCf6TxE168RQwEBJP/ihx
r4WvS2cXEVoE4H8Bs1EC0tXyMOdIEa+kOikfijqyJ+NdbyLYI3CgiLG/iJNM8vOhZfRagJkLCPyF
/VVwm7mq/Lu3LXkNEuOUhuTLM53JKROqf+0tN0+IqRpGpdXHCIG/3b6fVGS/BFgNfUfFO6uPrl8Q
2qiU5ovZRKKlXumgaWK6eMWF+ogIFTJMoT1di9MoAQXkLvRzoOT/tRco8m/1bwbyMz0ZOySgEfR2
CdMDlqhIMgJPCw8bTqN597uDEIxmR9uU76QCxJfefd+corMNtoM6m8D6X1scN4x2mkY5xXZ3ENZc
9Mf+jWTpQqvYfdVtCXn98PXBKmew4YguhTv7dIQ850Xc0jQSoH/LhntQS4pSek7EvCaYmFLHyBSK
pjyQyreYlbnG9V4jGQlKGLgzeknZRPGoBCg+4YkSOH7pSeNZ/TDqRfCVP45SUWPQfRCIG3gK+bem
OQv6OQ9e9+KYhVJ3SiOz+vBqLdeSgbU0aqN76wxZYKI/MpDTzU5fgjQnsVHytXo13p09RfiAgVrN
D56TAH9Gtq2uHdeL+EZY7Chk7AhHiuwKAkqah49t8Tg0ef1GeltVqlOErR4CRHCl2Ac3SN4zNE4v
/QsLVzKXPght8/DrJ8rXaKyIxvlr+0hMHR+CPbHp8BSJXNoquIZN8pb3QiYZIleEV0HaxhbQYO6X
72qVuIi7pMAXe92wBTYsWwALut+9Ui9IJRSIM0IzZ1PrY6ljLyhxM2L9JqxYpWVuxzbDcg5J/6+g
tGPib38tO6BmsUTmlKIUfbjVxpWvuanDYzCfUxKXtutvBGHqX/iQwrYtbR8FEvSXUWTesY8WzU/4
cukSobi/8byd/UtNAbeyZyO2RGcXXzZCeihMekehmWdCtJmgMLnmQoYLeUppzxkZTdf03dEDiY4E
BOxcHJa3VszL0dlVgal5oAy0QTD0Ys70bikUvBRX6brQNa5assGyB+eytBSjszBBJkUHsO5aHGtK
a6hSOd9+JhZmyIPUkkt93fdkSPg8k7y69XTFLgSxNcNNYDAAg7RtnHLEso69gvDuasCSUwSGrN6o
me0WgQ6pZSIsSzisoCjGUI6w6Hci7cSnHkRinnEeCNu4ubTsQn5wwl+iimawOrtRaT4vETDSAnLR
EgfU4M/4pD9BYTaL40y+uNGHxZ9aIPYbbOtduqR5LpadYgr3nhlh/stuSWX9Ngm/1z0W/jPzbwJN
3d+RmhjphvKY27Mq+R0fy6nbQuGIvr+e4t4/ONfRJFEs6g2GF+IOYmO2ghFVvafuss+hFyPdhouX
DJj4rR/Ok0vfd+wynQDatNBR5lZuAzZ6VXetCFmhiNMxDTHtBRLEMCvRiAP2NambCaqJlcMBcBNa
DVCso0xryhHqT/4gm6aRlu6PAI6Bo269OcI1PUa4+4Pe5yA1NLsGngOmJV+sLBI41Ma12rU8zut4
RoBi/+T8+0JJpRoS4ujCKVno7VBA8puPsdxHbFxUjvlh9LCBNgIfG0m96T6c8fQN2HZvHOPugc6h
5Kfig21Nc6EuoJJG8Rni8BplUM22psBOi0RRtcIIQsiFH23TJ6uqaTr5aWPQxbu6Qrz6Ldx0Q+1o
4Bt2iATWdhU3uJ67bGUus5qG9g5BON3x5Ron3pFtdPuLXTSIXG0n11FbRpYzFg47Rlk3zVuY7yEV
vjJTv86AnNf/Gue0qEGVljX5WygiQSayUPuyJN7uQ4mI38VH4LjMetVIw4M8nJcBz47qWQwl3nWg
M5I2kG98U2vJII0aYbXvcebBUC67NzaTEfF1AkVoqTn8stbHb0kJy7LTM3ZG4np8IZFOtYsU+kh7
8m87RiJeA2zrW27U1z4WQiCG70T8AC6WvWCrVM9V/r9jZob48Qnqg969zD+9Vc0tZ2n15IJX4kST
fILvx0xDezbxYsL2gZ16tmVF6q7DFxTakGrUwIw2T8mGEaWPi11BvoP0A5x3pEqbwcT4EUJYZ7Ex
cgVCp1R8/wRnuWyJ3p+sqUUivAQlh/mcg2MKeIw4f7XBFxeEtCKzGCbkmc1WL4P9r+SSTkzJhih6
diFXkTj3B2Do4TVBBX+E5p6cZ6djAgGnEc9f1t/kvFl1dI75uc/pNA8wH8PVR0cLnYFYkgwubVjy
YwxrN83FxjTm9ifMysoq+e8GoOw3RKM2uWLS5aZBoKm+Q1sFm5mWD6XxIK7E9N6tqTXdsFg6Hn9e
0O7u2GwX0jhetTfrVwRO67VXQ8jiUuQitPqlmARsYQV2A7AtEe0akDZ3OOqdfkshdLSzwEYove/q
E9BXQ8cczJfSmZYcyi6thjY8Gg7jgr3iEBcVEB3FczvlBViMvJ3EY8huKEdUfXh4uLEh4BeSc9Yw
Xip2g38ckbO6TEi9qT0jhtY3D+64F7x9d29zrbji3qibnVWLwNutaC2OPqIzs60sWjwrp499XBHE
qB9SuxAdRdRpOf3Cl7SNlRhjE2Hu4ixJQkx3XZSNSarnoWyC8b/qw0Ut++xnjBa0g9sY+RdVd/nz
c3cOZxKAZe9H/resgC3jsAWRH8vrGQ34KslSwYnRVjZ1FfXSSSh17j6YalYy6AQKbUgPJkY28a2u
IyyyksEEg4uRuULs42IbHF4dyJLxqgM3XSR5jya7cppUO2NsVbph1yWDp6+SKqgCIZKQQbW92mIn
DsUtocfyRgLcAfJtGHnUllAB/6I0OLA6QjHih4QJnpPqshoCpI3G+zfNBbDud+7SBEF4GkH01rha
1066U4r8oAo9/rIwvC7mvoTX4ppS0EYkKbmwxCWjigfzQPOWzLvrl7C2NVakU11UjDUN7kSENCXH
4xLCo7IeQ5EsMB+qLA7/tsm08dwpOLZsIC0wO0bjsH3GhLnleAT4tGUV9+pse0wMkOEeGLPlpplf
whOLUojzYmUOswLkVRbx53TtNOWg4cN1okxh7ouUKP04D8BOljwSkLyVVpIjUV5KLxHVfaKX+zgB
j6Z1WulYod5ZritcuNokOQAaccEZeiaBFQZ5P07Y4kXcL4KzaomEf3Zfkmen6jq2Zamv5iq+W21M
sAVX2Bym5ifgp+Bz2J5iaFIQMNRjfr48s+DqHBX5ltvaQL/XSKgbtIkPr/XVX+up/rrMBpDNqZd3
zuQ/Y7y83WZiJnTIAGF+NnIT1+XYHg95YZQD3mrgauwGlGagDsVWLLpk/UxVmHHctqApfjoyUMrL
lvmvbYgktrY33kcfTk9ZVRXcBOyENiwWRaFvXIgy1y+4IcIsaNCYGEGvOZRgw5v2etoNZv66ZdIk
gShwBE6/PEB3A0TE00ydj9oBGkNllwz//Gz3RAzXJs64j2xxdCDWOFGUa1zfo6OB4G/dw8rvM3Ps
cEbw/IZ9zm7z9rQjwgflGrf4ko3IM8iRHaMwFT1RS/uuFxOU8QOOIW09J8Fb7KlVrGquOEO6NKty
Ied3PUXt/YUtKxf0HoS+nd98sRBa/PvVAHXgfnFrBfvthVTdI/M9tROHbjchJXVZdC5rQAZn6iVx
uDz/ZvvpMfnjHMhDjVA/cJuP2tJsmJdCCXBOhqIjsMXN6+nrgfmPcOpVINeS9yrqx2sXvQxrblNx
shqpPoa/cstgc7l4luG+x5yXQfFqsXQxYADnzU6PPgdcb67rk/kR7RRoUCj9QlU1lUC+6Tt00isM
qY8JfiRXe8i0OBsOmsgK6QwZNO36XBuxo3GkyLdYb6kCFowqyXyzUxEVckR+1+IL0jB7rJuSwbGL
r1hdGqRC76ZnwMDVsXLrmOXQbVgrUZL7c+yrO2jJgOCSOFwsKxTcotmM+/16uQPNE6yyLqQbPCiV
OWKIfgIIoBBMsWcptK+UwHgCpfxq6bkBs2NVmWg10axYCBROi4nS/BBdCjFxyNyPokGytitZbg29
w2hqWDwfX4SO+YA0YcCTaw6W2r9pqBW0zQEUL9x4KtExgdrork4/m+m2zUw/JJ9y/tUGicAhmfer
l17xgEXYZI3tyyGrHQxR1XAb5IhdfRz/tNMW5NYCmCN1wMXPnMocG65RDhyYEZ7wYxBsDCF221kg
GEDzu2oH8W+WYqUYULTK37KEJ3XK+N6x4oJC4dHVnyBYaq2metyzDPo075N+v6XurQ2qh2J6q8VW
kCid3SaONS42uRzwELdn869lV7xwjuDMxinunhqekHf5oRT99uos4OctF7y6hMSVv/nZRrcWKJ5/
2h6mVhTws1AZKFqEHMPBt4pctzu8XfExlaL/K53/KlRnzyA3DSUzaX5mCW/SHYYYW1HaOx5ue4tC
HiUzNsE9fh8YZFYdr+cmvMDEdUGjIu/hb7UJcwB1sq8jcxwWIvn0Zr4d56fIig9nekegtB9Iy6O7
yN7aA4naBlOxLliJqGv2dd5CkLK0K8akjhAl/mGmCmZ0HPL+fmj/aWaMsRE2ur0Qca9QbLTr1B0B
mRI3ycAhjvQykQPFAgnbQNI24TQB1v8UuTEpJdRYEJNiz6bMQGoJhuZVZtcWYR/RbZe1aJLQJQU8
9rDOgmMvh8HGGnb0NAnNVJ67Mu/x867PMM3ZbCSWMU6HcFd3UzbW7Lskb6XuZWbktLEh62JKiLgY
2+J6hI2mZcQ023yf0X6llO64Pb6UhHFznq/L9bs+5XTbJh523JrCIxXaDuW9KK32GGEgppj3IUjG
TZbbkUggfbu6CQ0R1e3/3RcIqR//11q7gT57sbyGtIUNzzBYGg/FDVXNKbSukEhjHROtfFpPfyq+
m0vgtW72KR9nguNqRmfOiKmvyioA96FqAyvTiF4PEf+/VcoFTZQjt2VZriATGBePGemtLPjEEuz8
69vQqkwuL4Udhw/28K/EL5JCBbq8Vgq2Aogrs8OYgDmL3GmA5U8g6WrEQGhYfH9vOPJIkNoLrsMe
SJjD+WboGIVjfuHDm8cyywud9Rag20uQNRdpF/cyvBMsvS02EWgEWhzsUSEYrf1xws1XOZZZVMfW
pl9BvDsK9crZksL0LAvZr7zYECmCbf852GpDhTa8G/YWGXVhJ2iClNMtAGBj2gBcTA6ivfA5SHbD
CDFW7Ne2cSKeWs9mgax3JBrnwvMqU+1FSS+SmTELY7XcZmvX5h0uOkIDOaCo5R6f/p37KCxyhqPU
8gOLdcIW5onb1NmuAbhJGEFPBJvh1gfZgwA3ir4f8R94Nz9VF5bHNL3jGkIqrUo+xbdbKQAd/RTh
mEf6E3betvEhYXhYRpDYpXefJeNxEIwd2aPJunn+VXobaWLzA2nSCW4q3cfy8EkzBaKFvZZY26ww
Usv44naTUCRiyDimwmS8uMbFXknRMv6XpJpsqF7qH+lb61BgUOtBXXaE17nw9rzGUr4eFoZ3OOc6
25jVM+X3iF+KRsDe8IEj380X2Lsg0PXJL7ZA+QRv/aJlYy1zcEQ8FoN78BCUXSVU1NcdGDgb2FWF
1A/IYhajO7p7DZvgueRjq+GP7yvwvi1A7XUg27xjPh/ug/FZR/MUYPKuPXEIfLbJl//TVuEFs6lB
HYhMPsLjmh1x2dHtWw00KQbNwCoK98YO+lneUdS2wDJgimpqK3m2rKigKQIYGqnFSeucwV6b+ggr
XbulQwZ38KpE7pNN8kjXEajOJBfWK29yb/3zMZUw5FtV+HQb8u0ZYkNOmZ6JsCauGkE3sdHJa/fK
fev4bPJBnz0ro+UZyZJmMU4r/LVY7NViH3vYqbpXuTMY4DRvCxm6BgvSXRIMTcNpNgho2f/8L9BN
BTGsI4o4GWYqB8IGlbbHufRWt69WOG6DSUXoAjr592UPzyBca4uv5np8/VUhdOJThNPgX4xPOf2M
cDcxFpF0g837MfgvnvspmDYR3fCQqyBz5hviP6BHHfG1tftU7uxg2nvq0DA+j6B7mobFry6l1qMi
go5BiNxJX3Wq7WomeT9u4eRM4HfynbEMdVzcmjPeJFdGTGMfzpjfKMlZsr+0VxboA3Qjyk3NfvCG
FVoAI8pjL8mx/hy1PVQC0w6qZG/4EMtFqE1jZn7RONg5RHLJdE0EsI61AmTrbhGvyksNSJRK5DFR
Px54VYg7ByfB3zGR1Qtq5FhztJzDLlmCagPY6GfTfuV5661DIFpzAf/POrhT3XHbUWEs61vMzFIA
7omc8avOch+R5xd3pPzyfphR7plrLEZrjNhdUK3wSYCt9IpGFmluuZt6lji1+AK7iQvCUko59XHL
sqpOH21o5RwtZrxh/FLWGC2L8jmj67VwnySBH33vSBvx7ieFzeUeQ5PVfvs65QklgmJr4kz6KYbo
/FzH3jSCZTtZ48hHOrukhisbzQ4d/3XUetT7XFg+Wp99mt89akyHZ95NnKjP2NwcIxTFjaeua2wi
BcMH0F5c4JAkDDqWbdxN4FkU5Pxx01H30JH1+cFKhxgZto3AX+DVTg1DXdZMoMEt86VDuYGCT/TJ
n2wLm61LdqmH5M7ktxrEz5LM9r+Wr+DCR7+IW1kXoWgkOVNjzYj1k8sSVqYvyu+SYrgXif+Eia1t
Oaz0xURnXmhzZb3S1vRkv81jKmra78iARb/QDcWL3iDBtuSEtuDeGWnNkdP02MEv+oVcKwi27LNn
w/SZcPBFnx67YSZpC4oDI4fb5v4bFsq7TVshPdbc7ApmNP6AOUy9ztqnhFhYh/Irw7XfsPvymNPx
zaBVeSLA6HOp7byu6U0+1FazVlurYvCXw0bCiTalHJiSNWXVus9a7XGkGzuzSKRjZ7xBx8rYwBOt
SGrdMUz6O1WlMwOraNUaKGzahSDlrxq1N17klrbVmNksYuGiQy647UyvA2TaUu8tc3rZwZcPZLdw
H1GfQAyBLw1vEIe4FvYxlhokNLSJbSBDbubUeP3tQ5jH1Hc58h/FN558CB9z6W9EWDSq+ePXnlXE
oQ7vIQqKF8z0UYMEHg9yF6XzksVQhhf1aLu2OajjoR/IGRJvtbfj4q/nIMqmskJ/Nt5qhjBZ+DZB
nmqdRK2SFRGJ/x0sfIDs+gMsh1TbuAlA9SKMrcBvvCBFwOFsm1l5WW7VkpSukJEWFDzp/C8D4AGU
dRUUmB/+h4Ydoxn+KMsjWw7DvuF6/M2s/27DPnJXlpaimnAIg99WlNNjek8e6mCY9ZN1QjHlxBVh
wKM+1sD31kXN4coPurk8k7IRUd7ZBKSvpSUd+5P8ZQOfGhao3FzJTgRG6CyH1DRFyd3T1j1N3Ger
p9TFQK/ewuVdgBpmouS4wzgv9Pj1l4NCIt04kTmMWecp5ELPvq+Y6WgqxiICHlCxI/Mjyx93ZXtr
QqQgq+kJfdFWFh8Fv4yfmy66MoEahqg+rR+eQlbIAUuVdmDejWCXjUYFKqgb3r/5qew67pL4ufLC
VUXPZ6M5WPZQifiAzdxYNmNdUlmI5L8MjSUYWKmHDK7tl+gkbXpQ5xODuigLnqvEo9qEdcdIoG/0
zAvxwJIQvB4K0dVxhd0Dr+iPDg/IIXFoa+NHC3vajAfwMqtYi96xGWloVaurOTIktkOv7ig5PY8n
Bdyl2OzJ/NpyQR14aXXQNp2QeZlbyCE1gUUQyR9K9pQoK2X1LISqO31ua2DpMdNSA0dJVI8m8raw
5fPF0m5Y6hgH+zvr/mjKHqvSmZMnSiZKshkZ0LdpQ6YVezqUZJXQBQ9EU/if6qlMKrYdiuCQ380p
18HkUrx/JF7+wdta7DkP829GAmMKKipiHxi0XGZiEGwn1P7IC56iYhd/7fj4LHlt8BSPnmlb9XoA
nSCUN6hN7k9Gs0jNECuxXEJk7fmS3Dwo4Z9BrBag7IwQt3E4CCz5iTEY/xtu5nE3wkYvhVAUf1fJ
HK5N8WMYHd60MYqKD+r5hlpxgM2maqBnRHW86Asu7bIuEdYkCQmcb75iDZAeAtqNvN1WN2lTvrIH
R6CLlHXxQShJxcWhF7MmXD0C2lR2GgWPxQ3rROzLWASZKgWhVYwRCNyMDxgRrrABQUYdx9zWF5IS
RO/QHRtAJneK8Vafdb+PtvoVQZLebJIFmre6t6sZRoXEzJjSowoKSWdjL3vV8wAEhhPmK9Vna+D0
0IxMDM6GL+IaA7mi8RCbRHgIr8SbZUjcrtRQdhtDM/0pfa1dNhzfQJWZ/ALhKk/elCn8WBl/rrM1
bA3FOeQ9Xt2EKZTf9MSIRZ6+9kPgstuFF2odKvyuPK5tMbD0raOmhzkD6/3i229D5Odr1zYaopfU
lXQ6IjzvHXl4TP+gEtZdbXR1FXuBHZmwo6h9KbPUCopc/uloOjMEMfwd9QFqC+sHTQuo1hySs2Kv
b4p8el/bUWbICgjOo4KXA18bjmYFtRHGzmUYtPM0yWU1GoJOPhlFHYeDL2R2rfOROTml9HKv55iA
2d6qDXAbG+R3W3AvpNL0Hzfnv+haXmxIlGDxqaYsGkAif67eIeSTgLc4qJFJC7XYXXxi8hQm7i4T
qPP5q4BTpUnZ+8uzbuOMX72RVHmM4OjaBaLRxJrRQ8tCDxb+kXiD1HO8+4bJkipvrDyQ8F7eypXr
A5NiL4EVhmCakgdRhRlD/krbJZFRSnZLL7X7qergyNQxYduCgInnG++iibaUWsdg/shBt6bsM/6y
HzCIxMLcOXDIKdOC8vXMCKHJ+7rCA7qJ91JH87K80JYO/uo2IBaEuOIjw62V3gRtzIyrb1pOV96k
3a3iMR6Xii5KY7uGpyoDj8naXgNVaW/bRjqQPxytQz3QiKF8jkg5wnzSaMpnqQ2EGs3mrlpLrH8r
WkGYAPaLahf1jbXqw0uBpmLK/+O9FO714yOWu2QEhGB3iQVk2GM//AzMFE/Ntcj0WvSlsxIhM5f/
gz34Ce9MVu8kHkxRO3A3x3LBF5Bqu0EE6fwUHy8sRK2YnHD7vMJ2FHbs0LKQn3zlcw+QFcTJMjFi
FiHlLFzxssNlD/HqgJJ7VQOw9q1QmxY4PBNKeO9/kQpTJfdCcIfy0PErjNMc+iTpLBPP8/kwM+f7
6ce3Lvi80fAZCOv2F8f8Ph4WB+8VKuNFlzxRReU7JAh95mknwQWO++FLrYi+0dlk5xLiiQMwECx0
dKBJXqgrifSxD52Stq49Zk5ctK6YlcZbZ1KObkMRLxok+BAGPtod0/Zv1RQ613Obo3iN806fWcRh
5667v1PW59CJaI8m7++3LRcbSWOBzSOVsQsqcqPt2Qje8gP0U4l/ed/SX+5OpPMdvRqz/fhVgrdz
g4oYf1OE7KNlVnl3F2l6pEMj7Ro1RFU5KRHS3+xNBStuC6NoHabZqYiOfI9azGjxpCBnqBheslEd
S14kEXRR93QlDGZEwTWDBsVquWHCUwa/yctpT+V8j3R0UH+sivHeH6R+ISE1aA5BkuloNbPIyfSL
JcYBW5qTeQfUjRHkrzWMN9rBHluSPGvNNREYh6NdqNlAeCfGSnJd0yVosMhhHzNL5QJNrqAJoSyp
nlpOMYmvbgualEA8DSFimBamvBe7DOVyjAOZcWkozj29kVB10K71tOBEml6ZgQSg12SJqveAqqf/
bklRq1Wr+IvJUoFMlKHyufb9Mn0JWzJ5A4T32lG8jZ+KCCnfpkAyB9DM7M77nsxF0sd9HEAPOPPo
azmCV5SYN0+Dc3yyPqa+IvWMtbffTfpTQluTjpUIvmOQf7W7FqibDW4eLMsa3WDAUtti7us6PNbo
4qQeEtvbMj8soQfMPlRaepGgB5snrUoZzsVaCnml18WwxIRUwcL3E76olwwghW3IMWHsgDgqhOOF
XRKPS9eRjFX/8gJOwBJiYzdggnmS1rEEva/4xiyyMVoDd+MOMgYm4Yqb+4yY6wnXqRJrsJwmyUIJ
ZDuDwML2UbAZHFgAkvRsVllJgerudeWZQ75lbF3BigLjSYaDvDKl5WCHLkcYAF+p/G+4auQ72LDQ
fbX4e5Eif22IKjoPHjjm9rO2GNL4yqRxfZGHkYS69FgwN8O/de00Gdo80I6zK81IKbpY6tjTEWef
ixgdCGIZJ/CB0xLq/KSFwzWzJKEy9JNKLGXri4NlSMEl7NHIhXExEazA94HNhGNKtFZYKjhbYpPV
NfCPdAfh5PlcC2P2VNL4woEcLOTCvRR5/AjhrZ752PQvIum5EdKWYWwR+cd2+oFZSA9eIW/6vAq0
JzOAJPE5jt8tSGGGp0U/0IJqyN6nOTbtnKTynNtg8Vb+G8On3f4GQFhFUvbLX5I161O+KoXhm3qD
NCZFTflnyRZTRC15mWJT7c9xappiq6T0OvfuXpXT7ieARVo1Va7TwP+NLEtAdvGCwxJ7mCQjtNW7
NYJOkiDYSmw4HkTqZGwhHI0y7VoZnRyfXSvDqO3+/lYz6xHL1e7SfGpFQvCH+cSt2Da3bi68RPwM
GTT/qQpv9eHVpfU/ZwZBrnPS9WzhJqMUYmIgrspLMiBBZdTxCzt/3PGhnaC22BUNw1NCpp5I3wXY
I0CcAVM+7TeWb4JOxabpDLBxE0Pvevu5R2FELGcRyjT/3F1fwYEXueQoAPAMBaEhE266HPy6eYMs
h7jAgvsbztijim59wmOqnPgU30059vHac3kbIy0K4oSE1PJHlAhocvgCY2iBbmxiryenD+ZSEPZl
RubfIC/gMWldJldQnMEl6moA2SPdAjUCOjNwGh8sm2SJ0LILEVojVcnlHtbTBcBFnTuNJCxL73DH
Pr/dl7DEohKV9tibnRAoOBUg6fn4qMu++VpK5Virf1D5Q4JOkvWgVIcBcq5SLuqZuWwSWS1WpzHr
6xKvms31n3M3kmFpgW73TtuE0v1xMWrIUH6eT1jY3Qr6xytsWY7n5fSN7OEej9atxAuuEJP7XGHU
7cQIrsXkYTuYlgMJUZ578+GtjIuN3gmFeWsVFVwXVbKxef0X4rmaaJvnFcse2GDmETPw8Ged5iU/
iOJIqIYQG8RDy4ZSOJ3x7tIiFxbtb3QiS4NSljGCAGzLXgIa4409LRlCJNXfzu34/MJKJdH4eLJI
+jXqvZAmU5tepS6sB241S7PE9pQE1ZaZAxIHKa7lS/t8BopEVvNU/WZ+DcWJM3biR2eFXuIcdL9I
aakZm0IH2xqYsgfOJdaTgL0A7AhgWVs2E9nYbHhKXBQDD+XnwHEAwjJnUoWtAZx5SZiO5lkQLYp3
2PRXU1PeoeK25K0kvuZKeYSdaOPHl8gyLHk8kekTsGdoBEBp2ksP51QbSAm1R5NbjZPq3mF9Z4ls
8DpXawlfUHWqeyutOfoOj+wNfq8g/W+QSHIudvVEVbQfCHV85cI0WgVJsPBM4nPtYhO6g8X8Ajn4
7Khsw89d06xPaJvjsTWLq9wyjFqta1pskNmEbNSlxwkJ7NJGHg38m5J5yfFLlhQ5/eUEWTt1PmnG
NQZwT33BwcDlnpOLesebiowOxTSrImMOWphoulUQOt1AuRR1MHD20jk5YsVUoaAPNWUWbvHx3zLk
EjB/OlYrdX9Nz9nCj/SOCjjplnMrt8FYg5rgXJTNXlKGURbzocVEociW0mXwqaNBBfkqp9zpYjv2
ag2k8J8u0tpxCJxwLuOYQS+LvOTcBcfMA6fgDWJ9V+ivcAZmcFaaXGK+e+FCg0eh8J7Y1pgEspQF
I16IlHabNeDxsGsUdM9mFZYYqeNaKSvWO6BUiMfiD2znmNMCsLwhAhS0HLMjOYmIJzEN0hMFfc/q
PKToF78SRVMFStxGsP2osaukm7rX+TFzbFkV9r7Z3W+OC0erox5We/0DLYdFE5QiK4oS6gs+zHvV
G/6moBOzF7Rj5P6bnriEkByY7M1kDMrQrpRthqt5UoNXosmymyuuojizDaaT+Y/q2yZMxMumBkuL
lU8QMs07pD4G6ZBuJiwbBPSEs8NTxD8IV8+GpjZiIN7II/uT5iz2xe+stINH+e8Q9myXgc5LtSHL
hsARXCI7hySJ2yp4c7IzzuE1yhCgo/ebSPUvw8UQyMKOwpDgLt6gFLBBtJKjbr68Uymszynk6IGI
IgbMUkrwyKV/5Pfg9g2YZkaq+0QailKCvJAaaLktnglba8VhBOe/z4k37DUUvyNigv6tVdrBffdn
bl8RmCphvr8xL7+yahb3HB/d/TtNIJLLlnbFARItGogQpoumh498/25ed2pHroglj+j1XGz3mgIJ
kSx2K8ucD01UEge5rq0f4PZ/Wyqi7UQxH0sTkfkJzpRdzdGVqatBdVHCbAW1Dk4UZtE4WA7hc2r5
KBrUpAUZ8SlNv/ibngPF3wu4IJ2/n4OHyUZ5l6ytFHVsA2kRqRaYICl1b5IGsCLVs3uWRkbvW+iZ
4BfjCmxmxwdTMu1MC1fNW7TuAYRW5nqqWG62Kiz/U0x2mdcmmcOT+eQba5bzhVc729i4StK44awY
6RQayTAE4303eRMEOJxheOegdalAgUMMLDsSgUh2miuWR6m9/g9wpx09AQVEe2KXxtschqLUAv/W
oAxlEpL9ONCKJE7nVhvPF/Eyxy1ReyRGnEjEYuSn56tx8hkqks3k/C3WFR3OCx9q94QFLc0lW7cx
gKocc/2CSPGVmkD73FSWJbDSiQs7LBwU708HhmIzzf4o3/C/VbcA+8IImwSp2bEbvzyHTM15b3oG
3iCNVH8jkKf7V+FOMy5o7vJQ3h8kS6IsmgoNuTHyW+zthVNkKJGdH0mbABwwXEiV6Rk7VL6gxfPY
bvxOVfcU+lCH040DD1yc+snUYyApt6j6WeFWA5I5O9a4lbXK1ACXU6TaR7LhJRQVrN3oV8Vz8yTD
6ZQ7upBWrSU22M1Hm25n7KwWhfDYtBgZNnHNWq/R29j7kfTCF44sxo83dOJnwfye1sP9+L4z8SxG
ISsZDGMYARUWTfGtb4x/BXTxK5+NgWed+hH2XOUQtA/rxG30MAszQozGUSSdhZTLHa+B0iM+7a2s
zf+d5IYgEI6IqJNPPiRtJkGR0KL5mYZZgA3NZzCre+Tvvz0dvmZBbrPbaDZJ2R7HeFj6v2YPNk24
9c5Ub1ffvC+PZ2EdlQfaxShaa+MuxYoEeBQM/6P76F6B3xA3b4mdB7rV47KcytkgIZX9nhP9Z6kU
uHXoNpMPHSnOQr2NBOww3VJkPc6MWNVsgIGOXyivpCIzHkIJ+xTn2mN2t2o67XLqi+snh9S+FX5f
ZFZvfnQc3wCYlK0hb6TYPmgcK0cQwvNiAIEOhNc4tr+tV+CxtG7yfiJJnB8fG7Yx8nFRHqsQ44K4
/EDva6TBpgOE5VsVFQl75p1eMb0Sg3hmavCJb7UZfX2ztzK6nQ+HUhn8H+hf3sNTYQkBCbh9XN9q
OgVe+bZdk0PaGjr2ju8SvbSu7GvM/XelbUjMECSlrV56jY2sqeE/r5PkkXxWImuR04gFOuu8YBPj
GLL4ag2z8sEjATDTpfRD8MVLyZHdz1+oPon163B4T+DwxhjhXpyNsbSexJAQrlZ6NWncBGzoomjV
34kALz6hSWqkUAoGAk7ZVL/IqpfKnK6bXItXNxINiv50t6wJetuf0PoDtLNrp7PwE6PvUtiNxsjH
u6lb3mUSqPv1nsmfB9HTpDBWwfo36/LTnN2OEhhWsk2mrJnfg4kzz/pmw4l/pwk/8j4PJsSZBNrr
9NNPe5grO0sHrt7SK3GjovhYBC4nMnSAmgB7a6kW+AMucyDI/bHE2gCqm+0HkMivXiu8Vucz8VUw
PwIuJ/ewvOh0S2Dxrozf14j5HYDCM0Xfx6yL8D54eLM+XIfKLUWSPDRVCDlgsaGriZDkHW3yIGzI
NmccHP/rmj6tFdg236BhWIWp3WkBxtzirNYipFZVSlXtO8zre/vd+ZGRBdCqyZDUcxkH9QspNLAv
XFbCKWb+KiZcqNjZyklr3fzYnGyfXhz0J6nTMZ5xRs0JuSXxxTRTy66RW4tewoYuQbLXzAHMBoCp
LwrpQHfUSzERPa8v7X1nBmxGZvrn+PXDkMjT9Yq5RZWQ9zN3SIYJjKLIcuSlCfP/53uMvMZSRX0Y
wcdgLE4H5UxqiuCcEzEO9FTVpoHS47q86ScuV9LXFLSlEWas5gMOGpFbbi+00KroT6nplAV6F73T
OYHE6JUswzojqNOCKLw8oq/YA1PYBNM82LDdTRXL4COBIh5Jv1JoP3FFK17vhZfoqcKOqQUJcmEW
cFUsndvBUeSjwxaCfnZDnhbDMNIv1GQdGiGsu1SqHkD9Od3fJuYkf2/5GHJmCVoKgMxxUP2cw0Ch
V71n23bGTvgsUA6ypYamyXHtI5FtJi5yfZoBDIbxoR6+IPtpI4IlFVCDf1UTqmSMrH7zhpLDcuhL
uyTtAeAmKus2f//CAXTxOF+gAPOWLCu12cdm1o30DIVo++Q1WBP/dZLfHPE/tlIHn2yb/ndYS5uE
OoJssoHEcT8ossh9yMEwufKrgnYkc2Ogwl+gNoQ2OL9bIZ51fu68Lp2q9DBvI/OsajjszRcSf+ZA
b21HWhT/XIMo4KTC2jlOMxqZMfQP+ZacxJiuPDe0Dq7MVxnpxO8bibqu6swH9jxIthie4Avo2ijI
IWXvioYswnTyieS1AItbMwaEXH/LzD7AKgtWRWsXozdjqf5+NJ0bNhnXq8Owp18pXmZ35sks7zZj
NDsV98eHEUjPzK/2oHjcQV1tnCQ1HK8WPraQicXzI2RxuFaPfsLuC88VvGtRDaOiHpexjDGMdPCs
ObHBV1NcGHGwbttxnuKgiNEE2QfTbHX6OQ7Dut1AozcjVvNTXuyC7l3wczbwnhsFuU7/oe7gtM4A
Tft0MOIEcPAZs8voxO7slmpiLzCY0TJcIUPLO2c7Fhea5+yveI4xxodry+5cTU5UWW/E/8pMinAQ
gWZ6LAvNdcEKZpJSVEhXXymEyb5/rH6N0bkRa3XXQy+fhI9z0Idpcvd5ljL1ZfHY2J6bD9DCz6s9
W4Y6jW+p/3IVSh3et8xk5vo4km3PAHUB2yQvYxIiNslk1u04KToU0sow9GqBu+O6pkAI1n2/7IkD
aBIsXKuKJsNMLZzte0J1eqIw83YeDfgH1I8h6g7k7KaWila72nTHLqakG8S1BkMG4JEfyrjJbMoY
oDOu65dyntIryDbn3OZeG4TWdaeL1FkELk0uXFGJAHYe/P8KX98BbHxUsAVqNSSGmsz+3Z1Pr11c
2II0UZvlyu8PofVlk4G1YExoJvcqZpi1rBpTIgYbnWaLwfHtPac1t+hCKTkSrjFioMZbnF3TkUTp
KdizAnD6qOvgWof3zb08MZ9pX2xGnp8t+GlDeTs+wk9VbwJ1v8374gAKJ6+hrO4DttCbLq/a0u9c
5pOR0ht/MjJEst4cV6WznqUWNN6f5bvoGmDHqHUfwENI1t04ExbX7lFqIDOc2/NNqTmk7MUKbWyU
e5bCowfOr3mtZppYr+3p/OLMsyS6Z10V90/rCNZPFmDl6vOrhN46sz8lHrvW3qca4ijHxlGvM39p
Xb8p+0XTNiEHMK6sFs2JuDehb/k5Vm6/+MEbnk2KF5EP1jjXAsjRXmFjiOfgJrPsenQb2WQH54eI
eE76ne859whR+AAq40ScAiHWVZ2u9b4yHUnEPYHz9kmk619azvjRsGu6f88dHrN792vi3J6ZLA+1
2/epwz3SmC/wTXJSf/eplzr+gavhR5HRS+p9j0tnyjbMATvjSzMwetHgUyTE5d2HOEdFbwhugHqS
5xSsc8KQwx+tHyXZLnLG/TfhhLZCeoiEBdyFE/l59Mn1FdPYhsGw2cx/hRuYoIskMvy1i75am0ay
DTGEYRVoQjCAA3Frp0tYZzKoy+pF4xFIycNi3Bp5Pyr7Z5a4NP2rKpWGXnqrrCCumI6RgFH1zIU9
V7K1iv1odeHsfqdZwOwVP49a5f1Hif9C2//07iGJdSvLETFPm8BvPOqO7eN0oVPC0zNfwTkEtAoh
fvAymXLT1YXdWjdqOZEQCnbnNBU9V7W/d7K6qkU0GDnC1LxzQDI3z7hIIUl5NErGnsbklmluhEuv
a1De6O1mcFqWNsep8dyzdVf5WcCKgNqpk4jxHzvS7xjao3IL4RfaBJDlJtCgqhfCy/JaQq6Md28Z
fGhrIv/quX7X4buAoeBacm+jULjuoTAk/ZianbNkLiyGaPLFCwPRHXfvZeJy4izr/h0cOalzTp7B
P51kZY2dktgSUHIBU+UH3yC6ZQCMVEZf6SEZMPEK1j3cef73eriW5X58wRJPXqyeAkc7mr9q49wP
9ODSiIQxINWwbZH9m30av2yfkb0V9fdwmxAE3K91uoiI3u/NJvVOuAbDfpIs8dKJEwMRydhlNqQK
7gPDjk+wHsZxD/SqugigX9cImD2VJQFwwRsdZqXOw8tm6Ymbl6JOJWcNgyyutCiobtx3qhVpNqbe
1sxZQfWgkx+WdV7gG9mgUyYgK+snQ7nYTnC3DV44l/xz+0Q9zVGnRt66NluJZNnMlT0kZT0Vpz25
lVz5GjIfOGaMHpvtdj7sZcTKx97t/27PX6zLZvwYYPw8GC85mxhHYmSCbArRqdB+/5+LSIG3pxFb
5/1MQ7YUoH8Fx2GsjqUKiMzvX/SimVqrLwWsQu6i6P5hLBCEj0f9Q4GSrPEALXfLhA23KB6JORpq
IYVY/mSTEAu7Z8CILyoKbaP2iyWGWlDTZB0VC428ldqFVuFQlylto4R1BSpXBKMuXFHrBjfimYNb
+McBHOcnMPe5Yyl30BnD6PTsgYcOlDHzceTdnFEV9jGvAkrfu3fGUa7UgaDbYzokjk1I/JH+AeM2
w439iAtSzftr7l0esPvU05mov1+XhbaJ/ry1e4FIdkRrxIJxKOlxb626bPxc3qi6VBo6VjmFwV/f
U4tcxzomzrkf7UUVbcP7g+F5GlY/Jipydy2RqYkDXLnHIwRLI+aQypvkNlOdA1spWDVvJ8LxrjOm
yu3TTIjqyBWSiCI9vKTWLvr999k5YMDnLW9nEGyKzMwimjvDUNi1UmyED2dUq9optA1rPa8NNJhU
5dfOM2XLFU2+dGsR0pdGWsbrET5VDPbsGfEZGZHNk7fIGb/8DD77wIs0afLtM+D2vWiNdqnY3OSQ
XZ9JFRyLycm68wz579CpATPn2LhPILJLRO9sGTrg/Y+7bffcJQKdzvu5LJ0kZ/B/qGdlr0EJDEJV
pqxqgeKmwARm7VmzJ3BPTNgeMcGs9ZCSgGasp3nIPBmV4NalwZLqFkuZVQH1wbG1sjI0iC+7Negu
bpaRo13E+iP4mqhwGgEEQKgnqjvTvOiLk9yS9es7M6n2dbDjMR41bX1z6gXhzq+1LrbCEVb05Y0P
fa6rtoH8Z9pp66aJX6U8PqFDSkpg+fyCjQZPG6lfBAkhdVrphl9RNn/GT/fdFVjZjVbjjpUV6wV7
jWdUFkK0/d8K7/3hE8ggoQbZ/Hn235Wd3PgSrwdHmAYtiAXcGvMcC6j34rGWTTN2IVx7Zq/ss7yA
H+o44tI58jAujCBUdlPRcw8vK9nRzaYlDjltU23rNQfqYXG1Buo1qTBkWmnKXhjv/VtWTjplcTd4
qqICcil8vilOMekuvt1B43l5/KF0fr3ufrqNCR9MvdR4iZ3pyxd6HggwK+u4mMwZYpHUl0y1+JAQ
qebM8cCtrQc5DTujMdSpWd1DZTKG4W1/lmV4M+yQeP99pY4YO/gCIMjO4DSgKV2FHrSvRnq9NDDt
LN0uXw5ewAKsBmMThkBHZUKAbiUUGT5C2VrtWfTpV1gPX5fi6vMQvrokxaM2tBM0qLrr248Ow85/
4aI7feJBw+ezKLmyvzrU2wlcjahHPol0K817KRA2VJdL/1MgyfpNtbJBpOSNVrun0kwtsdD1H6Ed
0ClIk3ALxfAhw+3O8ooXMBo7R4G3tZ3MQmv5d1LkgNFsp8gVrAVRXA4jampU44P4boiq99mSdxAe
dSpU7cdolOBtFlzWnI8yGi0KgemfI0xB0mSqbsUxyoNNupBuPrKq8QtIi+1WYzraI0vryQ401Y4H
s3Q7NXNvjGi4f7ZFOnny6a/6WxpprvfLaCjYcm79JJqyDQaN7X44qkuuDThyERO63e9zlbSg+9Rq
HdSpIUOj8X7eKwMfPSvAy0KjMBOLhWKlgibh7WiOMJ6iQbdHLnKqRZC4z/yNLrJd3zYRmsycIhPE
bIHSINkuzOCSgb+LiXoPnM9Rup/KwubC2luxsvqk34QAey7vgDO5NCHDEPOp+07hWtvFj4Ji+vDx
DCmAlWA/b98pPCgNvMHyZh5usw797rCF2MXcPwt7WCOEPGQjsjSgKpouxLB1P14nmQ7xREqBndCH
e9mDX1jRDsx96IsUQM0m0YycnKBjfN/JfpCz8EIEPnLlq52tdQmG3wdTqf3t87rsk9PovvdA5HX2
k8kQRsYWe8KIYZ0ZkUDAry+nKVYadEoGo2qOOPhBrKhqb3RgZsWDtkqZ2LPcGDthdravEwNHDjsO
sjLvijvqA5vqkKyCUAHDBO9XDg8xr5OovPFI7rUFqocaT0p3muq0R9pPpCT0RVmpKxlJ9KQgjjKC
a5ASASnAQhoua3JPRjBrGPtThWFeBJcC2ZykuTpB+ih2OcH3o+2JAJb5NHxDF6LY161XF7lmBufP
X5cSjaDrmcO/AxKtibVBEhS4dfw7B+x97dI0nPuwI/x3dAKVqBF0I5OgNNf3kgXDaW5IL5B+4FXH
/8AN/gmAP7dYgZumjF++OzE9uFm4kEtnd2axG9udHqE/ihAype4fDTIfpc+k08kaE18/BvUA0T/f
Uzp4W2LgV2IXmFiWmbcMHdgTeGNcnI7BwzOJ1qTKgG53o+344MHeELuibRTRiaY4sqqhXglVyaol
2qha8S50NP9+ze9x3Qh6Ix9+FTwY3FG/lj//ECgzWgZTBQK+pskINn4qdkQ33Awjw8QdofXo1IAQ
pmoYjj0OJVBMXbWpypKVrDmR6YjMllq3tfT081FFtv0GDaP93k1m2ZpUA/+0Pd+0C5KKR5UqvcP/
Ycf50fqzdEl5N2lfdHsUIl8McSpB/XfUU37+pbP5ikV8wZE7PUD2giPfBC/tStIVUiEui/b2KPFm
m65S1p0L29+3kxxMhpCS6AZNmhH1EIngMwMNOL0p18CeDmiM0blkVRyWQnZZss+kJPz1BbqI3a0j
ZiCwmk1cekp37E82S2JoepXXyLAiDGjCLdS98ZgC/fl5q0nBArFfBAyeIDnh/QE502GndZCLN9EV
uLbK/eGldZh8F3EvsN8LHCGMbB3VR5hNVKNRbHjynnhy+nNPkVkkSpswMLhzQXMY/o906UcmxC1W
o5a3M7LEItdt6kEQflVtpucCeK9i+7Lr2azYrDl3DjpJMqlPOoae4Xaolfynx/anC1UBLcjEfRs5
DYzfDJE+R4F48KWHp8hUhBcqdrJH+O5veblJ2jkuf98TFWBZL1iO08FcqI2GNjPe2HevHJ6oZi/1
6Udb8n1MO6STqhHaP4kOX5ipVt83nr9yikKxv3CL7GiNINsipn46zeD7/FGagawGgIsFVUWB8wDn
wnyo+kypwBG3GT1lW2hZGs+eA55lo72FbYqdw5ovoxjzhq8oUN9TtQoPhJnPlB2EI2uS1GHyJLLZ
iL3zQyBopQWlb4dGNi7xGebO9xgMzEFsDgW7T44bpnoejHAqD1Huac9lzYWGHE2FipDFEZyDZOkD
e6rg1XoxwEO+A0vIpj2WIFfRnJ3ehAj7YmTpP7G5q04ajNchH4ZnZKPlydHBtz8k8nmHod7br/MJ
W5ZTHLAvoctx342toxFzOki+S63jV7r9q6gduR1Sg9QFVMolHOUYBg2AA05lM7pSsH1Aak7d2R4H
1u7i3mV9hKBk1VwycO3I+GMntzpqo1mNR5skO854MeEFqZpOxAItKhNiKyZX4Pkg5hYfm3d0cfE9
4BBVg4+jmHhrZpsBVq3vWtYb7yTHcBpSmytK7rwodOX2vT8KcSCOLa2lQVby1eUZNPri8N78ttIV
OYpOdjzPSPX4kNww2J+E/MmDuW789LAz1Q5Z249qCGU4TW/6wXT5NLaI9rWexDr6cmz8IY6w9X5T
H38PYPsr1hm6fAkPrzm+SW/gpUIyl99WEToKy8wXxBSh7aF0/aOcqNmDg6s/O0pyXyNZT9MWnUtt
azWjXg4Nx2E6yMfue3esSfqajlcmMj0cuwtAc8qx8yTY7161E0Lj6LZj9L6m2nx2hOXOOJ6qlyW5
Wu715jkvBBrjeujYKdxh0+ahdifcsq4O/orsc8h+/ZTTDx/gdF1Dr0C/hWqE+woIs4Wmm6Hym1PK
h0aVkukk1uRVvWiyxVqy9HZGVTs9yCB54B8vRs2SVBdA2ERCBVeqjYhm9WIDP6a9gAa2SUf8+JHb
eFTQdQdm+nbxLsgCxI+KICDTaeyPlRv76nopVXMOpT790UXg2LUQfVPtlx6pdGXcc+thzL4IbkiZ
kfaeZL8epJm9c1vJQFfaxsiumvlnPF5Wou+C2TaJqahIK9ChSosi/VZxqvUl8aBFmPtyFMVtVe4e
Pxd58tWjv1i3xy1oI2CApMjn7KNqzQ2UqfYENAd3F+SM1HLuCSuDdNPNHqF7m+cJhhmtgXhPBMNu
oEbCaQGbG+vmoB92rEWV/0Yql5vgRCT4622Qz47D00CetP6IXcWWbAMoEYcsBb3SpGJVccsN9APf
Xj0LEq5+9HCCDC4LtHVcDbFjVvTAyTIgfMKKh6XcxzmRKQPqyvPSL0Khw65rP1S0UQO9PsmVF7rS
oi+64Tlp2AJCVgGLxpkdHPVt8RU9Rfeo5G50hCFK0CrIY6CuHqb+ZJDHDGlevfqOzK4X78p9jfHP
EFs8E/WCeiP57USEv1aLDZ7gGMLXofqfUkNQfc55nfDwJsz/QTC0HqVroODAoMUWRT+ncO471sdy
xgdksO0HHA4qFw6I9rwLZSuxTLe+WCZ2lglPjlbvLnISoIzfL79GxKka+CLMRu3CH3vkHiQTxKX9
cIxm1zSR9jcRxenORcj80cAToIISWqTdbEOd3Xht0lJMm6x2VoxByr9DA6HzpzEb1ye/JES9Th/i
+mHTtHBHX0GivSVOiZJtS6eVk1KPI0oKtQHgRl0RCQNG1w9oqL9MHx+YSy1fjmvZ12rk8ProfUsR
8U8O3PBTwB2pdsnLnwGMaal+T4OfmltM0DS8MbX0Sw1OYPGv113A5oYYOeas/ABY49bHLt1b9lgp
RpUIYAH8pcyA/FDXu00xhwmrZKzippl7f+dNYQBseeAAaE6TNEIclddLl/mERU1kHFbhr6r9s2lj
7rlBGT6IzJ6mH+5R0eloTq0fU4x1YCO+DBzs8anrqTcgVJT+qaWIV3nUdMoSh4Ag7KFYQRSfVsZZ
goJLE+ETx3V4cNwHuOhHxaXjgnvslo40ajAO9jp8y89GB+MHkLCnkf/rg9H8qZDwK227jDUwJ/dJ
1TftFW6cO5EiT8O4YKYUh+Wn1JU/xJeA4CpkNTUNP/kewJBqr3EKK92KtlrOhunlfIlhVjc8Tbuo
drAsS8iicZCjL3tA9ycxgiu/OsSwD8z9dG0rwVsbfFhq6jL7doyTMOdkDlHeFGq+c3Uv5biAl77R
9it3lAk9sCu2SdCr30qZ1URWwYuy2bciy8m9UyZR8AAsEvbHUTUmvLPBMTYOgTMYQrEwnY6x9dfH
s1AmStvSzykcy6t1bSTMsp+zHuhtScfiyCK5O1p/Lk9ZSje8LuVIPpV6ez1QCxa+NpCzG17MuIuw
8+O8zi0So78ODIxWyddXm8tXJfdKvEF7DaqcBqCeUafk29jZf6KKv76jQVng+5Z4DF+IScD1XAO2
HLOwvvTI/eKB91cfwia3/5aRfd13IhbZ78xW54jt7ilNTs0T3hwvNVVC41i8AKwBWS/ovRnrXQXQ
hhmG0bo5ndgalJO3jdY5j+zO6OykwEbcpym5PiPrEb/WSZh1mClueFOIQ7zkz8eEV6B7BULkyFgD
qw2TVFq4FXcY3JjITVgNssUGJYuZ0V/tzF08S2EgByBJH5H9vAe0ngOh4L4GyLicr+SG0IVgd2rz
ar2J8kLURWHCDQ4YGmswbNU0mZfHqS7pz2o2H9sFDRZ5DwSlwDonkQm0tdIMzTWRMBu5PeWmEJNT
U3gC2Ou0H2DvlWZm25Yhl5BWBb2g7vXtOabwl+OFqyFTM+gSXPbdyCBR7iZfPbXEZbUeDHNI+Y+u
ukk83ZBK546wd/yATQgi/SePlmmkCogF2GqyPEFjIR5Qo+KCLss1jSBVQm/aqiZMTGS42RdyTghQ
nj+tX8F1z9DFSWdoPf7NO6BFZE0hG++tkLzZ+JAvj0EqpZhggoGdPrp8aWCU4VO7wBjP4OCwjsLR
11RITadJYxcmBcEo3/KfxzwEpSHWA/APed8w/kFQkVc3hprqIypcITv97ARzpJcu+VIyKbWxBcrI
QGOnwxWnrBxOvm/q3V7SXOCYvulhnWDBFeX2zfIldW5vvKurMSwHWomKcMkAd+Vz8f53qH5+ofTK
W81woWH3RU1XKxPzepABXTjBhSWM5kLkBuPm/B6TDRxwJsRb3DhbPkDMk8IgYbLVZVKwLkTW4LYm
2CixPR6A4WtG47I++1H9mSa5szAQgZ9zLhJ2zl0Kvgze3vbFI6wu3JBTHxFB8StAJU0qxsDwmio7
zdP7wXE0CUE8PehwtmlIVprxVGfTBE9wJYZV4F7i17+U4sTxzGhbE73fLn/OVawQQFc/7XieLMVu
zV0ShYlINda16ePnk0gGd970CXebML+IHU5R2LrJXW7rL006CWOsS0P4pHi/6BOHXAhr58SNF1Zp
9ij9TeB+V9gygr2xFp8gAGg6AUYhb3A7lEtPU7U9glkgcu7tSwuQA+V05hqky8p3E6mzN2YF18eM
iUNRKbg62yrLsLTC+SBIS3gpYnYCPCQWDeXuxYFx1FPX8+rd7V1MAtMItIHrNNtMiP66AjCivBr7
kmcOlkTwCtk0O4UF1/mAJ/+Jys8t6S0m/Old1x1G6mYbgdl9nFBwlESxEX3zzgD9ea+yGzXkk/KU
Z2pa3bKWduKUo0YK/PaMMGnZA8osM8mV6Om9+0EdfJf8FKW9nZCs9m6PnC9wZClQX8QjnCRK00eX
7iVsAjDuagHP7vBSSn6uxKa/URdLnMGnUNavfGoIGzfzfU0oUFpCYVOmTJuWXcIoCemWSwcASsPw
FrznIMnRfITaXbVpL5THUzYnP+JOqA0Heaia36AnXaNhIX0Xn4V2nC4B4rdzp2yU9W7x5Fr5ZUn6
vsRu0027meKR1Nd4VoHriT1cFzg0f53ypU+EZHKJWAdJl+ahaspliWvXlSxNNWovTog3HXSRJ6iQ
aHMNy2hBMvzbeI9sRFw/O/KY6YGYxrtuwAKCjAEg/T08e0dBWpFUe7k9FG/sJ/cCFxEolCBH4v3o
4uTU9sTiYdy8LM1Ywt4h+M1ivNf1xeigvj5NaVfsAIpgtZN4GosCvHE4pwtEcEoaXu3lMs2Ike5g
DYHlywtO/RDUiGZWWCPdrZt/2NAZffbFha8jQSYjZOEdPMuN6j+9ZeYEFqdHWQwoEY1O1KB/Hzlq
+WdUWE6Y33++cUKPPYjESTwtZHRmaYoKT/2meACBbgDDA15AABLMJp2TLJvU5ir8guo6bkuXg/rW
wdUsFs5vkIvFpZo6XSPAXhqYN/RgohcL91zp3FPUfT/Bmk6dKU9IMIoaGdlNCcysW5rW8F2REUZU
syhmD6G03ZfzEyWYOGRLkm/bZKLPeu5WcD/hFlYvhlWVoDygxMVpv9SAjl1p8ku2Mtr9+pQ7oXPH
f8KOpKXkSWTHs8Ut+SqVSIxW0CArdqnRRFi9KXrUWy/YdJiUMxfva0Vm2ERxNYMP8NljGVwJuPUK
huo7w/xIp4yU9KYm+LBQcQvSWH2SzDpHEmZE8PLuNdh3ZOrX55yFCKtGzTwNFkXRc8/jjGYUjkOZ
1B8TVlA7muRPOYyVgAgFCQuWYhG6HKhwnfkvbRw3iEDrWPBiIPDxjLTQl49FeNntyu96XFg+xJQv
ptQ8bv88WEQfdaSeuLlJZgSAndKM/RncEzcF7U6DJFw6jxLJoAy9/J82aUS24zuawVr7OKcB7ivI
tC8mddFX7/tU68UMEkEI8g2N7lp/caUXakRsb7JiBV1jZzrqygFrqTH/P65d+fc9fOMBf0o3+XzP
0OktjPW9Iwfm3eVcp9zp97Q0QB43VTithCopbYbhIOyXIPDtuywomGShvjjOghD3VS72Paauya+o
4/aBgPByk4xZHlqZzJROkRbYOCakyRjQYb8Wvewc7tNNoEKBGL7N8+484fnhocvUHc0EleXcdzRL
5PUMtmcM+xi3kC5EdkPiKmXrp6CClfkaLFu/sM1j2LG4++cbdXHcdejufyaKWRiCXMEurgyZ94dr
kGu4Ni1wjM2/xhUPQEibtfx5H2RdI9DkRk3J4Fiwa2s43xun4n2tZHiyewhXawUlat1qHxARiBFc
B6nGkrycCxwadVprxjn8Ekc3gY7AQLKkBL33Agx6ghSKwvthmtHrlIbCxNy7kfmYSvlSxpNZ5KW/
2EaWsEWXAdDvMjrPuP2tK1j1ukkOhjUxIwAjog9l48O46fBTXS4d7B5JKINPuQha4IK87dv0PfLH
NMPS3Pc5MLcNuEaAl6Qz35rnkWjSQ87gjEBzHqMikV6aOFOCKSubpnJXOwgLcri0KHkO10gcXqwo
I5ouIYyey8iFUNRxmYbu2U3c/NiKQ/XGJ4ax8ddbGUtaoUt2hLpKpl8PcA+rzb83MxByL5C8b+bM
8pBAWEZf0isf4kHJOGcu5qWWx9u9s9VTpy4TShCBIfhJ20I5j+ZGr4m6pJxMB5pQ5WCmVm05kjMf
5wmuVjMiTklfTGuxndNB3Jn+SSTVAT01iJoxTewWORP3odH67KXFBDLcC7xfBcMwPMHzLAFGK4NM
6kk8nimoY02w5YeyDBGiv3N+Uh06kbGLVTDkSRDRcXIPLl+trGvuu4ofi81LxN7wkKrq8Lj44QnG
KUgEVQXqiXOU+HsuUBxPPKnxogrmLXB3j7/4ShplTR3m6pFvJ/C3w8ntH1ZyHP4JXzp5jXB6uvnz
CyKu8vDIiMEpzS5gp2hPbHFRVUz4S7GYgkxLOwTYMPvvAoj95eGlyQpCDzqo+c9uEhZgR9a6lxID
XDLjgZvs6KBWKGD9LMcmWpApZxFbSEJBOMZPWoJOm9bxUFnewt7JHWQ2JSduscHJU4be95Se2m3D
1slzyPecWyrFWI/dm/yX1cW2ID2T/LxGwadODbZDKjXt+GBkFkV3IEy77g6eNvCrSdchqyBMVzC5
jamFdTPmpgRZK/l9l93EDgqdEsi1RymRbMerw+YkG1jLCbm/1eLpryV7GbCGkdwNhIqb7Gx/aJSy
GO7GHmXLX9TTsjNL8fqNmkH8CTVTQ1K3k/Xqq4SEFai2JH/twhdvj56tRNcbWhQyb03EultUzJyp
tAFFwudB5WaoHVPhSd+vNSAz6P5AkYJ4qVXwT9rzHeLCZY9qiubEfIS3sbV3zPqEdxFGQ++kcyUO
lxmqbBG/Og+Fo9V1F3Sn7S/06098mfY8TsjGEJBsmnv9H4MimojvSV+DaFqpeXr2Cqw9BZZ4UkXP
RQnxnHHWI7cboHuvUY72+mYMsd5sTM8OKqzwYhWob+AwcwHJ7pZcwjt2sAX3H/Z/epIp6GaXq/Sj
RQgwDXXilnTJLsNY+WB2+EjPqEi2akAL7wJlkPtl1h9ELqogkMH34GF6nx/0Pn/BbJOVrSOFa4ub
pojnyaKLShIC0LYVdsR8U+blSDvv2847jqazbNcKQFEMoKCXXpUjqwGEGgsCCDaufqLXe85Iv4Hn
nRGVaa3OnPpfyKqjCJw4gTcWqYkWJX/pQuQOfnd9cFmY02t9VRew4Qm7iLRPlqwIBcwaFB6115iB
0tHPYIE/BOY7I+ukhFptCbHNpH4yPSnaaVn568nR+hN6HHQ2arWhsWqdHr/vdd3spU29fr+ANRIQ
Wb4w/HKkcHjjVNXFAWdeinsc80FiFP3Jt/g55Of2ptlUau2cRXSfYt0iohnxmj3zOBDiB3XtJjpb
p5ONqwjgLOXx3iE4FzEwXLc2dlL1qH1yaPvZAT59PyHfvpjeYdUt0GUCycwd/h09Zh+U43cDe6pk
5/hYIg1VPnxDrKZ9SK7crfQ7Ww4VhIjYlcKRnLLRLtpWOT11K47A2EGlU2vEWN6B/ov6XjVdoYlD
ZOkh44xZ8r9VxjwNPjNElHthsv6Qtk4mZgSYt9BZqoUIYgqMRsgnfANqnMG4vXC1ho15RnERikf5
XpfH3kbWez6Ntu6eO1Y8opR3F+Aw2uEv20eM7Yfd2DjIlR2z/xOzJvabkPb3jzPBNHLknEE3S63W
KYKXeAv+ha1hV5hMsqBfOh6e/syRN+kqG0chIrhC4dZXRnSYqJ5KpW7e/nYYi8atwvB3JSW/GTsB
R7GtHPe7kkUjRicUpnd4My7o9tTBNXYmtNG7TzxdrkdUU3SRIbZZ+loWYURdp41Og6jW8pgrh44z
xO8kvi3FUXD6WZgR3XrFfgTwoTjV8ATrf0YZsjXYmj5dlTrclWMHD2HeP1tZ9IKY08KnLB/utIyv
KIKejsHENLyKvzWcNRsRymmIyAY7tOrD8zPa4XTad+bISOCkdWHVjJBh1iSDpZVl0fg9WTQlSwII
GXo6oswGaMEGBmZqPBn6/HbprqWZc4w+pAuF3i5XkkQKyMdycQaz+Swj4ypln6ncaVCeEsjGKiTI
K1WarOGSL6Ce6ZKAUHCyBqTUG+FshBAOzxbj6/X81eb66jMS3qFo8N98zIeHoEr5XxPVQmejwGrc
LQy5h26riidEsv2n+CBfwkEhnfrHq4ccYslj1APHSXkuDkSl7I/emRDAFoJ8WfU+0xoBqycVjR5W
G356JxqGqgVd5BRoEYa51Y16OsuYY6AW3VwkG7NK34fh1lVQwmWmbfLdyeaXkbxxK32Mdb/r5hxW
Y2Z8vJ3+9bFfHbioGTEZR4nZQXmxUgIYqX/i2iPZzjIZcv5HCuxQ1OaMaFzvEs0+pd8nVfGyTCZV
fpJ/DmAmkwDJAba+2KFJeaig2G0eS1mloEOeTO75AwcNbnZ466KN7wHSGT/ukyD7C7bd3iJc4xKC
LA2391UKu3iz4dHSlFdM5MWT+ljqBCECS7b70rS82lvFo1hNxgr0aikilv4qW8iiFmHpwFGjcV8p
RotvpkVsMcEVmHKoGDQoQ8KoTBlGqYaPHylpNi8nHooFK85b4481Osp0dRjLvS76IFKu5/plP/kJ
UcMCnZXms0+oN6I3Z3rsq3cISvpytERn89YxIDe9qf/30UfGK/yO1ZoKvxtKE4inVnkHQSFsUCT6
vC2KMog8RFngXUYljirv0+N21Akq0+nxZTg2O7dv30I39J+t3SF7oBzY6qbjR3NGx5a2kcuzT6Kk
8LZzetNuKozE8ii56MRrOJ2g/pIWQoHOSm/gdit+8X3ryTD1ZphNtc2oii3MWAkF81YQdYU+99lP
ltv3gy/l/cSTB0NoFbvoeWj1ng8u1hBsPj8SOiV2GgUnUut2roiXtFlJd3sp25Hl28wsLbDzlEku
RJQ0pDX2Gfjx8Cra85Xl7w3gIA+5ZOHtqoQd0Z2BjpODuC4StukXUOoXgimqQXIKdCZv2y5d2ek1
pC7KGKAhLiohstPYw+/vAshFMz1eXkHlu5KG0f30gDzYS8+V3PLJkXowd5HKMOF7/Xhqk5/PYVPW
EjhWXPQLqGdo8gWCS/z9Wt/1GFYSFo0BSQoO8xomlSbrty47SHqidcCEtthT5+CSxYohJUpzjnDx
C1UoOivofusBxdYS2+Eovxda/c9P1fIRplMml+7jZtui0Ntty0g6kM/JCOZ4t4ymGtjO2IC+S8GP
b5gGG/Igsj8C1cvFmUwqMG+VhmCSP5dtL5FQbdjyAEX8GBvhBkBLl1nKk/y4dy1hDcweUZRnjLH1
K7u7djvydjtYhyQiUB2/m6C5RVJZTVSKPCM0hd109NrsMtFoJ9r5LtfhD1vZqY/kj7TFq7miQoCk
g8zkXdXtgWGei21toZyJ0AOPf6ExvtAAHc+KP+aOBBLXRMkoEnVqxn/iSPjoi/27nJLpahURLeEz
WYRJSLfLzXxytBpBxGs0XugVfSFM2wfyW+4itkUPIpJ3PyQ6BYvSRNHpUmumlP4EagkPNYixM+Ho
lYmZ37LY0JcezIJTQAyYOvjGWf9uVsgk62XrZdnUOCoruXFzyaw8wTmjH0xzWzyN/zpRbO0KyOIu
6ZZQPVIH4ob5cSt/8pwgf61MAHPslOUl4c8Ch+eKtg+knNBq12v7eKRf3nC+tt6iI8o026fQEavt
kykgYAaipv48T/I+b8mdJkZcPm1Sd3nop3nzMk1XMhR/XnULz5NQ3CbYCrz9pFFyeMgyEMGhX6AV
bDne1cTEug8KJCGxaB8xIOyqiBkJPhp6mBGO0aUwemnaimtwgS26JIE2rnt1IZQ6K9ZvZnPzc2CO
JqGKB2SnaXCoQEEf4xzGInHKjGAYyMbGMKhxQLJpfBI75TdXY+RT7DcnGwrbL24f+sfR9EoAFiFj
PzS/CKv16WJourIV50lvVNfrihE1XE9u0rUkYSx+okf37/lKAISK7OyBzMfZ5fl1cifgvajh4H3L
ijPkn/YCCEM2GyvrBkfc3NLvAAP2CQ1xpdxCB72YeoqVZXJV8ZeWO14h0oWguEJz5g7J+TwkZAZ0
ks/XU8LS+jvv5Uye++SQmcpiGkJnXjKZ3+8QGuymVDrruZ7iVCemlhSAXepQeAZybr49eggAZwCp
94+6lLa4wOLYBDEFHK6aexrxupD0PyCKKPxMTURalMGTiTZCAPeFQ9hU+UljgzkVZeklQywMqNTL
BQsu26Yo4XoUsTV+SBkWXMmimxci98Etx0/tq41Xx+ZM6cgFXO0gU6Aa3cTxCvyNCOQSJ65QZoXf
VTyz+vhYmCn9+wYFfJX/LgLXygr9PCyWI0k8azb9nJcV6Z0T7P2yEDRHjTOtnw6jmJ1JlRiYdHX0
hwkm0+p4ZrmWV2B4x5QHM5zgoi6VhlR+E6NoahlhvJcX0P4oQcC2CqKWrb6lWQ7eNmtvSLqXpKPG
4Q/wSeYP1MeH7SWPKqyQBP/5pS2Vlmz/b3n6SXa9loiEhaZ6E9Z/Ge6mYjluEv/7q7HFnk3KpcyZ
3HZPzfOWKdfFkQb7PrMDzmhlEL1itrS12xIL9u7gY9Aro514Y5xwaKukkplcVRJT0miMKoQ0c54h
Ibb4rV2KhpoAcqg9CloDgkctu2Rr9nxhHxbVy6JBuqimd/pVoplim7gRGdqWiqV/wKWaESyYCY9M
ee6yoEFFeNBuEl7ayCMb81L7JFUlft3xFIJj0BnBBQ8tpQXXyrM+0fzXNe9RGLP8c1eKbCAuLLRc
O4j/e64oqxeo5ZOfP6pTMhp1Ug9MEoXS2POwicTUwTygwlPfZLWjaOsE4tWXtGqoRehTd+qk52xQ
+3tK1xYOg7u5ZjaEG0P3fqziSGufiV9Zg5U6FDmbwqiK5ztHkfrQ4Ff/uZutmFHFZ2g7xXgkcKmQ
zHfWGzPDMkvQqosq3l8DVXI+SxYzH4Muv2mfFJdBoT4oeGZM1ML1gh1U1s3hjVdots7tlZZTP7rU
XUU+3n6W7VqVLIr0nQGxhSg8sv/czSyHNHZ8FMb4SYLz6pfsAziBabhOhZJccazx6W7ygyjtm2it
yTus/o21lVMD/OGpkbb0VCFXSIHzW1c/E/BN0AtVg1GJTc08r+DpS/OvOnhqBaXI6LLYWPaK5JCa
eWcRmqIEbMQpDeBG9XFj03Snb/nmd5NrCkKaONNoDWcQrke86mH+khP9gTG5acnB9Q+RiBr9Sedu
dgN1z0HBqnqzGxLtbMKNnoQ0vlQTnPLf2nHOdQ5aW/bIxEOMjGrDfgKpxrVBJQoojZBngt/pgFJK
LN2CIHlPibx9wD9mR6pKklhS542O7SajGAfVcrPHFdMO6W1IwkQSxXXYja5aS2QzeC27T3lDQJu2
fWk+iEnO/0kJ1BxUh0H3IV90Ej0w9D/uf8M/mM8Zr4VoSQ9gkkhm7oeeAMIMIW7KZiaB1yyK2Tlf
UI4PjVQU/w3Xk90GowEdebaASIlldt0WKb2JHN/wUIO9+mfLaWnhITp27BGVd7MhLPkaFnuLGmon
iIQJtG7jkbMPrlZg7sry4Ib+gxapZ1FxFabqU5DSi2irpRDGXbBOQDD4CkFC5HFyJapnqiDHQohP
eZ8ai/uAmSDg1K2JAX0KZ291HfKjUJtDQVY1EaAUOULsLuI/2JtuC/3MeW4CfvkqiLrf9WZydOUL
lmnXIX6wq7L2dBL5Me3B22n/mhMff5Np3TLEdc8UrAMgQiJ4QU9rkOlgid1M5OILMDk53HHRb3Zs
iDLY92E41Ktjkg8JwbIP+amUB8qMk0LXkWqDBlWiYoB4rCZpjLQDbjCharq7EHgtZVXKIzLOQBpP
vsTW7sbCPAleXVaHMWBDkPEq2ewMUYBNa2TsC9XA0T1O8f/zIx4VRe9cV2zpFqLslMU6eZdWGPpM
3Z53Wfzy2+uzBmuw9dbXjtgDkdSlDdRQCoCcJfZENt6Xj1lLtkCN2gGvJZVivxRJGT8pwb94ElVG
ow+SJARvV/SJ8BekpZ2+ZkFhQZ0E9QNj4eVjPRzVPK8t2pCfRtqp6UKF7OmbDWyvTGfAw5al7NqG
pkxJ8Z3+OQdBs4WbyUp/KahZYMMG93WzSTO/xSHb6n8PyzUmBKDped/Mk9N0RhoeXmLcx4zaeE3W
z7UTaDcX0Bbcf7d+L2ow+1Zx1dTnr17iuDBHigO6G1tbqlD6fRgwmlpNSNb+djhYQGfHy0JKNCGr
Rs4AS97v2asdRKgUeyVgYigBen80wJ3lB0EH/7NvjIVtXSDUdqnYbuKK1a9BIxqm9YRG03KEMYqL
VTrCMFUSV5K0f2L68CYPaZ9N6fuM9SzUS4P0piLp2a2GQQjLCg2QQoIQD8m/HFH7pVoSgbfNMI02
MA9fcgdTRoWgB/ymbms8O5SeafBwEJhB7Lbj7SDRt7ObMT8gQ0++OZLFEkGLymvUKlwXBOz6GCXR
CV+Y2OeCEj3ksbGBKr3khYl4BljkAsR6XK2k4orcGTWvT6d8SWG5KywPLvn+egVnlfips2yQLtNS
D5px9V2DS2ykCV4ioVUaC9cmmh/eyLQDaiey9yJCxVMsF8d/j6F6tDAgDMUE0vTqQYuux+1epPSI
TuvkgYXkiK8Imiu2aD/zEiAj6TDNYrZcDnfvr4P8kN++BdrCztVozDfdjhTBIbYtwUD921RImGQ8
Pl3inOE6Hd2Qzfg0z/Cpq/WxjjwY7sDAuHnjVQkLv0Fo1NC2rx7OxYOfojXQ5RFmv/k5YfVI+BkD
Hf9/A2RNZgmQR4OAy4jjk6VpKpQ8zUCiKrhU6VzsKo3m1YIlSluNSKhfCd7kC8dsiDAhjZAV0pwm
2UeDERxToOmtXn69Gw0dpAphVDyX//ci2rErEEP2lweED8LJrv2J9VBV80/6/LL78vRjCl2whR/l
lGZ//8Jawc6SscFWqxnTnq5MQctZJKoaUM56iWhZ2c6342JRH2hO9DezXgICn/K5KlBzpmc9w+un
KV3nwIh9l5F8bhtxmJRD9A1zin4WmilT+QBqOZlKMqXEkNTaOZleHqQOcsaxWyZ7MBBsA9V+cFCK
qXcBDaSDSoZ9jXmt8Y7XHd8SakY47RPnO3oKw4H7NHtVPp8ahYyc/zvPC/ka/Tjent9fpJTL2QNW
cb1yC7K4gi/EoEh96wzBtXe1uhOQ7yCPCM1VPQbsOZwI3Lt8jJw9NgaZAuTSqS0+Jhsh7rfHg2Nn
wVEabyfy7rKGZQG2Ez3oWG/NcfmbhKvX9alrH7p8H6eCIHfkhR1Mmx8dcehN86A8lFHfBiSKYKJn
hXP6pU8s7nMwLw7E2veFFG88Iam6xXwc0RiO7OcITl8pqEwqYKtkQTWu1Rox1Ze978wK34goFR3/
ggC+5xsUDComrz+Tw+72n1z6EhbfcNuJled/kwLz8k5Inuzt9hMt/rTrzPt4kqHHf0NizZBw2zC3
jPw5mCB4SLmd+p9uzgRFrEbm2NMab/gVpDh5CQPBxh1Kh3WUHykinUbZJxGICWLExRRmVlcPcVZQ
ts5dwc7KiyTUpJJUaTXrSC9ZkvmEHLWz9guB47OkgFvQHeTgwLWXB2aFHy1cgX1er2U0o/hfdkNe
3TGIt/7wuTlotkPG4rb3VwuXaQIXG72XimJhMj+C+MFT5CGjdrB5O2qiYvMff1CIFI1bqPk4SihR
Ds9JwG1zNyDA6gkAK6qaA4+KCjCsKYkkAv6biCnPZlRY64f/lXtVGDEbOvNYCamsrCuAbo9VRTtz
GpmkBH3trI2LK0NfX6lSYXpxDmAOQrV11OyJAba+ou+jjwgjrCAiijugh4szTdpsmYy2AXaXXfZ7
GNyhsbgkrNKBV8CwJ1qa8BIKBEPhPKouKKULoXtdjMYHmYpszBPGqBAYwnGcUt2wJ7FXTwmzArPS
5Cm56bxS2j8T7zYtq0JEB9+5RjeGb8FlF1YeRnZbCLySAukX2BV/2wUIGyuKXCfwJIYGWNMOeWDx
z1+HjO2CPDMTvcnJtNX9JSAIpjbDfkiSHWnDFR/h40zfGnuzHT8Np+ga+4TkL7lkGWM+XvCYLZrH
o+PIqb0SnBs5iwmYJmosnUyuZpx0Y8aSqFIWEsRe6xR4A98oYII9qEq/Mdd0jiXkWo2FoEYqmqWP
jrfAY1ereHtYFoRwUog6SZ1UPtTvvKoVj9rSnBwosHnARQCW0sEg1xj50B1z5jJEW+Od5SQHJGXP
/D2QjTN6k3exM6n/4zWDkwDIVHLRxNTEsPiv2XFUtk2rCn0NniioayMS0QasB779kbtBgU9oE/lA
MuxuVezja8dDvyjGpvw7aXvsdKovftrFYcsAbi0azNIZh40QP+N5+XX1AAjBKFc49iIse6MUN1NR
JIxet+awa2uEHrMHscUPXIFPwTmT2o696yRdtA4Wl1JglH4IzOup1SglE9+7hwUIEXDbdW0z++78
R19Xb2uPUHa4FNN367mMRWVTOK7AROcXbQ1rhScz3lOH0p/uRBNoh7amggJGYJ565uaz7KS/Bgbj
mknFdqOnKgu616bh/w4YYX1JR8YqFe2APvlAwTJwhvK1gL0tQZnQFoeVbHCSAeUumk0jV42I2yxq
OsAO3w1HmIh+L3tmV9QevlcpPiRtx02g+xmMwoAP7wH1l/x9W9gFDpPzj9AABKdgh6NgVmYrBgWq
uiY0dm5yyAOPHkZZ7BX0zLHGq6ME0evf21Ypnblatuf4JJjovnLMyuB0heHOMYnQfdW+pSjiMm9c
zmZxxrAwzy0lbTxMO+TusnoJGpfYKkKt3RqX1IlY4hdrLr8IsXz2XvdcUcLVEix4umNyRcNCft/I
PTItRPZsd7FET1faKc11JVp7/+KrihXWdNb1wno8k7xHrv6F5Fe1jLnr6sanCQRizQTt/FRcgmhG
o4geIuKT2ImPcrfGVi/VnryyliYPzOA2WTxIfBrz8qBJ3/7ibbvmE7V4Jv02t/x/3NkERgEJVP+A
PdMpe5dqerXHBsdgYW9M+sK+yhsaD/th1cvQ6iM/USJEjLK9gBuavoIP80WR0j+dz/6yspjazBcC
YN26ZEo5vOwCI+CgwlNB9lCLryYLUC+YA60KvknGqo/NdqDbSi8V2KDBTiY/UmPIAZNa/jpIBpi+
iWzmGJr0IZHknez+weJop1Ny+sTwbmFXIobfmh3l4MpnNCX5k/c524bk5z+QITDIN8zOU+LwcPJd
+zIr+TvUTzGIK4vHFVQLN9P/Rv7EHJuLBtQ3kLFNS2X/cFedPwdL6hKG5WapWAdzmVUuqJTQSLtP
wv9zJo5V3Sr4TpJcSM+DcmXdByPl4Z0qD45S/71d+zh3oXAZ5JqTdKVLeS4aqIApO+m6juRYnZ7U
eN7oFKBuCvRpEn0PWbrQXY67E+gRr6YouS89aGVtzvWXyct63zIFVqU1ZXmPTj7Xsf3+KlFFtMi2
QmTXc8qFxDyf53njOQjRSPnc7AbELMvzONlKdTqlG7Tkwc3ZpitG7KtVeScA1S3tVwnA8t+J8SVX
1lDHuNtUbIECx6Ybv1DScK3VGhNzqSETeyMeEuQcGMpJRsnCIQYQdi5+mS/fx9/eG124TcoiM4Cn
V8jonOABurHzOUOXH7zqVFcZ3CkBq2WTuFkSo3Ok7MznNPHc8UTgY6qK0hbbrCDbJxnW5zse+7LJ
aAguQ8DmCao5VICroUHSNlfp5E2VjuTKlZZt+q+prnsLgAntRqtNOj/HMxBYgVqXuIJbDovst7Xt
ls3MGZgqqhIeE56h3O+hgYQYlEcrhUW9p6hYrCguA8RPumY+HAZr4i+YEIVUcSUa2RWHFZe8prjA
1sojLxIrTOqeTTcy8/RLZNmRGdu6L1od4+NJHElosULkFq/CjCvvfJ9+VnQTCxuBuQfur3nheVhX
dJf5SBJFzPISG7n851gVo5a9W7ZtrAgziEjAxOWE6gQ4iCdOGY3Cf4sE7Oyh6ZoR83f1cBOVcGfr
g7BiVyL5qbx4vZvE3MVGtON//mG7IK7CGSNOM0IkfFwIh+OXEiWAHQiipKHRHXtq1BYWpyAi/gF6
Dea5+qXuRoCDAo1CG4VnbuC7tym6sbP0DkHWBjgDmBrXCwQvGRfTUhF6C8xS1UWyv15iXQr3gNl5
t0QxvWdtQfvDOLvYjj2F1lPE+ldb8J7Mx3GjGdTiRC4nfOA7ytbY0gY4x8YS9nriROzeP1ZKBRS9
U1cV8APHfu7W8bea8FnhgQD++kp0ytSzqbPqBZ/ZU+tlkQepwCwhzRY+JKt3MlGIKhRK3LjE1vwU
ozN73MqDhu8vBkdQa77dV4Lpiu4Y8YU8wdtMGgfTv3D9Q1BFfmw4G03fzkecRVWtEqoyrIHhZN6C
VO4mknNhDslovQgryC88Ca2c4nqSlwStgbCl2Dvth9TIPHmmS0gQ84bkk+NF89VhNMmiU6EwdbYs
0MtfT/wQebEKRN4GuPpCu/q5gqyQ4S2bZ7uFtel456LtTZaxNgnro0a/KxmWWH939Vx26c9xGIc5
o5uDABKnqq2hZPKZRXPF18gDac+Z/f7zrAV84x3A5XmF8FhlEcbeB0xwjnGsuYcojngiMJhA3qxh
+JVdFJs1D0duTNOd49VnWSIC4pJCCysGeuRLLzu/ZhsA72N3pyFVyIuRXLasuZ0dkkO28b95jXGi
W9zeooeyRUnlcqCs7maH10vYVYcFfriSm237C25kMSYLkloJoLy0xIn0c6bEIYDDo59sg+cl3VLX
BdYnC1sP550HR8X68Ox0fUGx57u+g0A2zlZVujHlXhTGjeM3brE1zEC2VZNooPqwG1OVtA8hmnIU
8GE03RDkGtee9YaAVRJ2AcnoNl3yDKvqlsqP2+mJb3cB44LCLkfFpdI5ciST023p3aFasMeeoYE+
u6E6CRuAXHiqRk7wWpXiCOoUKmjSd9p39CP6rdBpkyCcmPRok3qngl9IjpqAMieNoCCjeSZFvrxz
79nC1u46a1Ly4CYfKsFCw7EO6UAznhPmASYqVUVs+y5rONLjdwlncuXeZCZJIFY4V1JLeilWqxBP
t+rSnFTd8yNhH9XuqkJ+v1lbgb7LMTqzHN9sPwAStlqhQlNzR8SErHmw4uqwZhsylaTjKAkEwv6n
6B6poJsysPTxtkOrvXmeK9EftUzdIsTehoASZpXiEZa30EKcGY8UM13forMj/DJMz7ozYlVnpB3c
jqM1ypTWH8cSX3HnKCYi7fu/HjQTqB+KIXteZPfgK6vKh6xfCi5+sTXiGj/ujQXrZcSoPopGk67O
RCiM/TeVm0aDU3Va4iD0ezpuLMIe6zMPXcUgZ686X4PKE6ZbPrCUlZttoC30WcsmBcJsgU+VP051
oOUXwSItTXPqAWuZ2FVLCUttqTz92uNDW4mwUIurkklSv/U08EXORPZjO/NzIp0Im6fN7uRZ5F8M
VXwDQQ6tjlHimoQjz+/PXXfomuroNtheHw+pJSNLQ8xu/vtZg3u6SSSU0YdknzyTgMYMQjOhoXTR
ZRvHFU+AcYt8v0aDiUGD7KzvJhazHROECeIfTp9jNZh5VV+7ewnlGQaI92o6iVbhYlyi/4FW2d8z
eADUZXFPpH92aiJbk6dqMrAQhSwcbD7VM7F1zen0Zsh+n6jYPHuc76E/4xtZQ27OOJJHxJoq3DoF
2Uk/zwFOQrTq0YUY9WoPqX+i++oN4Bjvft98nazfsOfTPvQ1RZUVDWzOSvzT/e5xGEiEFRX1uM+d
3TCHhUh8rzvpJapFCTyzb/ogRlT9VYMgWGXcFKOcWbV2KK2QXa6y6LG/1gOe8ZNhj3+ykJsX/ku5
T5fjuBdmrWsbtzDmWeK3KpmmCCRaM2yahLXQBCpCYqR14Jqe9FzmmJj/PRveELd/SHpnog8slavE
rw3T1D7zIXaq3Y1eENXSyqAXXIdedDlmBrR69fvxsLdO0V+Tn4bEwtUX6XHwLstrK8sahBjNPXBU
/GMSKjjeheAxq7JVj34Gb4VHafEIfOSlmwNIdeduD+kMOf6ADl98Xm7BxBmf3OuS8z86NE7gk1Vb
b3BJE3Yne1tE8alIy/ZMhcHWcExe/q0K8/k7ziigzi6xkCkZIm4wWb3c+4IcTzA1EPKyOe18vq2w
lWuioe1f3riBtZIB7o6otJ8Lc7RlukFiQf/1C2P2PtxUIxXv52SPJ/XS/EU47fOUKb1XH71b3A0a
5nJsNRWrGZyF9IdtNRBJKqkOopmPvBqsd/8uCcxd3zYfDHkNR8D3J6pU2iEfWZI0sRPoMTIkURBR
MzgI0kNWU8Qx3rac/rrvHoEf8VsInEHFI9+3pNcy7jSqAD31g9+0EjweiVsOi4TT6mBf3SFYui3/
i1b8HZIEP72wV+B24o7Yw/qQ5UUf6ZIXYqI9/xMXAoMsaoMyfsFAVHaGWnlDKYcHjAVYhsUydKbo
6mfb3zCecaUKeOqd8FS1pyAhAlSFjm9f/G7/e1D85iDbouPjeIQRn7ZJ10QmqoFhAitSekbMh+2P
rJKfw+p9wfyEDmvb+7sU8GvoyT1KbjLLaBYrHxKr0F4HC2OhOsoKtj/m1Tv6O26G1Z1cIIclRn94
H+6HQcB5i6g8tmzvFpaTa1R3nuQ+XBO1uKnSlLFgdIEtBygyhTaZlrxtzzy4UtLDdbUnsn2D04h5
xZDpCUAZLEEOFB5q7CQZHuFzvAERJK0MJHK9ecFQkcWpsqLWDVsQo/qCX9jHEoK20VhWLz69gSsG
iDBforWUanEhJwaL5kBIcW7GiJs0vQRPAv8+gDHVw7DWQWv6NKMn0JYN5w0jlJDw1TEaqwAdV/p0
8iUXXkcXm8FmLErwgGlH/yd0vQnGU1ZcSeHkq+imjTuP01g2P1buC4r2TWGsvW3VYGg+CXgZd3T8
h7kIGVH4lipBxhK28f1iiliR/jMGOABNCLdM3wiS7Ar6c5wKz+npHEyIDwYuEPK9Bm6Q0Uhc8ep2
rQ30JBQGwWkEOIglJqbxmmH/xb4bQDlErmV1GrSwJZ0DK0muhxQpM5EARW8hRveE3VtJW0fR6/Vr
/ScQgwf/DOqac8M/ZpT8UXKZHml+F7FewValG0BDgFUjxg2XeETXa0EygPvNUSvmE7ec1jNxaVen
reIMyFcDNUOTYh7Hh5i2pkelUprNius3CP6kAH/DJcvPlCcUmRVxdXGW59Yf/InKy7deedjTYk1Q
JBuB73x2Xp52dUbKsP2JAzgb8rZlAhMJQkSm8fdzonGA/oKlByaQJrFQ6BWeM7rvZqsi9ROr1y4u
w/+cSdKJurvBUFmQBm3V8huCntyw3rOUn8IlHOWS2UKveR1b2/fTGP+FwlDLGFYrPoDcUkfaRrAA
TfVlZLD896OSeQJdAs+SP5VSarxHLuVtIuatePQORO0PGX/UwURDAW3yiUTBHu/3KhPMToMi20WV
xUq5Cb8xHm3pF/4p8LwOsyfq+vCNsWF+OwYp7L5eZXBTgTlZB4KPG4vteuZDmHtcE6lkBnCn2Qu9
7k7uIdaSnGF9yA+PYk257u4vH1cnzbdzBODZNK+FH1bBO3SqGj5Tew4BgR42IhGWXgoivGKSbcBO
m1LUPXISV78zpUuGx8OO9ZwBbgzHp2qBNRKuTgxoJ9tFU8JHlJwe6IuExkd95Cu1hod/UpaWjY5X
HZc3WVjXAi7TeJAEB9Axff0+oVko7qCoYqt5DNZfHl/mNJKEXDT28EImD477grF8cghehdBwrTv/
LrQ5h4BIvTaZVjqIJGRwNd7Fkwtp+c7MmIsfQTyMl+/XTBLAMksQw7XJgnNCE2CUUogaAgklW8OK
mojDQAVTJ7TX2Teq5sjnHfxjRTCzDCMCa4BoMOaUI2AF+WoJ0xjHJ0fkt+kJEh2AYmq5O+jGKN+P
C0lJ8mHe8MN2gOEAOcHflz92dgHKVEYQPtmW6vJUeGhCpF6LceG8Tl1gp2v/mpejP2ikMkAEPavp
iFHo+HJf97DGanRu92mIze/NV+GaywGr1VR9w/PIRICw1r5C30VLyFPxIpBOmjUm2h8fXh9jIQmk
eSp4+Z/jVG4FS22ZV88Pwbkd3zjg2X9P5mVqJq8FgkRuhlVChiW5axpGYBqdc7rxFioK3K3AQwo2
TYZpxQ2+ptx+P+nCfc6MzI1gEON7/1stC2yhrRWpn7D5H8h4ZHbFywLWUoYNRVOw0v6S08cEnq5l
9gv/4SVx2yX676DTLEX0AmpMMEJxe88Kq6fHIZQZEfW7FPLnopMFAoS6p+s6K8I1N5lpC1KI5ZkK
OKSUTHRVlucQkZfEaFtPSTqkerqMHKAW+bLj/lvvLg7BUn/cKkskgLSD0Cd85qBadcY1+WxqZLba
Q11/phJePwz1PMxamTCVL8mS6iuv4CyCduMhlrfqEIXK3iD1MfH0WzEl9AR241hgRp1hv9iiBfBg
eQiZuVZlx0m6fKpabI4yvUvp7nejSRyVLbtNW9P3ZT/EtN/TcU/llQkXZk5qrymkNt6h8gx5yRc3
MV5NEH9DnVj1+7KjKkk5+ImdLlaMkQyC71Q+Nxoa9WCNm2EUwOpPfZymQYLxf9Fl5libTEEvoB4O
oJ51UdUDAd6yy4YGHrs9TJFzlojCHBD/GqRM+8KQLPkmvjvxye9Z355NxgIjSrObIqFovlJ56xAB
h9LW6xcz2OaUUe0EsyJDl+cqUWfFsI++aFhL0m5PrMSBWECaukdeqpexu+KRoun1dFXqw9qS1qxq
9jg/uOwY3DVOI5esj9JK253AsQsogzYio56PYDePOiTxz7aC8XN1ClBMDY3DBof44Yx/u6GbLs8Q
AS8nL9A0GCjnZ2aR/SZd3AUHo3pOtpa1qNrEITgughb1QX3bf57mzKRr6/ZUz22mBfdzzgF05mWi
1HCT7d3lozfHGKLnhceK36PyI2sbbg5mHRiyFTkg20OO4RfOH1LFfq3eIkDiiyCUToagUlBmz5zQ
PWNE3BlJLpTDdZweYjZ04gVukWV/3okWC9R3wd5kS1K/F9izaPLCLSS+nr+Vl9gDbPDF5fAVA2GX
+0AY4pKfHeYg0YlQhBlFdisCu+2+elBjB/0m06GxYJ5dpwM2oycgTpT1yMhgbNtjBdq5AKUOdSMv
QXOZmQw/r1AR53UeYjc5tFP1n6DzsZG2x9DHHpgEf+WTSxZgnmf6tWkH9senIMYg2OOMtXqUKlJD
AmCNJwPuAXFBH3zMIdYY+PHEN6dD7dD5wXBOtxAH+YLbzj3Av9aPe15MuB1+KGVZNDdtj0P2uhP2
M1+OVXBWaM89dmQ/gCi2VL0NPQuw6MvURcRD/cAQbJR07EnQ3DWSFsH8FPyXW12w/9wGv9l+aQhr
O03h17uPoEAuLdQQDX4ahKnOXNFU2OGnxjaCore5HpZSLXoH8JjTtGMtebSnZ94n0P9aoRyNfE+C
FcBGB/gXcUtLRjSH7hHkn70/Tv5aRBHfdvSFeOxXByoMCGvK+wrK5Go60OySjpxs7jH3JKu5q4Bv
tb9yN9+TojW/AcG9wNS8avfli88h9s0/7vy7dqZVn5Baujh5ZTJOXGqpBhhFg767QTQscCRAvy3n
tPgQ4cQw2xAFLhfgZeLp30WzkmUtUg7vFQHO+ZS5RjXYpDsbRJFdRnHvDbnFHM6kurePHUebgPq8
BaxQ3vKgsc8teRJcEIHdP4xeZyRqrgIB7N/gIB0rCvejTioX2i4k1pwujRD8LHBi7wmweclSDejT
damvDV6nniuIzIiQji1HLWWgLN+TvJ6Jv+4PG2QJHKSDHQq7ZXjwtJNHcTqhPBquXRYJZ/jH4foZ
sGycu6hAn6UMGz9dP6L0fU84YvtZVG1CV2y2dn58X9b7cpvJjqBMvfCkW8OtkylPSqHKdqJ6YvxA
t6VmFPHRbyc/cMnlRLtwBghb5BG+rbVj4QLbQeaPIlVnin1rsicLCCGOcxjPlJCP33WC/L0f+yhn
ethc47w5duD9x0+VpNIez5ZXAQyo9aEvJzy/PZx03C5I+ya75mKE8iteem+iiWsy+pb0HVWdmwDQ
pflfGEVcgnhhOP2oS7Hv55nBLFrrZ68ZDkLURbnG8y7O1cc36baUP16uDI4um7lhR9JfBo/+Bq/4
h8ov5HJPLPg9/Y/I5vTkZV6wXPWyRZ0/eq2Fi2f2omPvWHWJgRN2FUIM0WRdtCNMyUbTJcPR7ZmJ
eBZM/5oE6NHY1U0C9zVrejtCkHC9sSViU1ygCHiSgKahrUGmMhrkDDmuu0/fWGU1Rq+khaVIdapZ
j2D/0BYWaqRu6aFWWutXLK+l+u75+FdwrkvaAuirEUt7Fl2PZktorkB2e+qOCAkkyukhXvEnm3CN
0p8zU/ouUeApzk5xo8JORAIXqWg2iaKtbCEbIAEkmrWFw32zTmIH4Srh1kbJP82QFr73Y1im/gqx
Dcliqk1hl4tqnAZxcqEfU+e1mG0dAWmlDFtm4NncbkST+uAgVkSwJYssZcUMDV6goDZbtvPscwwI
FRFdumhewwMgFV77S50Je72//Q5e1cxBe1CfRO4dKcmWkIL3xL0cJA2Qhzq/HAy1vC8Rm9XX3zQy
FmJvq/qRXECpxGq3Q/P7PAW4B1k0+YnuOQlaAXvYBJFpOjgYO3av54yGCm1VFGKQYDAxMhec7Ryr
V8GjLSE8nRSXwdqqHkLo523hGlKF3Nn+HdNeB7hqAQojbM9UDZmHOsvZQL+jmzZtDydyCWqFjQ0x
Mh8rarxRm3vsp+lvt0efx2qzTY8ylV2EkuSIhCQHigHhMdyyt25WHTOitsX+OrkumTb4A6KE/slh
ethATSV0aifffClYBNJbBLu6eEP8HS7zmSd3U+tmWuPvR4ZlZ4gOgtKyPqtXdMzfVaG4DhZNesCq
CrPi1TM5/4LUJXPZ6g+WVvoYVEfeC5JQ/FbsV6Rmbc5NhzaHamzizg/SNkvVWBMThV40XjVM4ySD
WT5o4pgIxSjzdlK55mBaE4N5LfNQg45T7OQKNOErGXxRv7edpwHs3y1mf2Wayn6Z/szQF/j7dkft
y10MegRNPLT+i5hzwRl6Oe/c4LbilJyirbMNYsbSBdoIROfbNyCeDL7wrbcfgu++mgO+91Ahc9ni
pAKEtCnDH9Lx21TkxVLsFm8G6JWlLkGBFWp2hHnWZivKpTBBELgYn4Z0pnqCtfvuV6LbwQXZuVEo
W7l3of22l+Sdso/ZK8tkPWLQmbPguhMDpZ1VRT6G8d//C5mwlbBxihO4CHUc8Ue8fLCw1mcv4srQ
Dkn2RSVK3q+z1unOJ0kRD/+oEnOXkGcyFOFaox0WxIO7E8Ucdvwm9amV+PM05S8RZrMQGN1m9Yvy
0VascmYpoZPTrR24efPbYNLzQvepRtecAqeCupd2YMQ4PkxC23TsnPpF7TKWEt+HBLWHwuiMzPmA
UK2cgde5pj89YhuDPN4Qw/O6z6BMWDbzEwDQRMRA5O52D/ASiG/KqHBzyAKD1XnN4+oT4XUKNMDB
3IG3leZaR++BZ8vdtAfj5odSbPwgKU1Qv66dUFwBK9fd8W5B0PjjlQdrHVJ7/cJ652NAsCy5Exun
T5diX6aBeM+4azEY5dASXI/dthxpoAqTCZxLSFQhGTogxb2Tt0JFtKOdjFmCsmL72/LJ+qK/DMnW
2ragWWYpXQlBWK6RU2pko2kPMe9J/ENpBSRfgs4LG9UA9ABdmGiILW9zW/qx6mfLlvJe82Nvifiz
Bthx8APpnBlC/+MexuUuG6sMtuHNZkC7qBjy5d/QvzqZYgeCdkeMlfjJVCHB3WbhoNxH6xxt9EJM
CvcfonmyRquUFp1aIyQqsC2LUQGEA0QhsKoUjtl6RXYIH49D5JRGil+bPBWsbCt4Bg7N4lJrgQv4
95ckxwJ2nPXht6i0wZVdh3HnL8Qg/vjOxMZDJNJNEucj66nV9TrLReyraj3B1rzl5qo2iVRTgu6y
NNKEWs+sJaWSwS3jV8Jm+zTjz9P7mFKnC94ulU4m7T96KKj5oYJrn1Om43Uka3gLuYak6Vc62gC+
wFv0lBjUFfJGf8+ThKulxPqMR5axGBxM7lqmXpHrY4X9AiLWKyRNS+Ii5ushLfWY83WFm0xJPABO
7VAhZv2589H4rtyFF5oS2LEkQBir8yC9qtjDWzYN5/5aK1Ln4qI1W08Zi1/sMMfK0sSkQLEDjp7k
NKAqnTf0LaPgyD02HAFaA0wraYfjKayBjtSAnCCAfNPThDrIXxzUjbCr3VazjlNNDVea1JmCJYeS
LRbi5te09Kzkr5eTJLR4khxVijQqmTQAAkU3+ThqqLbWoL3o8v5u2DU3JNRuzchEz78ARw8t0JOR
ZFh2MP31G0KEHrxY3NGH0ZF4uEbVfJSosFm8wHrwxbgNS1DhpgeQ+KwNGEXcJmgkFSfpMLU8nS4K
oIW1/JUbaHYryqcsr1IrsmLrhPucwvmsOxn+uEKKplPpm1WXHd46u2kTD0jx5h0n6ehxe71AVtJc
R5Bqnefw1h9SVe6xqWVPQ2Z64h1UX1DJQ4+w9V3NG9VcGI7l2TJMXKkTbEnUbCKmP8jEn9jIqVBZ
2YeP57/Y+bl1VRaATojWpKJPkRtDT3veCoShUwQzySp7bDBCWmdKOSI9+sUD16rLJcin53iiS1zP
MI2pQX6JgjqsmAHHryUx0tcfIHlLGciJeAhITSN2i9RmwCXxdR2DOoMA4uTbTQ0Z2E4T2K3GTb4A
dVDBZxKM3n+1vZ+gCDVPFAYv/q68EQPPsGKVy6d9i6LnELWm/CrOWWLiG9Fkvxr2lv1E55jfzUQu
WEyZEU8JYx+tZ0Dzj/IjDqv8gCwLJQFv1L4s/wDIb1neZbYhsrEKa7Ree5ceRKwcA/Of+eWQNjL0
8rx3b8E/417N+KPvjbTptG9mJiXBRaJUO7zvn3+2EotucYQupj/NPFJ3xrARvZHjBDEMzYRp5qPO
iA5UJx80Qu/CWTHFHbAgf4W1TjtY12rlY+1TZPmOXobX9LXdfYv2Y+vDu/AFI08+w3e6PqWwej9C
u8TdVV4MlaJAh2PMIGwR3tPudhK4o/HgyjAnuoZAVE9TNB+fdLQnDoNLlYJzP69awLo2r7XY8gGt
4FDRsqkLFnwgKTJb6Pu7bNOz8Sjde0Fgi9jLZ35Xyyq2j38vd16oLogyQ+oBZzIxg7G1sQf2lWWG
suF/0AIPRbiVUHKDjyDdBo6+zv2TXLE7FSgUSoW75qQKfFFgwcGi1sljQZEqoWRea3MqvAHPmLhF
2mXA/jyvs2GO6c8GzmUfUxlmjcf37VXAvsdnBq3ZlJ7+OJS99dmqZ1AG75m81vmkHmOvUoE0vjBa
F2ez9zUp5adQUFVI2GkANosnMDO+hOHydKi8uLV+yiX8BvK/TUMkqjxlr3S4/YiHvller04pTGa4
PAwj61UpVdoGEwPATuPGbAN0CaV7ib8XA/UhTZeIhuDvt09LKUhClnp1MfBXs/swxab3oRtOwRzY
4XAPbNSWJJZZZUA8IyVIBTx0zi31o5KPYJIM7IvS0ytk+wL4pHRt9bqWPlvOp0lFsWRbzT9ruzpH
iQviUHdZzPzY7JjDHO0k86AieQpAFlK2G+mCU+DYN1FZF+z0Y77R0arM8QpIEz2qwgfBvkaw0DhE
bxUiIsm+6eeynTK67fmaUO9+dEXhJ4spJIwXgaS8YaErxdOw9s4bOfesoQPdqQ18+0l6yDyu5EU0
oh+VlHSvTAX8oF35n59bcXdWIng2awk8Wp5GjMjmpbqIaRsN9wuEeJMUEvFuTpW21G1wklU0Ve0e
zIO+gI639cdKgVx27EvwUGvnZYGB2z/BMTLKKcrcKimGxEol+QbAqF1eL/ppS2Q59tZ6f8uZn3LY
99aYGW772VfoRi7YilimomOO0QsDD5PcLksL0qX/nLc73ncPTNfenUYuYl1xJRZseXj2oxYscXR+
eJn39U2ofI2Cxb7fQUwpmp7aWm6/SLsYgtGxmpXWaTnpDIwM9egzMdsVnL7jQVlO6Gj9oXbwZeYw
ALw7QuIwEmfnG+7nGH/xM5i90+RK9NUb4W0XJZxcePIzH9Zy7iRuPdUrXBJqmd/wl6iD3qOWfzs7
6g8xPOxzRVk5917gC1OQUqE3De5ltg9/UeE57kJJj96dhUDxJdycitLHX0kfeHMgrlW/vy6LlsFg
Hpa4zWb7JrXtPObsTeclU1sSumldqk/8woaLTwykdCvk9kmGOsWtFcAlsGGGk6ohMdlcPeZeTxHK
iPbDi/xnJXZaEqbz7KZB4SAG5NlqUnhB8RuRS4OP4I/sjw0bdFxgneIzPVmXVfxA7m6FlacGXcQl
RPkK5QvfuxZedgjlqOV1GyMFzxq6MAJejCN0mPvresC6aBCOuJmm9PUDkMiN4vlDB8iF3HZ6gAYl
jyBF9Ud8F9ObauthXBHFd6AYz3ajTljDUdVMeUOTjvtloW9HNR2DSLEN37UXOoiy4jkxuYqYcuTS
z6ipSWq8Ucrx/NJVC+IlfSCd/s+mFRqs6013pQ0tnwD4GWOiavK1+I5PSiLIgiReAR4Tuj8TY8Sb
2fryYWrWkCH7k4SAcmzPZaWe7c6iVFwDsPf/nqqkcj+38++8yGWgXa+USJv2vN335vxlKJeENshH
hVG5kOunPNrEEzNR8+WVcU67riWlD0EtwzCOermf/MRWI4kap0L4STxGM8iW0d2/pE53tQpd1Azy
vMEyCbBrt5rLZxTPFpeDmLDDuq3ZAZLx6Bdb9SFALA5RRRM6zyQzlD9FbYjTfCjEYAqCazJhQaYu
tGpDDDLzmlL9MHwrQVlKukdk2bK2nvdj+7kGc30IbDRqPg3Y3S18L9dpQqzwuVbrJn6DGCft/Qa8
wLlAdSuLMhT4bvi4fG6tbMJpC5n4qIMl/yVJSgf3O89moRid2blKX1UNnjQD03ZPb/FlMMmEsemJ
hrszODftWGIj3VU4T6m0b8VKBC7HYhUFWcBUhPQ7yl7ufpJBZb19w7edklVQ8FiF0rtv25F+iT0C
PnTA53XaTzDh9o4UkjFbJmYrGF/cAq1O4NT+17F22dWmpwdAiud9nnykNL2AyeR8K/XWHr0+sr3J
r0LHmwGEQx+bBlrGHJ7R5T7wAGePkySD81hbY/6V44JKXAbPk5U6k6/E5brK7tOLB9auloz0XBVn
iK+KcJzEJ2m9dDID8C1MC9JMYTYi9FQ31hiQUBLXdjeN8y5PUaaXAUonnbK0tsqJUm7A0lVcxd9o
GewtKxit+InuL77cyUmRc5UvKjda9MNPGDTw7cUQr4FsSM79+hhE/xd4lbqbgVwgYMGlZmnJVsm6
Kh35qn1a8GnXPqWSja5MCvo8LXMy0Aub/Vnay2sKzJcIv4SK0s8L+6gXBtpAT1WQIRbJHRjtngbL
oC+TB3KplXDO46r9OA9tj5S/e41W6m2Iu0YDWWI+URb0BXcdGD5NW32saOWHIQxEpRfJ7AHjnMwL
ddcwQRSnarxaFJk1eFFsFrHI9TANwjLYZOjW1W4oWt8Rfyq4L/aixct7r7ov6bzpl8qBXDg9+RKA
ePISrtQwQ0zcO4KVo4CAUSzHTnpAjspwUYdbdAgLFLVRRaPDNkQRBdrSu653D9exAaUPvXaT0U0E
120MuMgyIulYx8gdShwsq7ISp7mmAXuX//ruFAOJwhR7j8u3p2a1yR/Oru2Oozu3f7QyrL2xnRk/
sEZtfZuymgF80jKgrUlVFVztPpP+6VB3MJZKQH5711n1LIAvv9bUy2dCJI3Tzb06rZFGy7TjC3Wo
gnh8G7bjcZww4JLZj+oWxPeqpQmubDFYY1+INxdgREwrAhcu+nhB5mpsDyiaaxRQVjpGREgftqQ0
AgwzduoPnvS2/PI/VbXW737zHE/w5z87Win/XIkoBSNQvQn0XMyVKZfxjNBKxWvwKOo5fdbCqfBW
zbr5+Y/RrpefyGtfjeowra9vikRjFm536RCYqK3y/j1kIuuGOr8wdAk9AhdobN1X9BsRlg27rXMH
gwUfCQ0Labx1E3F6TJliYPEvcr+9N6dXsp62CsCRsvwMz/I4WOvBVE/29+mNxlGmwpzYCsFpyxkf
OWZ+1K0tRjcmBHVB+djEguAPCHGjWXheoTPQPHX/rT+gcNX4YKnLWVZ1jbDg1yP0nhuJB8WZT9bo
G0UXP6BhDTTA39E36w/lR+5CyQp8Do/lEilPzYCpdtq/blNKidRzXSAjGYmXOMGhCylN4Gb9glgf
uVbhgtkk7F1Mh8cks6UCe5Zy9TjBQx7oF7sOdAPMYDHmzPtzUfBN/JzR4yEKsbZq3uhD+t5+uD/9
DZCSi2WrXqGUgqxdJyOrAkdIkfWW5neMymZ6jg50j6gxUP9a59RO9RyK7tdFX88DQuowt8/vUmnn
hyyJXU1FwnTMQyXax6iMaZ0EE0tz8NPvAYrL3b4mQv1VI2PWD4tlsOvnmatW+54aXQDDja0UlbrA
ymkuTXmRMoveYVpWL8MPt0t8nGGaa5qJQAF8yE/GRUXNDgDh57bQyUu2R7Km1UslwEcQbAg6RH1z
cI1JIod9J3MTO+nlI25HRgDF1s/Z1ILPfow9Y4Cn2YD7Igim4owZTJLvjHMcPMVJgxnFVexkllvC
8xISTB2eC/40J0ULiAVXko1S6PR/RyPLUrIvYMN01ruCIR9HqESC/m2ZxDOcKTEcUZNrWAkQJQYy
gHWW1T0AbveKo8BfPx0qjFPIY8I3AX+8BSAUpurtyEHENioZ79r2OZCXTVc3NTRy6j/OTx40mx1+
mJi+nHOpKycpWHmMC0GbjAvfdqYrrCD2BkwrkST64D17xKNz3fJQsUt8On6OJF0+c5MNpU2x+hIi
kdd5R7caRjS/3kZ4seVHeGH4QdJg+pcBXA7afDsHsXtJB/no2a3wgsGuEuwG4JQa7kbS2RyewzdD
Xh5Kq1d0PxjfE3rFX5Qy9Dskz8jpCLSyAEs4DFQV/QIdEfSIYBZCk3HKUnYHy6sZ3PsGPm29JnZV
gh8uldE/skvuO05YLUML7X6o65IbAhu/n761c/E6Ns3LG/oTu6kUp1vGRFnsqPV+5bTQri2iRNMr
oRu4Gak67YHb19IXZHz//4ZRCaD2RYdLTFrtB5r4tm2VDX5/50sYicfdEId7MM5DYQYstEJ8ibXn
oM1VOnUKRZVAarc9v8tbLJEkYMXl95K0rbFsqMXFHK/I+OoOkbihKdXYg9hMIpl7MSlptXZ4P8Pd
hMHyqEYmoPhFXBOSvVaDoVZZqyZ3rOBGPRsTHTuXjIhHM7foxjugNIW3Q3aMvx91waJftNyqNjr6
lRgwaSLMx7PN5QtU9TvAYwqK7MGsiZQDl8HRb+Mvx6mxjEbSOCde5cqxpy2FCA5c2g3aQzoXmOki
ltwr3KQYuRFCMzn6P4tMNN/qCjxrjqFfPiAkLQIRO0fvWToIghkCGduI50RzVAoLGGOhQSzo3NB1
ReHaMzgy/BY8m1br3x/Bq29T21ggYIJOAxjZskfVGL7dmlzoVvQKeJvNvZafCoonCBkiOhEfTfMM
iQrkGCopsTUcLDq5DRG1lRbCMp4Jq5sgOyD8zuLMgb5SwBxi983Z5UV1FsKGTDGDrv2etAyQCTya
sEsmZIqx9Q+DLEOBUD5ioJbmo7xwpKJrn/yPi9t8kGJSn8sixoUghmU4pl2874UJVmkAAJgaghff
+ED2k2tMB+2Opw18uQ5RjZhI3C6GVkXCPLFAeXBVceWTHsURQfPbTnHB93Z6sTUMW5VTpe807Qaz
H9nLlk4HUY8OVQhlgicIkFBqDYM23u+OtrTFMj1DKt391SfupCTMDdYI1syfGGYaqO9UE8KA7AFv
MPrximsTPPaam+ZyOWykia41QabZunjtxqoQRnCFvaCGA1E87wFdVGTKDwMgR/J/GfMeyL53okq2
BL+H0SZVW/mqCeRip8yRYwR8/6EiOY9SAxm5bgaxwtxet91IdWM2Bed53HHRqRF9Fl8sha1ov3+X
wPdOK5XNzUwLTfpBJjoVSzw4L/Owu0B7rIVZuqFp5EKqKH6LX1L40JcJQYwop4BuApDYbU/du/qg
qzrgxgmtQLODvhu6Wafz2gJp3dHX0uelnJzeiCRS9evgo8F4RFQB22S9a0jQtkcLKpdHwSkgyyxu
e4ADXQEsbYXCDLCqZpp5i4djWj5jitx1ZXDj3FYCWoJ/YMGEbsO7+Mcr1GN7HbpaElkU6ryzuxcc
QVPUHup+IiYhMEemXR9EjrdUujPZgtf9i2hQpo9+HckDIme39BnUrcNe2NOePpr7r3RIPoT3MVSD
F8CbF7rXigwnBuNNmfS1vXSwF145X3zg6K8C3h/f4tEbOiZiiehY6qX6BXMLiMS6/WHNUZ3DwVWM
jNwLAlhyJZu8l7z7Ch5+PH3zrGpOaAJGd6Ewsry3bonPP6PJwuKJyD2udk7K1X0ifMtodAkFfZKE
Nt1OZukRPvBT9q5uetMdCz+18rwHXzu0djyB5Jt6TVI7fnsjswGKUdNmuPTJ53k+FpvFfL00/Wdc
77pGuww6DH+CDGAAMnox8Y+/Bydcklp1phpXu+5YbNzfb8V0GeuDGA/FYr/XTpzaFODzPeFs9c+m
YBvdV7Mf/l3ecGJABnyjSs/u6wIP68HAXLfOHTMrhkvMskTKY8UQKFzpsiDy69G8BcBoJq0cAHkz
gE/h67REEWZ7jq5Uj9rQd0sKZ2bwtBrRPIsYh0/fY3+Vi+oKT6gTWAelFAmslIUO4CfnG9B584YG
JNpMMBooT0tr9j6323FaJEuIpastIZi7QY/TNhW9C12jEbbYr7hJl4hwaoO4x5yJERyvD2/XfUeX
HQMk+Ov2LDlyM6+Pgh9oZudSitRxnLlCbAmcHx4ROC6iuDKuMbnG+ek7BMFYwC7BPtOeYx9hFcOH
udWBQYyNazm+jEb9MrQPj8/83zT1csJFy2EOqZsZBchMTaqkpYgEW8unsrPhuy40uyx0d0qDVJ/y
+EQBNd8UO2xOr9ia6wvohp5ivfidWinR12/m7odQFnX6x1e13KhP2kYZFSZh5/N6309Furzy+obH
26DC7EJ+XEGzM1AMwTARafzIeZAZ7tSrDB4Iftl7TGGgEH8YdVQzO7hR76aZPDqIqEWZfIwtVzp8
S67/allU2dVhGugCEM3ZZwvjnhkS7/ETszcEED2rr1EWcbjTz/z35nO5tAvLPuVoNTDK60G8PAP2
R5UwHIzZ1bDqN/AkCyxTf7FOq7YbvItB+nVtBNfyXl+c1YhrGM1tHbPT60uq9Xj0Cv1Bj3JKM3OB
WE4dRB4uetgnz9XoGjnAOYGYWmHkNzAeyqFqzCstkhkXturZY8HQELkAqNO4wp574/iGB+Z7EKzv
0n48f+kqDtSpRRfoJIyteadtYIPJxCodZGErGd1iDa00KIv/EDPWZwabGdW41HvjgS54aLj0UV8B
P/uECB2rbeLbl0wqT5WPDyc0hAnLMQ/GJ1XmG705puDdix0Iv1yEBVvXpLXlII0NIa9cubLSqoNI
TmNcXz9LbSmC7NTSohJrQvZhNj3AHrHQEcDqiJAzsOVWzVVH9nh3mEStou7BprIAbSVpxGAlW/hc
M0Jfw4eUievRQGAXHRxbVjcAqMm3Btj9xkCx5gW93BQiCKV6y7KvtlvSNuAK3BF5PISI7HIx5VYR
ORMH6QABSlwusCbs/Ft36wPcbdY8ZY64QxefiQ+XOvuXpYqVnwE6EH7BCYRy7nXKWzss6gStU9VJ
tot85CDqZT1wG9BhlIQiJ6X+5S89QaZ5mSBaBZ1HXiWMWQRdB83YHVs7k4d754TA2xotFBDg4uG/
aUwnledKDGOwvdYY+S3PJM13YLhYAg2TY8JBK3zMwF2btizreOUAvVg6Y9JgKdBXpxi8M1XegPWA
B+WGO0mOLif2xlylLhmup6yfwp0RMnfTd02sha5tANfshu+RYl5I1uhmG/+hMB2iUf2/VZdvXm7d
Djg/EDP+gVPRGXAf7AGY2kHNvtWeE6xO2z+CJQwA7U/g9AqATqzH8lVvhAZ4NN7+xEz/JXGg8ebF
AjRPtW6f/9NacHySjfWv+QaB+OsK2lR3ptl0UJAONeH+vTws9fMEoeDbKca6DuMmCmtwEBSSwgqY
symaac//OEFgGnY1vgJYvVhbphUkMYdfk31U4evdGP1KZbHPNLyucPApAC/ZfBkwF4Gd6ftrKijR
++mWNEAs4wCnmRLm+yEIKtaDCBN+UdmP8PciK681h801AHqNIPGmkAPKJt1ThpPRlXfNLAssD53L
EFbROYOJa2BkJbxjMJfDi/k8I3p8wdPh6PHJCrXfcwYr1vBcHjTE6oRnR7pnl0lfm+EWj0pd+AiX
v7U6+DmeDLawO28f1YEXDnKQ8uYz+R9WKZnhI+yIuZIf4VQjqFKGDp1DdkdRraCK3+yaj07AZL6I
I11bauIzP2b43ULGUrO/FCo7jvrbof9VMyH8P6jCB9sfLFLHeScJrU/heQL95EASqyPdRt0EWQ89
82x3jwB4g+h/qzbrezOUo7iHKNUyn2g6SvJA7n0Dbgx0MrriLMMQtL+7AqCB1VxQtmHdOqYEzyrL
hhFqKIe1OT7uCyuxSMykyX27sWG1PHpUz927ruaTSZSz5jxe/0br+Zf/7vphJBYH9b6IQdQSYZXf
UXYhp+EDR+hoqdz0H5CYU0m11FW1tAH35weFJYCyMosNFN8oTdEWKH/wmxdQcgvRQqjznnpx3Mzd
MljRWc5UCrbmrav6CLD085DNdMcxF5ZtoLJUBqahzh5vPd+o9Rtf/9MyTr0hBkEVPQp/AHDiq0l8
aKoKA5qASwn+P4fsK6l+34vD7OUCyhpQ1xX8S0KE8HCEeQJ5JUOmEhoBnVzAsAzZp+8C22ZtUSFq
2FnrTyc8RadDCksnZFvBtQnVADiq1e4f/VpNr0rvDP3ewCEXPz10B8zuTg9paBLOQ0fbyJwyon5o
7+4YtP9m6P9XHH4FKusol+q5d+G9WnR6cIWB1jZX+9j733eF7SDgMAW+KbM53tpHeuoafYc30tXS
dP5HrxU1U/VgQfiEtJ+Kg/BKM8AEeZk4nn1AAH+mpxhem/NWxRPSaSBtRTB/l3sojT5288vs0iYi
UibRMQrKwC6ArZjP8avfahG1ttjGG0kypCu1hIYgRhv62pz51Jc4exd3qyASJIU4tA2Dmw7FSC+P
MYejdmwoIFzoTay07hHVvDw0xn/0ZCnAgTohsb529Had5rRX8E/aDGAFTS4GlNHqKN55zXwcJETJ
1C1gSjoelnCP1w6e1EWxqjcyCkmfEcocl1kmRKTGekZd8yNZ7cze7KqQkcgd4zAzr59/Hkxcw/3V
X1ahriHCKebEymdE7CBVDq3QfFXUFLxQQGhhiWZ6upQV3GQwhvW0RQgc9U50n5V1i24/FZSnBUYy
mWFRSdNz5idfELI65lyAI4fVkGcncSSdIyQ3CSIJVWDRAPG70azNe1nH2dylTzTSvH0AeTFvbI5C
TFfW1oyd/t/TskY0ploIPhVzltmD8j0DhO6lolcycYa3V8tZP42nthg8OVm87zwb85sg/q0haNrK
s9J3VcJmmlE8jDonUQBaw9T4G3sOMl4uHU/3IZ84Se8PJbem212W0LYppv0zX2jHlqwXZo/tQnqt
2ieU3kAcyEu0pLL38DEYDw38Ilp+QY9gJPoni8hvA2RGxXUPPuw2knb+kG99g0Bz+eI+RRjOTdPu
FDuqN65+vBvQw582t+YR6yW3fk9lxx/QPxbcn+6lOu8ccoGUOUqUcIKkwzV72SWhIkudnQdI7DGI
szLReyE1EMB+f/unAzrlGwEU9aKgBVas/WCxueSELVzJ4Vs+sV89FtPrGtuVOY70QtfAfhF2X8TI
bsbXgcqdiDxGDI8gMk74PUW36SmwAYKlbCpPU5yB+w8gt+v1Cmww3+SSxy5r25b2gokmooWpFhGZ
h0OWF3WzZnxYcH4xYcHqrAQxy+fMr1yp8X0+f8zDv/BF8tiW3f4cyVPSNuLtKP1VUzgluogLpOFY
94XX278eqFNojlK5+UW66zObPj8xNajzBoBBruiIvp5erR1MBIWJOnRQeGaYx5l7Jgv8nNTfeMg8
jw3BJH+b63E6s8Noyw6Mo6RbIRDZCEjQNqkuPdigb+AVrP7KltWvBiPjQU9f7XQCp7abwx8jahBf
bm1fcYa+C4B/4ANGzDpZ3irZYczu4d8KjDfCqgBoK9IejaOa/2+6ZUrsYqTBiJ9MAtuuhO0z6gN7
p/NZBizFnVWREBdXSuC3k75zrJs0oYQpf6mE1D+dBHugnCJX6b6YeYsg01ZW42Y+zG0hf3WbRT6m
f4PssRQBSW1sufnvqXxsWd48IKj2M5iNr/DoO7sCdaOHuJAnYqevOnBwSlGMdc4lgsWpxHpP4c1D
d23w5sYBGN6JLPruHJTCtY4Dcpw7CIhSXjP95aVIr1LGrJCXk6TT7qdGOpZI8DwcmkBqeCzVa+Kr
Wx3gWkeZKfqJtymnHOJydzwlYTu/BdKa6k7bF64jvNVQjgM/RsUeLrKtrML508hWUUT2ilaPO3pP
8pMs/AHvMrDGqWUEn3/BZesXk7KgRFLf2OP1/yPsTrlVRCJwMKICmy0kl0bpm+R3hhTgvbychuu3
pqNsaF4rEkg218tKYgac3xaEPEqDuATy0jGDzmpjUuErC69xdkcl9dF5gLBCefXy3XDV+D8Z3nuu
JVSZY3+00GbSuXbYqSZoSCXJ3vyDZrTEJQaEMlJyXtNs0ygO4hjQYWcTQALX9E132r3lIKHWiJvd
OaHwr4zO8+qgx80uPVcgsDYflewJwQqTea+Oi4pyXPS0askJvNcdK1Qpq3zGeEwjSztpjd12S3Y2
pQu+9cDhj2le8TgHMtlNCa1J7bim2/iWelSeouX5MIXnHSlEp+jvkGgdLWhHuVIPwBZEfzMoYtnD
3W8n9+1fX/qmoTkBP7ws8H8XUIfZ0pm5ggj+v8rvOVC6gNDSGknZDPPv6CsIWKhLVtMDgKPqZ3Eh
/mgRwdw+mXFEOZYrojSkG1SRbZVVjY924MXlYUjHK0JDdTI4u90zaf8mPcahlKuQHGOL0YSNI/8p
uD0ISy5Ebb82E/iFZf8Ak0v0khv/wk01pZ+tppcrvWvGq3KzoJhKh6gqSqhzUq16EJj0f6LQwnwN
w0PjGMP3vsG/Ol84rhhQbPqV9yyq2oXtHniYIXYNXr/AMhJWtOYowy3NiaLn0WPvov/z76S1797A
/DSgKJqyb2mKJTN2SlkdsJ8EYCd62mCpMmEbLJbz4/T99TFwKodOMbPz5dkNjZNA3KKobonUVY39
/amvkUB0uhN059dnDHPsuL9eil0TKoE8gCFY1Ps5cD2VqQJWFNdgN9uL6prlYgUuLuZSYQ61jgMb
fx3bWT0cfujpx3gmZNyAsgIJr9KDuWxQMT9IzWCw3FYkYToFUAK/N05GSrMR5ABqTAvFh15pWqfo
y+4eJO1HB1XkbXrub5SBErbbhZtBqdUCg89LRSVOoxry0pYiVFn5X8S5aInn779SZQiLR2IqBb1D
gg3CYqfb9niuLzGdXpY3cyNmjTe/YuwCa78OrQIsg5jUkyNSAnd4Ccq8TQJdG8+8n52tQW7iRgIf
XTbRtA5OwT/Qx4NlSnyqH/Ng0ylzt/NA+DTX2qPoUzxY4m8fpGouPyUO1OTVb5pzUzISZOj7MDuN
6mu2ycWjcBuiRuBNLh1ncrwD+meW5/8JHIjc3ZPm+pY1d0FqWG1qxa+60hoKfsE8dX9VX1HChvk6
EjlYNrLz+vEqstsrdAjgukx5mxJYHkqO+XKPnXeL4gFHGfJuYoYRflDoVDMPxRe3284Jy4iHjUvS
bVbHhHdN8XMDSer2RspzKXlGx3tZCEWBY63Sk1jzpDIunXz72ObbZic7E9//akLMDGaBOUSImSgh
F9Q9TGiVV6MnYKY9VK4Vo8SmVOWyyjQPfAqeJ+O7gsvWMKbeAq9ItdLm+bovcU9gP/hEOeYS1GmE
a/pYu3+PjM2Zd1bQfA+ZMoh+2uQkUw/wxXxcT/1AjaqQYuLiAk4tsQ++O7FrzgB0I5RdClBHFqmT
4raU1/D/V1LC6Cyy+lnxIq7Skwe//sXzJwU7lV0jZQqkNtAnZ4cfZnMuuMQPd8OUE2OH/M9TatMA
UxKvW3s5LVwo2E0fARveEsWpQzbCd82OxIMgwnvIEqColll7GyiCsEUNq6M1j3IObpf8cr0iRiBV
TY4M6cgfLIC+losXHHcIKKhwIHVkFWAFCiPOcug9HukTDKKMkJTzy5fzgu9yR5QGrimsoP87Z/w/
ErhqcJ2f4maWI2Uz545FxgL0GddReY0Em2XCEiN6hRhu6R8t6imEYphJJ0h5K+aloPGgenrjWNVG
13OkmAXEMU8Do4hlmRKP1r75TKQswWtMExvpct4gHALMc/9fodxXql2hfwU/Sc05ASc2oZz2txFa
Wx3S+XJ2FJbCwaKL0gllGKVYXlu92RS29v8wcJzGf2XPb2QFD9ARRmYUCm1qlIlgwis3NodTYEPj
MT2RB8koydV4fKplP8/RA0cUPMQURDDVbCua8YMbjlDJOPGgsH4JmxXaLedpuUuOMPV57uwmvToK
H7Qec5VfW37pOusdtA+725pBuYvHCuOGz6VFs6Uh1bU6TLBkTg4MON8SV0Rh96b5A7HfMpWNM6++
Yd+x8Royq317zd280rsWkG8Pod4+SnHepjKDtfNdEB3YkgLF3voALfD33TcITKaaKtRusYHWtbUD
Ny4XIeUw1Vm3nR0LaR2xNmXRPuWb7/zbbqr3R2SLPMmxxF4c1tj6SA1z/wstbmjs60DRcRZCQi8L
cg9Ao/HAUB1oJhENTUApuKu8wVU+PY759uJb+GBgsaah8CiA3kLg0MejQkdrw7+kVU/7zoEdN9Od
sbM5JQuz/NQX/XOqMrMYDawstxii+jVFV1WDi5ASniFfW5kKe3iVQRR+hJMuLioqrHjJYXK8cFHT
yborRjms2SnxrbwhMBiHux2Mft16XL/ANCFFC06rqpcTJdGGWcxVxXOT/Vjd/DxnrU1wcilfKoP1
z8jkCXuVujVfbUTKTrWxGOFzlu4USDnp1/Oxul94vV2G4YIEPJJS/K3JimCHPXGjMYoRkv0BxnLN
o9m9axSgp1knCJf26xi4Nwwm0nyTKpWdbxy8nb3NX701Tcizm2c4nV19XOshqbb9TMIpt7gml8Ek
muwuFtBBuN/IF+XixVrt2RD46P89PDPQ3M/Hhp/Yn7yUDiv0NgViabU4GFPBM3Lodo9BY6zA44iA
GIbUPK1aT3YmhVclb87RJfnfWxKhuJp2zwwkve04cfRpAsKYbLSmfFva7axTaGtM0J1lXavMSG7R
jWpO9fZc/DYYO86gn4KOR1EtBNwsstZBtE6d0YdRSFPQhtCD1qrj04a5IGaz9pOXNlxNAo0cznYZ
/89pthXXwuDaBq6H0ugpbtxFsxP8yupn+6qnRiNEqvdqSXPzhOI5wlUHJJ+3VuzwKr54zRVh+O0W
6SOXdp1tCEeUcUyWWSs0arawj750hsMEEAOYWQq1NutnpwlpBYiVc2HMIl5/EGAA1JYXQoPjHwbO
JHBtqm+Z1VzEqGfKzMAi4YV1S2V7jG9jEVPkYr4dMWUSo8EbWFOm77xD32B3oKcpN3TCAxwPt2zZ
L5PKGOW9PPDNF7bBsnpYwaYheSZVUOQmpUodK+amHoBekjhS65VN92boHln9qNgz6FatrjVL1MOE
O5CY7zbWSjGox3TJl70omjyZxzi0LFQO8/KFVW+oaOd+xUIMsGeAY5wiwmkLGR2e/9W6vSZu4poq
E/37/Kc0yXtPi4JGOJ+/mEpTMv6hiS/tyu6fq+lDAZ4rmL1zj7CfyeJTJZ9NBn+pPEKIcxgEbCE2
y6VaFpYPPpt8wusehGJ9s3mfr+fJnGdex4B1kfqUjyPguqpLIU40hsUc2u0xTfqgLeUWdqfaQF7G
gn5m5GUdA/10WGYn4M+JIR6ItP/yhGiGRBzpUOFpJbmi9K7a0k5nHr6VOBjkinKvQUbRO5mgWdhO
YIp3tHfMuMA4mV0e0EeE9mBNZZrmff4DN/cmwLa+T4FubNEpqCZpEYw3nBSyJVxY5nQphvQcveAI
a38JwqVFl7m9FGqrmxmCKEUkTNMS93CWYL79LOkAJZL1d3+KCtLgbbd3jWjLNkYjPsCWAPjKlxhp
Iow3AmFkp8f0yFavIyTQhrmgxwVduBeMUoNdC/QRUYnGE98rmNCfLb7PBvs07F9reXwzmo2FQZZl
0XSZHtGINY2S3nzEeEFo9s/Fch3z544B2RKm/I0JofcmUSY+cWxDpglxyG/4NmtasJYqGnIiB72Y
40BRgWLKYJFPdyAcQLTmz5nFiDLZuqFl56t1bSCBAONrf3INUbNY4ngkjng8td+dfPJ4gbp8YfZz
bjy2QMpwSW94WEg0oZ3VncWQVCXhXoTn74vXp3Sl3IfOEDVCxNbV0Om4gmFhKTJrWY0yMyrZul28
ARFVVgMQO8JD3YN2zWVUGOtd499khIQQrt1xnKS8/MYR6apjxJjFqCPdWmwtmo9Q6oGxqS8XxZSs
vUKNtfKFpyKqOPS/eF7LH+nfHneWbj7BHA/P+6Mrm/pwzXUZctAGElQhu6YZkOA8XnbaR25DdhgX
DL0ZqBlBnCsU9rJw5txzqsuM7aX0+9suNzaSrnHpPPg0qVu4uEnExXT4EkFc/xA9O5dpbIzfWk9s
P9kLRXvH67HRMysOCQMshqhFItgjom06ezjeS73GDUA2+1psID8cr4wRotp8KrWgDflInkYPZ2Iy
u/ovBl/HE/v7gIa+wLepaLYf2k+ju5FG0Kfjb5kzyqUD38zlTfB65QiMXPpKM/9y8UDmR8QgSm2D
v3uI+61y69jLW1VHG3AiX/wX9SKfsp+aKSUHi0yDYRKPw+gJTBfdbaJHJYaBxRFXslN0yKoo96v6
AmHnGQ3LRvaarQ7sR2BTOv+Lgmkel1TOZM7Zzc7K5s1J0fyd+QMZ8ROtz6FKUa7owduhgenqawXl
9qsSaFyuKnTIS9DOluytESc3EQq5SgA+qv5Q7uIED2alfZjENt72G+oLyZAf+8/FBWtRc3CoH5JZ
6IooTtiiqL6+dVAXYrB8STxVAzTHylOXeLZhwatqYVx1zPXQJz5rJyV8saDQqfnd5WZNiscttMwB
PeCtkxXcP6b6AglKhgvxj9qRfkiaXlmjmLRBC4z6cg8zNqGSDUEmE+L2+KZHZ0e3mCXBEx02QQgx
47T1CTWjpZhR5/YZuSLya+YpmHnqTTZR74LXuy4fSeGISXP0Enkb6637ew4K9YM2Cj4v6GXlTLnD
WX3BunoiP4kubR2mMJRHIv0tSWihd2liTa4qlJEBIMkcHPWb/UNmw+KWep1Sjs9JEz3Q7Cqg9CAG
Z+Xu0qXDPyTK53TOv8MsWQm6kxCMTLtbl6Ndvdmx81w3HbYoJlE0Pkd+BGfiuF3t9NZXg1myvxVi
9KMjP5vWEIarBZRKY5Rkrs9qUxYGgkUyxSP3AQ3SptxEeqNXBWjRmOH4yRiNKf+2o5+WuiSVJTGn
vJ2Ay/h50YdweW6JxwQO8T/q9FCXuXuwVg1jYKNS3VBJA4yTAqlrB5xbP9ZWq1ze2PnrmeFvffsB
cHpsQK8BIzU745BxORXn2Pb+qC+7yxVzPZxAW+6rFagEUhqH+CJSJDsafwVj8UO4qNHbHoFlkKGk
iL8mrx7Tz3GdeNm8fW2EoHLiJwZ/zgBszbbYwdBB9bSY+/0NhiElGuiX9rS6yNfFaQGn1HAPjHBN
4cQxIkQbdEfJ6ed+/TA0VJIqPH0YwiB5afjz+0d9vaZReY+ekGIHltpMGFwGmhzqCrn3aDRSzr+t
IY8j66Y8Ug8IDlxyjiVVzfHlSNkUcsb4TbB8a4gbMJOdOh1d0P8R5Aks/S1l8fCoQPSBC+S6lMvk
UaGHt372s2SfVcaQvIRpNoYrYOdsJ5fCVZGdKUKYBcR7oZSpRJ5ntMRBexXVCzf0oJsMvx8Rw9pf
rTriH/MI0BaFXXQH37kG21m5dbhf83zWXPXNscNkPask/le3NbsckmjoHUkjktNfh+vc7rEihVlQ
oCAp/xuc11jtVwXDFfNhon6WtOh7yOLpxTdlJCdosdDvWDq/fHS3jP3BlBajEv/Gd3/Y6ta9/wv4
sS3BawQJVr05AOPqX3U+DM8A088D3sNx2d5s7me6+C+Znk58ejMmuwBxs1OaW/ALyuccfrEqYUaJ
yWqjNyetItYdeOhmw4dIe57T9kAg+OChLUSVK1FkiwLGSixbXvvI/S//RCa4MPsqVsBq/oYjZM3J
kKopa1tKy0z/QKGYRDFgG6MKoy21YaryJmeFIQJtGxEACKL7TqZWMg72JhDUmHQ8KxWVl0eWBtUw
NkneBOHCnBuEYIGwhQ8qRmV4uTkhl77EiDRLyn3arjdf5HVla1KVKvAvQRj3eqy9dqxJTuWbR/st
pT8W6/BoHzD3R6+cJ70sSt2pSuSKYsumsTZIOYpP8A4u2DY2NpNvQUex12XgV8yzaWnRHz//wsbb
XmTwZeNQNe1EWmiv7uGws+etOYS3nLwYfRwBtwdLBcHMx+Sg9XsLBGtxSIyZyhuZNBMelPi5X9eS
LTokrJL4BLBVUC2sL81ZILmKmKMAxJxuwxU31ItbLdhAS2WO8N70LGfcgKoNJC7tCSGc/i9nSpBw
5TNnfIlLU1qigdVFMRFuL6KhT4xHdJzvqocYpRwiOasN9dCVAfE8t5Q/piKS1PiyhoodgSQ5cA0N
3Ips54vveqyQ0wYOFhNvV/n5FDdvhPI9DsE092yecYZBqaI+sebleY7+mdeDdAF8sylzE3dCMnA7
p3rjW2HWzcNk1fw7jDARGAYhSSCVdafFOafHeiZK46YkYM19y/uw7KLE/7PdPHOus8asxxkLWpLG
mW0SUpFQnscmu96YE0ndqrxbJEkIuJE7UXHfevs/KjTQN8a7WFgOFXXxr0EUtcEzDqCl0UrRJxeI
X/678UPVJDAw13t8T4ji3TOyfT+bZhxhoCP9Fu2xf2Lu30V50mg9BfKlZeTYiLRW8EqmH4y0etoP
ayCE/doTZlszyKs7W0eYXhpCNorTnOz0K+w5ddTq8b8y8ReuxfNIOciDcHXi3/shKOVtFC9UmElK
BfZ06YyJKu/9YdLb0Y4WSsJsJkhWYkk1kwGME5yrwkAjtsR47ScbIh9twSEctoyzTwWKdJUqDJ8W
wZQoJ7Q7Hmr7fnpnUdcD1AfRzr0giOn1eDAdOS0yrizSHIT55aV2M4sbZyEPtNebKPB1jrNBvgJ0
eIwbxS1mEP/1vXFbFPU2tOwcz88bexZcvlOO4m26cK1w1U6XNyxmcZjCoe61sQXTbDrmDQ5VmozH
ruJ/qlc4KtwxsfuYn/AieAZ0QlNGvhjXAAuOdZ/oAZH97OKx7pt539Cxu2Ag5cwkkBAWauKOjDV/
HoDs40lQY0NFsCkha34IwYwCEm4nf3jJEJd0UQUkGas6S5wYSe6NmD+Duc7wG9AWCwmSETR40xoo
gRc7O+gkf+Hdf4lcBp6qa4jZz2DD2Tr+EMrmEqyQczevlHxnTIzf1ZCUDwCFz+pCm3OIwc9yiANb
5Cv7ZjCq6rlpflOSOt+Nc0c1N8G22fpR/hWcrraz4fgse1DLO3R/5Zhp1aPzEBPNtjGHRgdVesS0
QyLp8XmbwHu+9ZRFA69Gu/4aWk2+98GLSQK4oKaPrpMNSA6kMx2YE6KeJvpAevBGwuwMHrfgjMG5
yB1X9n5W8DWUjvsvP11+gbcWzgWJpxTLUFNl4gMunAfm+syK4XEdPGYWFW2Qjg4D2KXfvvUMatTt
9UwY8Ed1I5WHHPWFcmHhTCgYBanFFJjx8b8fgFTEQkCf4adzpkmT6o1cGn+Bje5yVtV/7/ACvoOl
SXnosCDb/pScQRarPFw8KKn0UbPDkdokOFpnNldS9bsJq3wSIW4aX0z7Cc+l5qmua9V6N/fIbdty
q2uUnTWrlskuPnCB8HxyDtPak8oMUPCSdx55da2EInVeHaw6BFol0r6O3Pe+0UFoFGPrvKXiyi3V
PS9qUZJ2Op+XGT7W9s9dsgG4H+Xx1Nu5nvANXegGNK64LmBwYCL7+zxm16t8JW/4XJCMUrFBRq57
5UEmC1pj+DzJqa02TUCBG4Jp7/4mv7VRjinoxl+aV2dLzICEuVX6uzxTt74oqHPX+s/3aKA+5CD+
+Bjsxj0ER+bE6ITgMOln/p7kzsMqbSapk44SpGlZFLtQRbMvVOrwwFwdS49rsg5NmzachnIo5U7A
GmU/Nd9/7CYpc7tISCRLiDcGx43rI/xCjOnEAW45XgVvD7V6q84WCo4PoBlPPXIIjl2rF74p8SrX
/2qaQC32Qmsdx/7z2S+M0PIckNUQlTKF3FGQU8AC46BN+djqWGzjSQ0162BQHuSMiHv6csIN0MlA
E59W1dF3yyVGOqA7vnfy2vvrKVnJ4HWuhokb5awzixxanSWGT/jX6z4QH4Nh6/smPtPgxp40LYkK
1xKUSUSlyVxJSTVeHKQ2y3FnqswQUOzk7+Z6n/IUlkBtnveaToXdH5MoMjGhp2O1ksbMS28X1KgK
SyxKX3zaSslhGI10edSH5EGFQemyvEO4Hqt/1olCqHKyeElz522LzaM9GMawuuOrFLhrmlJbrCQH
KqF7/H/g263QL88FiQ3vgoLmwdyoAXwiTCtz7iW1w0RncXKwaS0UY9iK2JJautbehvrVIMpeUAmO
f8aSGd9evkM4apntcmQOF1YSptaNXwxqo2HuLwiOVN5WvQ+VXlGsyqScyURjbjwyyQN3wKtl6iRF
NNKh/0TjXICm6greN0uVN6ruLWZqsTEK54oI/nJILGs9lvzO5yKKIB5lHBAovzcmdZtjHRxbYXyh
KzDYo5c5sGR1EJudhHRuRnLQEtTSfD+psZcEYofAxSCXcr+1nF9IEyjetN9Bhgg8+8aX+CVa+4ay
jT9lm/xfWPCc6E8E7VXQ1KRe4WaMe1mX63MDe0UIE/9oNYLoXUxeHEkq/W/vShCfSdBvl1ksSwWT
usZ7eraLD5Shw8UBjOAZwYQ3ojmLMAo418b3RTV3g8ZW7MJbuxZNCTN1Fq6PD5obE1I4K2v/bB/n
rw/YnqzIKt4MxBlFcUUi9CN6XM2MEkkXiz8VDTfznK/6OVCMBDF/bB3BOXgUWduZtjBTpwRfh75w
Ucro9QOPwUGURe26qDTCZmbpNx+kEou+bi0F/HmKtCRULxBXV522zLrRIHVcwXp0P8CQbbDfZYf0
45lVBzIe8J4BZhdPjIG7n3sOVha5NsFEEw434mm0L6FsaHZ2kJY7PryaE2UbvKpsKEoXvs5k4QpB
w8YkeibBvugU6t+ZntOUfW5zgIQN8XHsMl8kizPdrkxGtzaTFE0MLe/yU0UJQRPZm9CxN8w4z6hd
58RMiqfSw9/hZ75qyYAMLOBqn8PwIFg/NTdHma7EMUYXK4ImwpLAZRBs6Q/HLEEsyC38pOG9KO8i
FL5gZQKVZoTdrEg7Lkcoo4s/UdYVwB6MH/xfQlpxOSGAymzhnDoGoZgB9JjlSXsoGVKZezgNHJZM
xa+vQlHVGumhxq2rVDrYiQgTBHfkIufx9r24IQz02E7X+ynUA0A8r63JtgI0KaAFAmmCIDRSY44P
Dyd91G1pZEakeFyn3rDQlUY7hsPKF+DxO7iR3lS4sDR1XNTjT5eROhigyVLAzVGChztS1qy8cvgd
a3t2zylN1Y0Pe0fpLsFJMsJllWc24EnBecS1rGzIS/lpl6pfqK4OXdaxU97gmc+PQVzEF9iIY25S
aghwQV4sU1AqJLQdYOH1/BzqGlKgNo+XhTQ3hkreAep0GktFbkM94D+czEfoRwHQSW11A/tNlJTb
uGrSKW2XXBIUIiJ0Ft5q+wHL//pa/uJjfk+4x9U3zM8y4sNL1644pzi/Fts8ardfTCP2kxg7UopE
gnHmv5GC2uCmW3zaVHE+xK4t47tSWnYbHcpL/h7fe34GwgWptgeF7Mi6nCY6tkJ5CfZpvUCTznt2
eRUK/qivrYlb9PvKx3jDQMvO1y0AMD4vtBudtlvdH545kvLtU+MmWmU8MQzUvj/4kihDfwrfj56e
3YVESgv920lSPYvjMo4Wy2TxAopSAvPMedvMx+E5FUXBRL5zXEL+QMUqmzlbx/3b2xj2n027qTX2
HSOt9lvsQmbmNTvHeQsBseTfV5+XsLdX6BzMd4MCj0/z/asvyihqOwD8L/KqoC0oQwyZvxVUmuVX
cAfJZ6Bz/aTqFZoaFBVMkIMPceoyYYA4mW4l+s0aPMo8/HxtOssuIKCXD700CvRlPtO1vcI5+hRk
C8J/e00Sw1CVEkKn00IY8ToJI/m5i//7hgby1It95sc5tJACjp5PTzwyQsCirXxVu/UCRZ7zK+b3
EkOeA2qjN18ChQUX+z/CejZS+2LeTzbhEvuUUmLzxb/KI5QrxqK8IfmdO3X2wxKsfp62YRM1xrmB
vANRcg2eGhX1lCh08N3T7ps91vxTGdKAOZ2NbmEgox3nNj+++RDMU20xwkRkZd8J68bmQ1Jv9dZK
k9Npb9JF7C+Ggvo9EJxBkdu7HiR7mXUESxYmEr438GmiCRaisx+c4bi7+3qCsYTD2wFNPDMPdnyR
bWbo+9jxvWxKM2yLljrbWAxX2JGvwc2mGAGm+R4SgehQs1TbrJXOAYBQRuk1J2T/wb5DeVe3jvSl
L5c5iAXxWuRlk1hbNBhkpUrPgHtd5yFOfH7L37l29+jSypEnIXxHWMaHy4jHR/sfwrPQjVSIdpxu
Id/+lD2J3YethsMU3T/yqOsYgOYKanLRQPg+y95BoU7lXW+O9LsN0PWHhfLGT+ndrAFNZwIHnGdt
zvbIzKe4T43Bg0r8XeUm8s4MU8ExlW/v4UR5QVpCRUsG204j+dzz8t8bDLjSmEvcWjkfPz2sO6VQ
kBAkuFVpyeooIkP6B2Dyn/JFwqvzq2IWubtM0hqMOaapskuARI+D84GcIoEgbcfURWBCHcD2jJti
+azrpUEIDk/k2wifAnED9mpL00nYlb1BpvP4IxkAtsuhvuzkyNVf4WVvf5sBz0ctMbtPT/nzpEIo
JFSmdzrwxY0T4lOlY0+kSxQBNOzhp11nq4DewHSdmvrARn5MWVJlcOLSHTv/Le3dB+WMFMeM6STn
cjs4cxSs+8PqXlZwQpvWnF/1hIK51P0N69z8X0EBcWkTMpVZszRVki89hdVJDu4NovFu9eGf0AIF
3pgUW8lxHjjLtO9BuvXJkugwKJmTt+gTJ9SVhWfHnI5VVQzdPfKwTecyWWZdykS7uDYfVaxL2CI4
5FKxyK+HO79NVxobOGv/SB9yfga7AliSzFXsrlN9Xu4MsRIZu4g+fv7h3dcdGPjmj3jUw3J5Pc0N
h7PTcm6Yt8/coOlrjqIwLMG6PZjAy7MGDrXJXHfcpAvEIN4A15SLlQr5d7nmdvER/i+EckX3yoM7
67Q28XL726EboorIQpQEGCt4YYp8AiEuSHBeatqSt60foVuvi599i992d3dnfLjr1YEg3E1L7nR6
tAUXTrem+Mz0dThkDg4/l0SJ8JAFTdCL3PCEWalYPNo9bK2Z6ZX2qDJvAf4DEGWcd9i2eG6AXkM8
+0NjW459Uy7cOZmAASKp6elAwsUNgD8gl5aYN+d97r9B89W0gKlKYLwyoWyLxLnSf7iv9TMzJgp5
G+Aw657PzxOyLVeTc6fK5rbIXLQ2tT9hpt3SjrgmK/BfCBfb0RSHoEq5/0REsRDnDI5CFM0r4dzS
3KamiOjyxr5i75dZVJjbLtAza76N++tw6yzNes0cBaWSx8KrsE81gMfrWKV8nnBxyRBmvfhTpaG+
5hsxUqG5bAssW/LgbaQNsOQncowXN5eVh+nWrQ+hVM/Kaxe/EkTFjSA9MI6Z31Kj4+paZlrEm9i+
2L4tTHvZX4s3sHl2H5S3+1Xur8o6LrQi8TE0yLqskQb/g5cGdG9MH/f24X7ACs/opmNlN8S2nyLd
qIusJ56+tDauA76cR5DlzTmJUVNy7SduteSLMJ1FMVheMYU9fXsXY282y2omODR+9LQ9bBs+Vqu0
iA6x+IGn0i+3IscBHRSD9RiKeckx9bYKCO3MKJdNrsWBYmZ1XDryG/EON6qecrNl+r/l1/URWJBJ
+F4UYWDBYQ7fXAxhNjSuXYDipQcZTpF2lYEHp+lumWFybnY0upSm7hNbQV5h/et3Ii+1o391Cunt
RVZp5QEfvChYYaBsg52TDHqHmaeA04OmohwaN6V9RwUkoqQuCtoft53a6nE5mH3/iFukeg+DG/Gq
VltIzBd0BzDpw/3l+k2w2OO8fPqeq86GXQsq5tUfLWn9EimYq8JoRctILwVcNRf7GCFApViS5t/m
kWgm8HW+G2KWXSN7hBuTF/jIR9VgBdVMALWqDxPJzlWLS22kkWVlsxe7/uEprRBXshV6x/Q+JCCm
amca9GzwBZl6rNB3IUwQDZbpL+ZOPMyJvib4+1YoxLN6HejTl6nl0Hb6qDM6qX7dVA7Z9wuQcPZn
JgfW+qHmq77a9nhL65vhHENca5OL/n2p9cPtbxXX4IgYmGywh39oSNS9psntGhIL/HlnSp34ZLnI
XTkSb9o02Mi30RDis1BLFFORvaOLU2A8Iv0xvT18BeY/MevHFV26/kKcpp1Wmw2a4pkgnMHQ1WiC
yILUlvFp+c5No1mJ0apPHfE9uH9B4RCUWfMY/t3v0oxitXElIVq4K2u1en1cqvV8NmLhaUuaZxhM
7X/yWtsc17q2SFqSqtTBBLkO5rsuwtw0HL7U/qX2/PhWPBKghzXwK3Sc/GncCbiktoSzVKsrUrXK
ibnPhEzif7a8PZdDYyNr5nAsiZWP/LzTR1SUitg/l8ZdKRT9ddHR4xx7A/tuVWH32iyIeF8tqdi1
dnsigNluvpGFW9LC+swhzDnJ+18CEOleEUljkzyanPDDkGvXgxLvnhvTITlZidEn4VRQkD/NMCw5
otWXye7Hyk708MtOwjmHsOgd4MDPrOtgUwWoZ6dK7cqQ6BED81b3gxSgrYnwnimfKy64kxZeEJaa
bzag6OZ/8Sz7u9QXjMPwGlsYFu7mACBRyXeHLCeKPDy6Rw+aheHu4U6pNuyrnBdCldkTKUkRqptD
ucP54fhaJBGJCabml745GYmQCXUKz8SleK2CqGK5slX3pFOvTGH2elTeOQ2UpQ1emkwcJM8CjHmD
HSyW3bOcAEcI5gxFN5uuZLUB+9iOQI/15pXPeH60A1DM8eQU/ebMZKZEYaAiNE/d6lAwPrLVV7Tj
Eejy+KI6vUD4V173Td0PgqbEM0O05Wog/k0jG7KebwJNxeoCm2rroNCpqflh+6gBj5kCAodF/xEf
jNUM6MaI1k8DANwO53Pj30aD/FoRFRRJbYA7soKOl9v7FKBtmsAH5U0o6N4FEeVPLjI8HN+X+BQh
F+ztbBkVacF1AWoReCEgZlyqdnsymagzrmupxqeIvBZYVyQ2KY8wo3peyojef4m2zUbBkwCmVa16
SaAwk6niVWZ8XgaqZiD9B1q1WyTFBhzH89u9FGCrdCoz7ahqR90Z5Ez30k0wxZP3MkeTNCFkDEwv
rZC5Inn8Y4vvb2ba/Poo22l8DZ7kZMte8FSBSgPp/a2T2kN0wBcqq9NQvCrJ4yGRI+gup4vBeVMZ
Jgk+rmtOQvk0WxCjsTPCZITR+e538z0fo9xGVS0cXWfS3/R97uNUQMoQQ8WUPiAlpdGFL8DDjD3w
B6Wv1qYzt7hlwx/aRH7wffiFShAIn/6mlOc0HRWxRoKZVJkgls9Jdm2OcZst8vcu4nQJ5PSf6EUS
SqHnJASuJs/dWDrOb11QUHGpEAm/ndmv3aMhFnORva4cUgAPQDiApvGCwHECbB8BJX1y5WQskHB1
f5xYnoOw/fO2nS+ziZ93pV4FdTEFF2L1GCx9zLGRthVIiMN6qn1owkAEC+B9pyrEkAg5IgIK/0m6
6JZG/KppfgYMbAMXsh4BlyDhRe3DT6SoQ2z5vdIc+qlduvj87L9rig1EadLPyC9b6yPWVxuawM4R
uZLTvoXcASSeIVAOykxQDZa4nJKy88sonbDnzSNFWJ70THAjyxR1zFRlXuQBZGzKfiudEM1mmzob
/qHFTq9eMmvwHV+XKUWWGaWydypdQuHyVmGuvXSWKLE2j+VNyjMr60EotWOHAthWL2z6zTOkjb2l
8GhxA6PT4BjP3x+yCtGt69kH+ShsWGhZzvWfA5uNNh0xbNR8Cef+IrqxEgdLVYcAQ476Rc5LrPmF
s2Ysgau4iwPVeav92upAP08/PbHSLDGCAl+BS1aNrKZWwdOFqjvMsty+iDODpjz670jXCb6za33m
V29NGXhcqOVsm0IvuNF4NfBFXZHkxEqMk00+82QcBQGiXYhnyC+YYfV5ylQ2aihCF+T6OG2VFAZg
0k5Kjy3XSrRuACflDsvfmsAmQcPqwLCZYiFgZAsb0mRzRe335YYBQSPRbM5d021wS+pjx85FKCbb
odx3urw5V5LfqgQokKxBUxx4/iCEzVY4DiAy/+PrstR6zKRyHrYeSg/LQhOaNxEsmt2u952XW8tc
AfpKK8f560zvetgu0L3v2n9gyOrJ9t8qU5mMgYLw8XRT7IVw1X+pTyRm03Xs9qgxWsM4IvmxMHSB
e7AfITlrBE4fcuzUn+6HQAVqK8Otwr3uDeg4AXI08agMt3z53FsNmqUAy4QM9xyRHk7rPbOzZWy0
N+B2IUGVK7uF9it1tdPQ+Rx4i+TqgPRh0CKffmOnBkKykHpTFzA7pC23eA1x8xZH/WFlpWACWnox
pi9NnHrfcuP5Gx9DVomKXe5FtMyHPEbUCR3YYwFhJ0yM1oKyzFJrE7cT0EXvFSEaHWNDeJFM9Fb2
5aqj1Mtf0+QBvQtCkiyK6tmUFvlncSi4PKvgrSnJKxug8lMOOWhQb8ldq0B3t8Y0hLZO3yGcR0kh
1ZCkGXxdTqxrW2jY9FEb4I3PTxRR0kACeYzFzyAI9QopBuVlAVAat3r+Bkg/zC7MclF2Q9Gfsclh
55hRJ0RNZNK7BGzKVXILK/NjbRMSjCbxbZV4etcLwxrWW4nGLAixMhEqdYrrV0+8hUzc3+r8Vo/C
YXsR2Fi+kxFwV7i9vrJ0XlIdPrc2QigebbP+SvTdcRN+LtF34R8JcuLZuHTN5FexanGC6ToIEo3b
8YrM0nSPRWmn7TPw7zCg33XnlK2x3J79RVI9QoAGz0EBkxYjqvkHCxwisgZAdYL8RbPGPbLryJTu
ht+OUArQq2SJqseTyMrpTtTOHtihkxOU5sPaRs65FfPDyvqiVeA0vff/TD0rOOhweCxsQlanjdRT
lEIWvOK70JuDPFMDiF/cc6VkxIXW+79mwc/tsgMiJ/o0EExO9k0hLA5vArRId7/U32IiS/rniUKh
HuBwNRFZc1jrML/RF+HY6vIfAY0zyeAzMf2YuT5cAxoQyRSuFpGu8wGN/IABkTv0d7uRuMCczShR
mW7Ni6XvWMClBvmgEwSK2RjaaSNDgmGvBZ7BquCkDFMJh8c0balTaZZfR/Em98Y3Fm5z53nexgqu
QBQftXoUxZBv6rQ9uLC26KCPb2zkexnyoNrjKF1CIYWUBCHa3msXwV/4+LDxIZa/AB061LOnayx6
DLS3EIVrqlU4MPZp3DAb4GZI1j7gU6Wi6cQYg1yXJeqP6gkrBBOz0/G1RTYtjM9no4eTVXBYVo0v
SIt/xGO0B1lFCyxQnmB0FOa9NukWVDiNINVZZ9QeTncnofBon4HCmd60+c6ZGG1tWBNai1Inrh5M
d2fgPnBIbrbb6Vm/bMOCIhoA2DY/65NMTpydEkR4r5darkel4YdTV9lBYoWfZV+eQxhT8LXM0fi4
vGdaNa+NIoA61gtl2RvuD5oNmRfIugUSV7rMIGY/lgDVkt/zFyHxRigPURuPaz6QNLFjMhs3iB4k
A6/QNGscUFokEfn8NKwsYI7SRX+VH0lE7kpVRVDgmTDQ82uXcG4wH39PlWpWrbDX7cW6gA542vRL
m1tyaA0dqnAA4BK7ip6wq7E2BPpRIpICdMGYnvIuNpXBzAp8BknvDvIYXHWpjsibLKgEA1w/PAxd
bj/6LfgWEWLjASa/41oiiCVsU/K6MTE7PNMvHBnpteqkVBiKoTNh7TEI3YgGXyy8V0lo18ODeq/p
DGwyBtiMyq5yPy7l4kUKExCvN+ZLxsG8kPBdVNSh+YGdgJPLZS1COR7lKkAF08l2uusKbrzCgVEL
JwgrLURghpn4E5EOSsZdC69OMiI7kTBv8/kM3U0VnvUnqDj8fTM+fO0O9L7F1DFuzntR9IzvgSC6
OeValqAlOP/e1/rxMzs6NiAoFWTC6J8nUzFQcXeVZMqdT+e/KVgnukAkSLFVcfQ6VOli8BdmoaUN
5kP7R7ST45RtyOzbcZTXIufq1r8qrq3Ro2NZE/8CXjhnP/Th7OCQTyRmm5vnqVXZ779bJSKmuG8Q
gxI5qiTjRs/bQb84OiYriqhxQ4w6Ytaq8peLK6oQYZjGJdSHATrBQeMFxIrxgaT9CXF5t2taIk4Z
KRfr79ukEVtQCaYWyoGHqnMxIlezhiFUAwap7yue+jjtP0E1wi/tqgnLDmAQjcQaAGZjmcDaeRPM
0Th2dtF4T+bTX3DmCYWBDzyWxCbKyvDDv9MA8e1jf27UlA7KvND16dMASzfKaV6esOdUhEfD3Isw
B0EXsixLW9Ypf1GQybcwggSZ9M07Lsw2p1FG41iiZyFzgDF95bYzVDQx6t3T8oV63OGGnjHHlXR6
CZzHLzSM2Dg18T+DEmKcpeuD4ynSUyn30xXtQi/+wwi3qvqcPrPI52AfHOyjlX2OkvAOaegtHBbg
/UlqOY/DntU1xgXMBzoHgxMFQkqordKwZgtCz8MDeREFhizS3Ne2ox+nbanL31ISsjkReG0AJBTV
GtSZWqZrxTbq+O4F4pIzV4KblcyZPXvrVYIw3tbE4x255KbQwCfEvALVzCsMOsCq3+u1i63/Q7qu
yUdQlnuwBSmtM2tJbHGY0EXR3JUvvNzbbjl7Ka6Y41L/kD02TStmURiM8Lo3LGZhkkFtsJ1VFUiY
sII53EFoJVxi2APhqIotRChRldtYwo4EcPVA6Zi2FAdieE4zSnvOsG8c3r4WiBFuiAIQmZVRpdLm
1zakisY2tc77NSfkf68T7dCXpdQvqtY2Hy5q7QIbRlbPpGyTAx31S7JAzCMjty2JPNBh9fZqw5TO
SYZHC2QsepNzXPtnq+5QwFGau2jN+vhLj2EiehEeopUFYUDE6wOKLFRdqPCUhjy4gQG9vgFoIApk
itnSOaXN1rz0V1gaCKnGJqejQK28Mipv2/kmQU52UUG4PdpnUHA0rC5AMx+4zrFRXR3Y64JYoYOH
5UKZyo9n7nI0kuVPzZAyseNZMjUY4cUjhoBQ8Fq2m6lzbXPyOKqz+0PHPS8K+UuQYtWJ13pPXrc3
QIPBeA8wU6WhdMaRDVPTpHCvVMCL0MJrL++K0ACXwAkWTFJlUcfaW1TuGzBJH/Ed/MSNmq6kztuO
p5iBgHi8wTsikzpN1DEa6cQ0BHsK/HDxxA4rgtXeCRvmDArkF/0HfTopWwOS30JmuK/C+iqkBglT
4C97wUgiwTmUsrV1ZeWanxi60SmKzZXv5vxPED9ontUw1CQzDvMaxTdEkG95jAW0qK2i2fMXF5nH
4YBBXJe/OBVrMk6rzJMZTS6rRC6h/v3HvWiItaRYDxfOk2r+2aYdL7U1x7/EZZ32qtx9bckCWk/P
BGhdg2We6Yls3EmSQBbL1EyAdrS3u/nXoqS19FN01TMdbjCcv4hmz9tg8PD2xnbzp1jLqGHdI9My
WD1z2D/rEmR7pheKvKP/TejbFTbMqp4EV8/ZKrehtE5/V5FoOmHWrJACB10SgtV5Ukl6xYUmV3WE
I1oEK8YtMAWZ6e1gdvjd2Qtg15HsPIrw2dw8vUOWQ5u6JtYGRjmjH/cVtFgBvjMTSbqOvyYVK5Et
IAPfY6A34bKTqOt6D7Zn7zXtClBrWxREVQQxRp0yuh7gFKQHxC/OUhjPfuxI6wOBOjwBy5nmQTsk
YNB2HWogCAQj2e1fABk4LVfFDFkZ2ncXpbgnuhbWj1l9vNjgg6n5TE8pcBB87yj35d+LQZL0Q7Xp
GUvOeWaELzUGxge2MA0BKXnMblwfqdVO0bD/8D8R/qPFiKofLfLR/SpyIC3CWKoq3ddCtB4HxjrB
iYeZ8l81X50Ewqks+XvFRqtPSMLURQENy5ilr8GTwxpB2cbeWZXtuCY2ldVAwCuB/utLksCo0oKD
8MwtrPzAYuSBaJIoqRt8kHFOB5DnNci7nDG6a2jrik7Kl02V8bXlmXml387hLYtCbP50OqHlOV24
Nynic40WXqtRAfMYx4m9CUTWVWE3CRQA0Wid3TChjja9K8kMCNVX75IT81WppE5rIgq4uMvYlxcM
kyvb/4O0BEJXGvPnhRj0FGi4s8NhUcSEvEJ9LmYJ7ZRux7w41d2/9y7cNcH1b0mUZ7cEk5fVrmaz
cT6Je8qoF6DdV8w1Xm1dqbh7BpEXmJI7NefG9ApjAr1CnGE6Qv1br+C3+txI1k1Ja3KWiIAkA3ic
7HjA8TURjgZT6F8lgRCrfR5hY+iTaTTOlK59Vqsia768LaCMWM6TINdlTyiHa+nYGj7EJeFmOiio
dloL6KQZaNAQrVss6D474JeKjEh4VtWkjPMNiq0TYfzB/vThyke7fF2CBG/7gueoLslIsmKt2CYn
hJUOJEMpHmZZD7ZGJj45TYy9WQRX4VKOtNccLYSXkSR/x+wqKyvmH2nWNf98eJs6jXqCmvyGuFLw
WEm+9RApZZTfTgNhv9ROnqu59VayO6coHifNH8Jx8TwSfrXbDsgY/gNwomEgoOLGeVh4xE104W37
5puaxnKMDEkoAaRJRvjtoUYGlEt4ockievqnMk9zZpOXZZvho4Nj/34hyZYN8gGaiTq2lrnycrDE
l5BVI9s3V8KwxW5gAF7Um+bNH9GLrkU/93FS8j1mx0E77yjnne+MxJsy7k1Fg5Rzxhd28UY8hAa1
w8wMkwtMYAh/AetMmG5TgaR3SP/5jA/U3CwsbSKIldGDAt08hPv4xzO23biaKNSyMdTal9U9k26P
yqsnz2BQ620ts6vT/KpQ+/ULEgwAA4u3H+vjMt1LdPcwW3mI7iOB2X0kjmCc8nKNrsKjuHqRBOdh
BJ/c4WmXxbbFWMCXEiAfnQH3h8irM9j0dbz/twIeM18UCo1/mBxgGT0Ud+XEMxrsVKAC7Y9Bl5dL
ew0O/rbYPKJbmfKi7lO3oO4Hw44ECpTmd3YbvTdGIrwjc/46kVnmEROMae/VyiJVxCJs+WlXKd4f
nsYQN+FSIT/cjovEm5iLsE0O1zcc1C0VdBaCmAr7urnGQVpp9aFGDjS2vv0yxWRN4vUEAoIT7IBB
OM+nz7xGCfgVZuAjEmsTJ85WWlsU3PFxdD7V2uWgGCo8u56wzTKiqs2SqwAqA+lFzZfDnl2xUvct
MQgRNiG8YTe5XylqYKWN97A/hXGxR3s6/f9jDt8h8fRxUMSI6G1KRTakA5SnKUN85IDQukTL8oup
04/7fg7bTe/wP7JY+XEUmkTrRPpfh4BqoH3MB/9aDoKQ5oNRy58h/eQjC7+fcoP+Uw9ACVOpl68m
AAcmZ2nB0RjvvIubWaF2SgawJKFl9jqIJMVzT7Fus0NbUUNsFBJ1acaD2w7N2EO5FzgN57um0dxr
lFzVWyoCjQcZnD1eTd+j1Cqfsxwfzwi41PAchAFzei6WLBQx7ETiEuyxvgqAXqn+lup/U5YE7SjX
f8OZwRq51TMtgoHUqemobkG0oSpUUI2pRgwrW3JVa8DkHmJhqXK1af1dxEame4wh9h3lq7+Xy66M
p1fDF/MzeGOUTwkvFAsyjMKtGo/kQ6qv0LllV99PGGziHL/jgDRLW9Qh0wpH9GQqgI8N19xPgRyH
QzloyZX4+m6Wqwpm8g87w3MWCj+9s+dcAON5suno28dtETICX5PILIaJt4XZm7IioW19AsPFljNk
9rsuDsOSb8mNR5Gb6HtdiU0FHxHyKmZTZoQ4u2x1jsrwDMPoDL3mcmfLv14aatnhiEK1cZBZ+15L
LzW6VlxcufG5ItBNv8NKU12J/B/ZzRC3k1WIkVx4VfiMDmACprCjGkktZbBudGzA9TrGA6eFFkez
S4oZ41jhazeKzcbaS3VCNpbKy6pKvl8Fpb9SIVYl/lrYJqLFgTkwpdRG0XpdZ/bRAOimoMNT1fAh
s9cJakTxXmwGqL63ZP17dqZkOVYDEAzZiZSCr7AWexY8/FVxGw/xnl+amxNJDyxFOQNfwfXsbwSy
xuAVdyZ0s1DM7XUvOMN3dhxTbKoO5jLAHJIzE5pEfJyhH2AntY6jeL3vGSaODZLADLJzAUBQk5z3
6McH90AZO2YdD2N+EGeqps4DpQFLYHslezYq+TqGFN9s3MHOPGKwTIt/eJdPyZa4qZAbSI9hBUjM
yC3A/ox5kdO4qcT/qKtehSUbKJ3Q61KSyY03rKqzV1A3IGgaXsORfk3a02jQsUJKwROcjY1N5yrd
hMLuUAWf16oFNxvSBd77XgNK2tTqxho/ZEppd/FtG/8HmKep5VWi76N8XJySEk9IJQT1wGSiT0Ph
XpKFh1pDachbaw+drUhLK51tWoXHFo+DnVwYazB51I2S3sqEGP187EF4tcKo+/VC7Q3je/ATbUKm
+7tnxbx4JHhJtMscAkggF0l0p8krE+APBI9tc68zdQbfJThjQZJeWYrjzeRDU51C3qYQr/j8U4uS
R8hU+z7/p30QcmzS+bQKV+7/S2tbA5kBki9RY3YvymopBgB2E0UaPi1IK0HkKDncmoa0d5rj5RLI
UZJMeXEXZZwcRUBT7NzqI07b3HloqmnInn93Vyr5ZYUpci6dMIPl/MROVWdzaehRjVLFn6vcYhIh
INMO2DLXk+JCb9KwjQwpWmoVauwfP6jLa4lWzHeeSDOhk3amf83a7T/ZLndDuaDks+eyUc+iyCuQ
pfo1cGAr9H3T8lnS7DJItPHrV6uJQF0UuvzXb97/3l0W+OX15ubaTChZ5s657SAvSANtr4JfZ2Nd
rE6ltRq6XZBwhv1TS/mGehZ2nbOhvO/lHVR5wFCUM1pmbqyHLbk2Y4B+qKAIXKFkD3pyLSDKUPNb
hfF5zcSe8Mqay22TWjz9musZIW5rVK3epP/iprAj33FKyaF/kamPV+uccqFJJyINFh8RRRwgv/Lv
oImpPmCXTojJ2r+nkPeXRHK+z8FK15UxlmhPqkAHT8QBlCI5AIW+nlVxcfIVXp/1S285bwHwzDHJ
qo1fYBY+9vx4EulMh8QaE23HK9k1Lnh74JGUew9gqypKF6Uk5CJviVWBJR0Z3j/61+em7Xw0sx36
8fGZGwzsxjxctEDcUTaiAxuxpR8lPdEKZF5keIAjHhzfOY+CggGYimoO3R8QHBAatyDFyDsWF4aQ
eEIn1P03Nl//6032T5TluCgV/zxfdu2Hi02KsPy0/5NAPkfVK6KctYSOjBqs9zFF9NbwZg4jRvMd
eOFAc3m+MCM7/PgwvGSxbHEmaqyHxyG/N3PWHiq5Zr2/n1EIw7kOGkrVJlpNnT5zyLzBsQQTo0+A
85JYqtT4/Tr3fcvYkylyDhXT0pAepeS+n5JzvwAp5zZqgTUZuzI+TQ/Xwu3KbQSb65K+Z1caibbf
QElKvtkpW3uv8FidJu3YtNGKi5DAdR4BLMyqU7mQ7l127A++M6U2ZczlsyU7qVAWvqbhIyDpPC6s
lG5rQQadnhjqR/bQkvWKAVbeKokV8jHTr5GuKGzdvj9bgVOd14cVD+7rRWePhoPOJZ6Y6D8BD1Jw
GL1LejvRSfg4Yi5V6tHaVK/gXGWAzGeVIDXfetG20h7FklnRUS54Y6zkyd8RH9V5+rkosV5fPo86
fOJaHc8KeRS8w5B8xWXB5eg1sXdahM5u/FCYgjYtcFnGIY+hzWxjZJjSkmIIinTboC/Q7ZByCTmM
OMLj+kRqWTfGtZtlxJmYfj2zRXTy8tpL+Rn7pZFxrh1/zgTyaukiUDKox+3t7o1E84TBOvn3et/X
lUooDJpPjvoHV8SldzA4ojqTusrDd7In0g0/Ga7P5ZsMIM23cLJqPW7xeJjlDuKi/CMQVwOtErD5
zY9E2jS+TK3zyCtTkvuu+488w85mc5z/JmkHNkEX0Ni3fYSxb/jcMlAIY6m6DRAq0JaN9DbRkgWD
XZiweOM55YJExgn2NCB7d7v3Np1LdqplvDSs8Lx+bT8q+n6ihOmEd2QeIhfACiQeKNgHITvbb8fR
AhtA5u2qXeFDWZaFjSFqSN4mOOQnhdRLS5saaj8A6kOEkfQ++3/TACO+wKgQ9m9dq+d45AOGkR51
CTcStiV8yZNSrDzJW4IuaG8Y44zBAE75qVnlFEXVM3QWnCgRTCp13AmfzNGyp0WaXvBzIGssUOZA
jNJN0hmvB+eJp9wn4AKh39+tFYD+XvyBvOPgsbOXWwBUarWHQPZai7wHBioJiAPyy+prCEu146I2
Tgwgse7bqbmKP/PNxFDpYshPFIkkzaNSQcad5KRGxKvuVZo13MfSlLKeVXK26N2o6Jv9n4m+trRX
YIC4sVI7pBZVxx7tKmh5os0qC+hGBUyXtIezeZqiHd4MH+khFkLTrvfBjM5HYSf9ITfchNbmgn+l
YoeUxeTQM6c3GLKsyETMIfd0KHVKh60xKwT+7dDkEb5l2mmyNExTldePGNyr4V+QoSxNqfna+y5/
2tk/6AB0c41hEbMDD55koqRNf6xgx41mo3m3g9bYLvg0ILXysrF9RIGI9xK4kiigXGLBfh30T+vF
pc2YBk7W6tFiOuyNSio+gA3ycv8/WNQSGA6nA7qsIMqIioM+8ra1WKJtN2PI7u/T94wqRiHysSXR
LHaog2ZeseHGlB0z+SZPekKWTHKaI0TbC0RpVN3Ro8dsCcFVeoxmW5qp8nkPcbPlObkjm3PW3Jpu
LbcyW4r2a0y7c2RyFWcfdImpua2FhLuWGj/pS62Z7CNMs9mcZy5b8RH2M90J+OA0RkqzUmX4PCV1
qvq+sfwhFul/AYcfCO7YZzU8ahLm38sgezAo8ihFEhoYz4YNU5rQC9cOoOTCCYM16CKvgUzUJ6sM
3o+gWHD4VaPccA7ExDJ9bqH9TLsqKM4NBluRKTXoWKp82EvU6cB/q9mRoLqDVJ2oLlTePN4tsqLB
hu9m3AY5WUsECFqWS0Gld2mkRH6KU8zYSnpjVqm5fMTIuejRCJQQkGPqk9aePGi5jrp7dqGbaRye
wElZ7JSzuOZ0LextJzo+kWZg53bgR3gUmbavtz/zexPPO2+FfFHW8nKFsPKerhHwwuT07OxYH76B
BOjS3u7ncJTD5ScvHymcEmXIMGUfEFRRqOvWv+Sp3WJuhDp3sKA30q25r8TBbAS0cMLrCObkelM8
Zco4jduO+Ftob4q7rrQWKoKVfVU2ZRASQp+skDxdKe0fzmdlhMy7gER0Dee58eJ3pd2cySTKcy1P
YiKIRGq9D8/swjm3hjfL8dhdANRG/D138Fx/DhlGcthVgzYmvcWSvst1J7Xf4hpeeUgNsQEGiOCz
TkhYBNU+97EVepp7Rq4oNrsOobBDP2Gzdiu9QMminKJhtD2pLTwIp3EcwtfRWwgTt7/+bEhNVgS5
TG9ps2ZYqtNfSxwjC+dM/Wh+bQy9pj6pq5fotOIHCitt+UlmmXREVBbdp8I4l6rGY14928vJuWdp
0v7ykkdzkpltUmYpKd8zZJJYB1QxFJahyOUse2ibxgtlpbljF/cB2uDYhTH6YBV6qvD8L87IU/hs
GVbAaqeqo9k+OiqOvfpNePiUdhfU9uDZOApBp2NqQXtHhsEoPXhv2+OyOyDgbIxpz7nWv0NtgvxZ
qRtHUGFHUR5HmW7Hai2MYfSWmdItJ4bx4YuIyg0Ha1kC/TQoZjPwCzFcpkxgRZXj4TjZObkEzbt8
kjl7ma5LOxNAFi+A/cXkZIWXoXmYcMu24/MqyyPkOz7wwyldIBHtohRHH5fPXEx5Cww2qMvFY5JJ
HZ02EF6zfAq1naJ8ZAQPdwoekpt/jUu9sK7On0QtdqiOk5wU5Pi3c7d3yR1QXIc2IdQV5Ft+a1ke
V22yzDt4AkEewQMOwzXqgdVqt/InP/hP/XbUx5jfbcf0ZHL2fgmSVTitUKSaFEtf+fWGX6T8W1ys
lo55ZDJ5UkO2LEU3io7xcEzhDrfrvQszoRfgYcmeOsnIgK7qoiBNBaalIvu7mrGh+h/BS6btVMTc
Q3GIjP0jHLH++wwypUHC/tL69pxQrmVpuEFKLCUhXWLivTgmsgcNHSvP3Ri0uV3RzcGu2BKLltk4
GJfl1MZDtCO0H9Jqhw2mFPERRJDjB1EpaRstYesfp14KG/w5MNmtwOrAqvoPZho3Y7zSRCutut8m
8B7UkxLFqr7twOlX/5JR5xENjkYUomAUPBTlv9CB9uZpiszyZt58Ts+tp6hLatDXuVIF8gTIF0PL
HK3yoylcXr5D2KQE9sVv1odzDJxOlBfeyGLFulobQM2wcaAK7MaBMOMoi85v684FHLomXcPaFTxy
cKf3p93plT3B5MxG/6GZ3QQjqHbddBFrRc9plRny77iDxLs0jPEn/ME0R9M7JrUM40bOiPE9ON2C
n5NHnBBqMklQXW4UFmq/E/YFxwboNlaOGc2x0hJdRFD1SaX7yMvmTOouwYAD35AGWL0cg3Yz/xr8
eklPY6qEYS/ehXT2sbSijsN7LDBV2gVQlYXFlxcpFvhkz4pdEplZDYa2widgTk3HEIv5AlcYccp5
mNS1KFsQZ8Ry7u+xU/VK+4ivX9bA1sIjGVaC9RfJzgduMphBM9j/eXytos27ZgVNKLrEqMeHRjBS
s7H4IFY8wD2X1dQRJL72D49nvwnJnlRGdkTp4E6A5++7bC5UTnz0nh8IN+ywxZ6ZxIgdO88bQeHd
xVvbkzwkNQiK2mkeSPA0gc5g7+cveTL9O7k2Q8Xk6WWIWJ8CMwRfb9lN849lQ7yn4CW5F0oUgwyK
TZ8XsFNV8Na1UJNRaJeTtUKLxbA8iL1N52MakYdRB61zD57S6AJibjwi4BFf2a96fc0UnUaDn4Qx
r3Q+8iWc2ieJMxV8wRN7a3XuHmdntYxrqZDA1acaBToDr/BceZF3cF5Bi41S8zi6FjSHVfoedS9A
DKAwcaHynEtE1cUuLTlJGj+OdgJWWLhvdAnWq6Tq0uUHQ8oRf9iATLxe48q5VFOm87ZJVvupPjfO
1oaGO9Hj0TLFQrudOX053YScDfL0A/LllD37gARx8HU0yvRXI4TYFb6/5NA4dhsxTvmVwRaKInP0
7qwzGZIJI4MpdIC8SZcU/lVIBEF85NyBRJgwS7fkwCicQ98NeSnnnl0d7vxAHaabC5J4Hhzm7qNx
JHPH2XbKP0hsvOSrw5xxi7lKH27PSc4yel8a34eD9zi0WrF1Z3fzWwFCqIuSeidjrLHFmr2Dd3Q1
33rOLR2DuPto7epEpHMddyYWPPVRoIdNFmcYJKOkDZ1tirnRx/jBgxoNb94AZlmnPq34ZTTCMH70
hvMI2csZ53lWVrm06fjhmqVZnfmeOJf984ygg2berDGPgmnl/oKo9hxy0ED47wkXGwwcrp3jRnWT
3IgncFVkj5uURnCa44p00TG9ya2/BcP7cXbSctd6+oqkmhu7gQXm7kCfiShDJ3miFoLv0VGSmMzH
DVUJ9j/7xe+PBDpOjsWAjCbmHP/JNngR8fp94SuwSca0O+Gi4uye2XswJT41/SoQ/ANnyXyOiL+J
k1NQlxGtVqPy02cmYd63Mi7De9s2jLx0hfr680TPFZwby7iTGBDiGJwuV5Y+aRHHtoBvTWf0NwZe
+tg2jFqP9HsmlepSgRcSt32NZgrpIz520eYVSHLLP2npCJZcpMVkeUCUepcRv9rZFYFqRbjLvWDp
oRA1iSxbiOyHACwcGNVzCBnuKxy8WrPJd32dlfGOm1dSVy6efttxJ+NvDoB33isvl/fLP5qYuh1G
muMVte6EDDPVBkOyT8CgUpgs6NZlg7P+6tjQDkZ/uUAPnhuHSq9pgVfGMWd+4eIWg0ln7AH18qPu
HvErFL3iKWVhFKYtgDrKMYtoCb3p8TAOYDyXIUAXEeLvvsYTwcxFfpGuuhkLmKBqt7d8HZ61H+V7
CI9J7K0yAKLQolXQgojo6rOL//LJoOrHvxDdn5WfgqTyTWoJPKK1f6l2J2nzjvCSq9ZBm1mu8U/Y
nQyReXw311FBK1zxEv+1fhUPKtgSUhNeZuq2pmBrACbT7NZNpXhhzMQW65IWq0vjOU7q+0BFDOGP
USM+7uWP2eBEF66o9CwqGPCC0/V0kz166gA75kebmqLisHjr38Kv13OE2B4b7lreTVay8GmLkMD6
RqYyePXaHqRqD7ulDB39DXyC4jcicUcT652pHDd/m7nIA4tsvwPB7Y1ZBxYOVa3U89l4tt7vv0vF
Nucudxg7TB0vVYi7isfzPC1LzAgYQprrm4rZQyGnbAHzVmsP06dlJpuEN6aRmhGC+mbpwvymlTV1
eaY94DQNPHr55/+qhHLKznEgNVOGxYE+86tkU9lK8hoz1iiMVg5UDA21eRH1EmPfR3UHljiZAv6c
H10HW0NWgJdZYqOHcRD5fcJBFaxNr/Wl+cRk8hkr7SINbsslyNODSlcvBquNtKKZHm2X9KVyDcqU
QB0itgp12Ti31C324+e0CXveNQcoKtYq3tz5t+nkBWrSrfgjXWCXfXqhcePtHgy8k03U+obExga9
sdc2xfFA16chiSk6snzilS74qrjLBS0AkBK3Hn12GKhN06DoZi+oLVEjxlI+GHHm3JUYWe3fz0NJ
QgZdLReFPNli++i4CMohlrk12WIv9ZFMl9Fy+EFQK6V1ENeXa2OSQl6bWMXG7YokdSEoF+V9g8Vg
Ei63HV1VFivIyKRwH6cmM5ezCgIuNkiakSjP3L2ykDPXbaPemrdUcXOgnjI6IVYBnM+7Tkf4VT20
gTfHVcfUsdGbjIz5cmSghjDN1tf3UvlVvuIiYmkHaT7zGXGzWJsyO8IJnHdIjbDuV8ZCscIlkx7+
T5k/w+pYJkrpOK7Up0CPh3yCGzAc0aZLOUDaSx60TFwxZIt3D+6aP7C7GpcY3ve6qX5DFSV724sx
6hcXYI13EkPNVD0JhDRS/j3ZXZSEYkx5CxN7xpSrQyJFloDQlF3tgyuxLWI2Q5d/wRBHf5fBV97G
Rmyo9qxrDsmeHGXIx8lF6lk6DKnZuCE4tjGTCQq/+tjyeKDCp1gFrUuGxYdO8WrttJOT+Oo93UUw
ISbk12/MTdWeCT9cWMlV2Pz/kygEWJN/MSaSIhw5VTI4wf407m66KpuFXOz20jMA261pYO+Qhgvk
eaUrKzjH+D6/8K67TEJBHiYhRZafc5tjjGbveS4qaW/nVJdb1FcVb7JkAEksCqUucd5HODELhmsi
7jBknTmyd7Z+lzZ9PAG5T9pKIheEQn5lKmD5zfid/+j8W7IywemGlNrxPpb3EvfR+DHdgmG76MxC
LiPQcrTYVZM/s8ezyLlOlTvRVcwSz5hmAXtpQg7ESygu8CHvn30gIvWhtYemsuSsensFinXp8Wxg
YFnJzBGkiM/Pl4txZNCz1ZpoeYkiVZEpGvLJf/yQjn1BBvx7hCfJFU5wxoF08iRMwE8K9RDv0aZP
AGq6zvcgsgHk3Ax04SYOQ6TJXkCQP5uhxuKTM6yNfTJQCUm4Mpb3dz3gSAy2yJSGgmsuWoq878rq
TdNLR5rcLkLWU1qGz0TFtKN02NyYwaTSPvDqdL9tBA9Xgnwvn1ugRXYsAgmNc2llyvJ9DsrqFF72
cTPk+sgI1muVbmpvhJp5NFE/IoxQgYKbRWSv/bsgqEmbM3p8s+oQWw6WgX8aB/sCS+IeQiw65VpR
TzHKfmI2E9J2mWQr3fcDH4Iq9ZNw6BKjhYj5MMwHKTyWiQX0By7rCF9zJj0VjDJMyfB0LwQrFey2
1vLjdrUHY3Je6JG4mUid0r6yMJ2R10xHoUT3Up5oaCXH+1tf0PC9HC+GUDPlIGu7E1bsS7Aml2iQ
JsLZJTWEWPWwJX9lcykDIsfIN5zTUVVAjcpPQfG0ibaUcZ4PzM3kBRjBFUFHDqMgHQkpQ1LP0Z+j
iLCorGfKUlT12Dpf5WrP58+3YLrEljn8NLFUaDokQAJ1eHHS44nP5Z2f1CuV1Ii6rDoInOZZjHzy
3QmQGPmsPk1RjZN2iqA/EkTMxzImPfuZA10lrvrl1JU98Ae9M1C59I55eG5rdlkXF34x5RQXH56u
kZpxFRmT75KpPiObViZhEhEQ7TZ7Ox2nRbXRrz+vGrHkIAQloVIIPl9rCbWLyEg9RbjmP6WB92Z2
kGw9xLRSCPO3wR57tcCLvfs6rFA/SOgcJhLBYj0U7o100rHkAT+jlkJVc4peXioN371u2jTWGuqv
h7YHQdEjoN/kpQkG/W1JQFibuMLp0KPczSfea81zeSUjep83DhEBHZYTDWg8xbfefk3AyInYq1KZ
7ucsYi3Fb3LF/5LbyFtHfAuCBmrJFERp/Lz2V3rY0TawD0POvWAh6/7+K1ecoq0KSBIhhseRN5GZ
JbQhmSWB4epFHvlzsacxY9toBvT6x/ijId/tPuivdf1Cid+uh87QCCqxqqArWhKkG/V9egSQ7fYm
p5yMqBcqNU9+EIBaKdfHlVnB5j0I97SEBEVOQDWLOAFvpsOWlIOaotmSfG9vlKC1otjXbSddoKi5
IljAwIIglKoKskB+HP+LJmq2kSEH7iCaFtdEARgzR7ViXJfCx6bzacerXpwQb2v5JBH7M+GKpvP2
XAsTVCpNlZnrPyFzRGt7pNm90kYlA1R9dXa3W9V+yc2ZkGnT4fhd6LpIfndITItPU+7O4Gg4rxCK
NJ8YicMY/uHMc23TV9svesPWTC4sZCY3JoNKu5/4QkeaF4cS6+Ed8v0568dFTCtBchzBUZNsRof3
/JdS6c2roUdK08qbjbYnsjbPGjR7o7uFtra7J3j5yGic6a9JD5rjZv4yRJr3TJlI31Iq0BqV/IZQ
sfp1LpX7jJsL51UYE7cB7sijrd01vIiHlBgDD0X6nBI379k8CfHN3LtBP+qEztR8gBDUT+fnXqHT
6uMBijD6yekZjdkMMlP0BPRH/hsoGda16PNjpcnMBSd/13oZH66xSmaMkItQI/0cFDn/pje5Ro7r
GGHjBhx26XDGpXQWBw11IpxN4pwPy8PqqV6au1Hxrs3+7OfahfNPTSXv0qy1hxO4yPyDUDbg4H8a
Mogdv7DJGfC1l3ohNh3sFgevUPGo+dyGJnLXD+mUXVxKb35J2Lyg9aDpXkyqCO2eqmQtLB+PqBqx
Y6r7o+717hwwf0JIHzMJvfbo5FvfOsNJ0uCyy4539eVJWE6dKV1VunXOHwskstpj/sVec3pbHKac
dHyiUsKLegKvw2wy/FSWo87W+vlbGf4Ka7YMCMabrZF7HKg/pWz9h1DbD9Xd04xLRNnCJL5MkL/a
JP2Zrz70N/fY3r8nFx+6HSimAr2RXjocbqra4poLNtW966NcCk3rXBjPudhbTloejczAknlZf6TE
gQuUFg5lcJAiLeSNT/QGcEQ+NYyPPlfJPsCkZTEtII+k6Q9jMbJWOk+BTCYicZ7/dbDQbWDkSt31
xJaAGKTreeNooNnPVHfBcCmn8rz9oZblAxZQVq/fBL0/+h1Aud8ecf3wbfGapZDzT+7h336rhDTF
2wTGz64EJWgYmyH4sTvvy9/ccN2Cut2mbRBjHirVPIhq9FD2vTqt6DcR2CLLN3qkcstgn0Qnrs2q
2LxFmEVahg6PzCmjP42c4tz5KZ+uF8XWpZEpYJL84ZzjaeY2fvXixD/NfeG9BpI2bqChKODaXRg7
niTcWuTvG+0aELoU280B5q8QoPZ2wziZ1jWcJgaSOt+lw7XYgviBxA8/6SUyDLP7TMr40Anu/Lf7
VB/oexNlyDinzI6o6IXEITqee34/kWEyawiToNwarJLPA80C8s515OjebOEWqxNjzGdsOC4N1Lv3
4B0q7CqSFAyQPVBdIV3338Hf/yUcqj12af8+FCQXJejLkC/jvupoeduH/B5K+BQFMFZeSo5BHotv
kLnwjH8d5wPhtnk0MK1RcVo7FCgFEwfpen0tdnR+5fdPUmK6bh0aFcKvm5ZffddZ7zDpfQ/2SbYt
Kq8N6aESctZaqSfUZzNZ0iFT6GbtrMajbfUT13UnZOPW6fq+vCbiZaVyFGXY0HlmnzZwGbKE848D
TcDQ4NkeNGvbz23DMx6F20+GxPwqTmdt/ys/n4IOIMA0pEMKkH2TTUrsVhPeqBu5qcOVBx7Vlm0K
lV6GmAVTTjOALEXTXD/ejvtMEIlAETewZJBFjyJcJakp3oCWOF3hGxzE03XHxWdtkCyOF2XZAltP
yZeWNVjtcUkrcRJQYdeV1klfCKhS3DQTFtmvJDvuaej8z4shlW9HzAUEsAHxYcjbkq8R1ljKeNpR
tLX/nADOMxTZSQwb5ZSxFDJZOCPhQ8jRKIuFViREbi2EIt3pme0cWG5MTo6VakBYBw0V5NaDK5aO
vCFlTR/VvSbKbnTPLqaTwKr07Ds0Hc8N951e8smEoxUlsom/Ir2emuRDIjDUEV2I1c9aouYhKNTG
pVqC1ZZdG/b1gKAH68mHk9bMeBDzprjPGHQ8mlMqOGukWu9AIQWmDUCrND5OBBiova5ZsJ58XGHr
pRVGPUOfOL2x7OLOzT9GtkOrh8d3kzxLCZAA5QWWLwQZC3nielFVAeY6GVaUHhRc52t+AWRdSVAG
faOGs6MZl9PEpYNGCmdUAhVWIh35OZDkkkXqwpdG2Zl4UsDebzpI6vcEEg4P3Z6OcdtuDWg7dEoa
AHx/OYwHJrPvXlyL1fiNBfgdozGORj6OQ7WiuhHY+s2fy7GwXbQJMDBMcPVS/qb4OmYV/ZRdaT3I
MGPCWtKX0vcBhuhQEGEupQbTgzLxBuRlKwxb1EXj57dvggGzRYwr4Jt5rH2eBSEkIKYlpwiFDBzh
57ics45ilSwzn4i1s56ZDDDmaR/6ZEejKGSbUOUqlGFMmsetDocxPiNeBxSyJvt46K17S+EZ7lEJ
paI7HGDzplfX39exUVHHx/yTAprZzVDMZwoTPVLNQ+bfzd82RaPVpkxJDoNT9Do6JIqYbk7U9ag4
6KjvfZ1+MdSV5rLav7voIxCD5C787Vi8FtAFCj5c6frEtq0q4tZr8brJ19fO2JjnkGTu8gZX3ZVo
hKLiKXCMt03CYXfW7rbfHX6s7dtDtfOCIZ/p+NvPFVnb43lzB3KwuRy3saApvq4Deo/uC3omSrWl
+NcRIUYp9bbBNhH96uRL0f6UJ94qyA7eykCg1BgX7UuPbGSiCdxG/bEp6HK05cram/6LnSz9/PDz
WE8jNeFtlAYIDdQtB8pXdJwP8x86pSPGrDIshjlOPa7m7sLfyqG4SUzT9bgeY/rUSL2YxSykI+kh
UBdSP7nbcJgThrgs8abkVSV0yivemG2355/cRLI5oB3ZE02FlFSTbqs7Wr6/EuQUXN8wx3NnGiPm
lefZPN8hsomud/wV+44MpxqALP9bpD+gnATEWhh9jWmoYuJZffDT6J/0sECzuEVZVX2j5TRb9S4w
seTt0kgTm45CuVGa9k9Jiiw76o/2C5PEtQBt2EUMAGQh5pCDHQTgzoy2sQMohnaSnNz27Dje5kMl
9PwyigegttoWKtkgYFbRqGZAVP98fNynbVUHpeSqwxXXPmgaeYxHW7bYl5klOv/9VToepMRFVT6n
B/yUSHbrNTYTCNtaezW4RkpfG1mfE4uYeVlJFFwDlJ8aVSTbQ448N0MSZcaCm2nCZ1i8FGzdjmXB
0c2GPRVCtqstTSzIw3oty0g42Cra5y5RtwRGrcGmiJiWxQQhwaFfSGZPBFEEcUfbJ0V3utgvNX/K
rPgpBd0FqonQ0mUa8HKiYu4ZJL7xOdpXB9xR/9i3v+7sf7NE3tlB0SJfDME9BtQ8lUtIBxSSWeFw
m8mS+Rzx1yArxDebOpYRt8/d/As29ZveTi1Big3Zv0gAz4iv8CYdgbdOzAkR1M9sY9BsUkGekXdB
oHyx4uB5mBJElIlgXVr1+XrwD74lsaZlmZV3HIpLPlabW0nXhewZ/VOITTJOrqCCIgKHnQKnzJcz
M/q3iUUjqgl0tIx8hGcaQjVe3I/kAh5jaMYQ8Pv3csCcWZNKpAPNsOMMQA7ONHIlAxjDFlz6vZns
6Y9vUvoB+0FPhf+qCAeS5dyoER5k4t6jkM0XO1SIHRBolMU4Xjycb8eqPvEt21PRAsv5Z4aQoNjQ
kbcWwxppH6FA/+7AktxoJwHY3+R1x0/+4xjqMoAf8PZAbvopBCCF3uWhDwLndcj7APS31rqI0bsr
WHK/xyv7Dm1DNgU3jzMLc9k//ccOEo8B03M9M6TeorsyjdIJN2lxk2YSYxFFBHfYKuA77izU6MPH
cCdeKxNq4k/6RuTETl0QqGxlbNNmpg4k+ROlAfvVwXRB1bB/CJcA+HKn/r364Q8tZv43gPMpIgq7
DHV6GnnPm8GGm1S2dmKOgrcrjEilzr31I87luRsDsKzsUYNHbamcZHakRCu+QF8lLt328iCMji2o
QvHB8cCnYt2rxN0gWOaIfY4hkbkqsuvGigku9aqX8FMriw8jy13+/NR0V8rDTMuDw6Mr7RUplWoe
GK7tiLqu12QQ+h9qq3rF5YMdV8On/V8jYP7eGIPgEGrdlMv6shPGbU8A4wyKwye7ZaA2a3xzZJpK
3MtkgRUcWzMuh/nC6A22sle0lKw9FRzELAf2hrvoNkMfXSOPO+atmgQ8ZMr72SYvWQxF6oQc6H7r
NyNAOQmPgttzAnTaPspGevN0ZtRxFWjc1TmGk0EAWOtop3U+Twa0rEhkq73ZQJNbFFVM+JM4bGZ6
zH69b/nB9wAMw83BSdk11vl5H8A+EbbQ4foLDSjaIvkTqJuupPKB4yrOJ2GS29jWUB4jzPbFrIVA
yk7L7OGHU1SLd17nso/NKJkNk2D4zfY+etcbRYPVF2z2fD3E0/4DE28vA0Ww4EoVKlNUSLwmUeK4
/qANrPKqLmAeypsN5zZLV61v/+Pf203iDSKihsuVkGo7m5ig7q+eYLViB6Gwji8NsaF+FGmoLf6a
QUJt1mVtkzNoasUyY58EsAzHnagz7PRNSTWzhrHfZh+wkGOXORXCg5KZfhtt41PA50UUfLGBDn+E
V/oP7TwIcVRDSp2ZAdT6aG6s09fUNdAHLWC3zioiNYY98YGo5yn8orZWauleNOklDvKJcja9dT+T
epP9p51wHf6srq+BujhHzj7QHbjX7MdpyuoGFzrP7YWpUjLFeiz3DKGL6C7qVcmoTcRkiqf5VJ4c
3W1/qbodh5RXlvmNCQikFhq2apLqb9iuxsf2nErsrFzzPsGyBZf7bVL3zoyBIk/8F0kKmrRdMjw2
gqbMQPbRaNAZJSk+X3HaOnRdWHBBxlHARXjPddzW/r3w1cufkBowStCjcEFHNZCoVxfBRayVxe12
Sf6FY1n1L13uEQ3NW+Tzg0zJp6TjTICqqFZUSUBFfvBYRBs5HkzYdQrsIbiyjFtqm4DBBlIhTI90
cVwXOsMzL85Aopen1f6/Jf0pF/flRWRp1zuo8zuHyhDHzB3WGVLEHikL5eYzeANlGjLw/ySs7+zr
oU+5Jses/OLGsIhnijkSbxDW/N1Eh4zI0fY86hDqZmrR53wISAF83lJr8idCcQDoUKNIKeAOs3M9
Wd+eoclBBAxmtJk18NnrrG+ZCDudjD2Rn+tIhLWwJWRYvOw6TcH/L58FBSoGyL7l1YrPJYrp1xnR
956NClpgZ6VSRGBRrQkI0dmAcqzn6Mz4L5k8+tTVWHNbknXpWHz7W7Snv82zM5Pin5PSZZNwmgrT
HXI31sqdIkyzlR/a48ztB9AldHW3MUmit357I+czWpdS4xhzHetIJ0xgigB8urItJaemnY/VipJb
uL5ix2xPghG4/X3gFLBq5/3sQe6KSDZImgaZHfeewJMNGR50SID3EzdWKScX5o4oN3xTYNrDfNDC
YPCY9pp43MsjIpq+35dGNNwPiUgAhK0iWwRj1bjn/xGttH07tMvWCIuhMaolo7VRSuuyesGtZxpH
0XNRbDzeqtOe0uhdnN5FEWF6Sf9rMxPuzHQwY72++Pi+M7cUUmLtGRXNsPZmXR18HIIa/jUzcqJZ
hr7jUH7J8wk3OyJePy1jsaZzrqG96eHKmSwcI/QajS8iI9/uRqYkEEyQxhZed/OmlMT8AowXeKUt
DFSKUMWqMNPFmkxZT1foIIIJLL/x6xOt+As8ubclG61LOZozOkykopxyuwrYJb1/9z+8bV68w2Mr
oiWkQhn/lg87L9bxlnXepQTqsWn527UJIFY4CjHm6qlBtzXVhsH53CXyUqmjTQC7hPok2FJBrgcS
/QIPrWKEz0HGnnpqneSl2UC84nou3lBJLgD+zHvrHSot2io8V6/lbnRgV7DtuoEQeZSbuf1MVLwN
g5DKnXw3FY+OEbhrjYe+NDM8Z65c/BlahGy0M3AkCcJ8f7neI69gJLlNMY4W9BGhe7J+32gdMR6a
fhd8L5zltK/J/agBPJ/hkcKJh5+UwPtR/uOfpYmjtm851zqVRYmUkP2Df25QNVrdV9kO63zlmGMh
gfOOmUgZ4Yawmb/2itc+brNSI+AG5oTY9NxtMvKsRqHBd0Q8qpR1eLNQ+6ke9JxQCc0VrxQmrosx
m/cK50zDqEPCU56Lk1LHb7tZhBy5UsODUP8xKV8qxJx5GggB49C9MJMcNOxkQ/HVXq88mgLDh1fV
yN3J9q1A1d/6GEsUiIwvslF/Z4GeEJi4O7Fp9Ykc8eZNcDqkDHZNgQ9si21XsNLR+xWAOEdkYSWl
qK2oDuql+YmhPGEtVTthOfm/AMD70F2q8B9enPma9tEwZzghZ0KKM+MCXBMGSopegamoCvYPg+J9
NqxkVRzzJ4U0aSrgdc6NWkm/V77r4xx40SHizvWtkyIzgbTCzSNqYnF/NWkVjRJwNIJgrzcZU8br
JL/0ecnAiMvs3IH/kxRo7xIDu6QiKvuOIlZhES6ryGEBY0sZZbk9NxOuNCD9wYw1Kqo8jmNwW9NU
6hwrMsQTMAtx3m8wsGwFpbx2WSomrxViJPdyOBIVSMi8h+nu+FFzdCtOzrlvCJrQc60mWXozaUZ0
ZJisATQiiVQQQbFw8UlVzcRWvMa2EdQS+p4kPzZCp/X1/3g58J2bI9xRTAoNTS/Li+YvCULhi3rX
9N7g0apWGP8C1XCpfRolTIhe039b4Mtjt0MFpvjg/trQ4rD4k9dHcGdxKQn/DVqEVlrtGzjCxxKc
cOdIch/QgsPTUkEb8kgZL1mxfF/NQKR8N5O9AmFYgcmfQ5FS3VWX6d1SzCchKCAbx7lb+KsfgDT5
qzYf0qirFaMNOhIVlkkXgrdOlvZdjCjzY2kMNXkSiBF9eFilYhgqUQVfhngPgjamc/Fni7Z+8xgy
YoWHRS5UuoJa5sj7w2BTbrMyeppuTmVFKfzg4K1zQhkRnYT7OCS+pyVdnF57l5H4mUnvo6IrF0ym
S6+U1woJDvfVVr03aL2+wLIIwRo1k/ASHerFqdhDPapSNRtFaQusKLIa0ICJw5BGb2yuzwC2s834
OQ0YLbIZuRRyf4a5gkzjC5SGyKy+Htm7/g3iUAAT0MFs+IRX9hOqHNL2CCNExAmHxyHwVlJvwNHU
EPKqvSGOSfCwDKOZaYgMTDX0VW5MWYgWFvkyBXZThFfIFyaonVXhyIT9+NhnAcwiaTBJ0jmaVbnN
J9uIqlxBwcS+HOUp3HqxCrRLE7tlXpLzMNZzTWI4Tf6Weq1aJaAWtr+gBP4+r/EIaUSdN/a1L8dt
/+XY2zW/uyEeOs6aVY/r8fgZqO3IOXnxuaPIXSGu/GMZlzxlp/FOAgJm8hk9LIAi3KdrUZ+aUupc
PIBX5PAP+hSTz1TI7y7iKS+N2I/nvt5NX4N3ASL1kYgdQ7QOmVvc93ChCr+svpUahLN3xGCGzlhI
WCMzHlas6JjvT0/1peNw4WR24wVT65SNHKCLWhfPQZGzbcE4NZ+1CgtkP0b/Z2kf/UUE2zv932eE
/0CRTkI4mTeaCZeLGzwxXMoe/vTNJ03l/iLw4GaZxuINKg7ep9fVUjHUWvOFqg3Un3vFS+ixTItM
fke/48pRXoSsOL4ellEg3mgvBsoGANx+heh5Dz9czi0/mNacsRc4PFjclpEdGRHGkgiAIFIuApOB
+Gz0uT5oDjfPeCzQVpXdb8Vw178F+4CBuZtpC5TFLVg5IOUB8HJiXcEj1zfKU5ofarlmUxCNP3K6
jK1nxoe0wacRHxKzVLOICjWdxr0Ez8j6/kw0nMbSeRC60CVxmSoF8fokHayxstWYRq7o9iqW9dA4
gSI//oez/MsMugHISTOiWEMRncx0CtI3MDQVXGkuxgGi+wmY4oEj+RDxLekzqQm/IOs229+EFHbl
mUkLWtLyk26TYVqhJz+l6p+q2jc1mxeAPd/P5U6DWSo1hay22nqzN1PWhgnOZDU01nClOYI7Qg/+
6h+3F6aYET4TdAXIqfQpaBtBedbTIukwFKmYOW4rnCtWXVfw1UWmyiLPwEpuxcxBezT+NTOMe3wR
AgHTaawHaAIlBaVzSJJfbv7GXrVeddsYF3zYkrDWj4kI717n6QUxsle0ZpBsuA/wohy8nKm7wMCd
ptcOlFM34e1vnwamjjqlWCwt5Faz0TGyqjjHJ+1/5ir8kruudnJNrhlp60eM1Ixk5S4CqifXntd4
Udu6jSKIYi12X/uf3MkycqkjlWkmpkAMAvJK+4dH7DfAa/6PfYWhxzxvSzcS+NVvq/vvwdNle7Ho
9OgrEsaBQV7YHCNoQSplAXeTA2YfvyEB0zqYBAZBXfxnB6K99W62ScAukaqC0d8Bi00icchz28tH
0ZFZo2MPLCgbbPq+Be68UZ+zahFQXWaEhBq6hUC2ccUSEN7rXlW31EUJxmhxUdQOzxDwXZgCLhhp
8W3k3nFy1bj9Z74SDouEAuXk9gAhydZxw+hl6qBkeVWkUKxBcHVJk5uKtwf3QCl1YHq0kWfeAhkg
navWZhhXSWnt93SO+XHTHNnOoF7W54ayEMtLAINeyIJF3R7EfzWqTwr03flMcaFNqyAvqe5hwIt/
pUB7PJTWjtp5d2N+eLx1haOCPKUL4d/beT/dj2OtGZRkInI2r5wks6/sqDgYtmjK4qVgrkCySjlb
0kmYQwQVI2PqYcOvLplOUnM9FPiZWjMQQYWh7w5YIn1uPoO9GW9qONPzYbrI9Ll9qtVptqQ1Pk/D
8qTeEoW/zqpAokYcmFERwzyhY8QoMsSOMYzjDmNSz4RLufmHd+fLVxO3IT2udajRiK/qsShGuGp6
eUKfhDhcPzkRuHPznbG9sklVYCt8JkKvlhEOvAtkvrT6IMIXsp4ogJX+3hEnNBZy/xnhg9BY7U6N
HuqnAA8m6pfcrOvYjyVMTGCvsD6iA3DUCzjkcf+kcyIVubzzlfC1WlsEH6iVBuDvJV/e8OhAErAs
uKf8A57b6mWJVCTCnYYQ/22Q5AsQVE3JKYZyFg67xCqQ2I93LrobE3SS+gJkSIxx9gkpsEGNmBVi
zNUlUjpALvGja91c0nTJDhM0ayJbm5gw8iyv4gZPhtrT9m2GFWG8+v89pI6LXp+A35y+V6K1EmIm
YvnXFGeTXE9j4GIFezUj83te61+vgjud6mhYsQSMs4rhD3RX7gn3e1R3Pr+Vb4CSLizeOPBdHGGP
Vfwc6+SvfHz4MI7gK1OyJzS5heJ/DqZPBC2ByTtELFIILVo4hW3h1AmA/v3+1jLH88AL8g2GB6nZ
6qPTt8Gpza+Av8Hm0eEJrutzg9uNP7C741lW7JbpsAj1obiV09rRF5uisCAKPZTewMI+ovwfA3H3
IzXvW/8svdybyGyx+fVw1YJrlSETLdOqf6majC5d3oyBATH2UsI39b1PyHqjUe0wYu2M2eaPJi2G
eBvR0YlKkWsAU4OO2IaJU9D7DN9xn4+rLWN3oZLY4SLQOc8fb+CcV9lRQ2CpEYnANbbhl7qBR67p
YjGwTv3c0gjGeglR6mIkVAVr+/n/nJIWWM8H9d140K3FVLtik8BqClsbU9NJJxecaj9H1XwgZEAu
/OQYzKzde39+qPGU2AX3K4foqhSZVnqWi39Al+p9EEDT9Xp9S4CNcVeVJsSf3RE1iz+niRz/V/3k
FImljeEcPDbcB9IaJhPcl1R6MHAtts3O6NNuJaVJl9DFcC1Sse9KEhuUF78Vnxa9nfMaNJbRIH++
9NvUInno7EOVgAMyUftjMlznp7P5VR1Udk87YqIFXufhkICx/COddrOXNNDhl3L9GtO6RglnjbKL
cbIn7va63RG4WJaI2OZhOeBm+Qtm3bcoLunsmopH74CLt20D5HGozNVNxr1N/ovIapdHVcw67G5Q
mHmhrIj1oZMXfOVMfldPeT667/d8Ebpb6Ggc15pVO4L5zPE0vHL7LO4BnZm3MtPRmsRmE52lBdbo
NIJi/aqQPvI+Gap2ywjhceIyRBYv39vypGOUoTmfSguDp8tKVkayFC3hZL3TgbgxOPE8CBVMji6Y
0/BMjla6OWH/hm6oTspOTA+qQW0zKcP9Emd9cIsDqoEBVL33KD0hS5pZberualbZYWCZXyU9qf/U
RmYGxft8rjasyqWmQ1C16khSRy6my+4h1+y6BqKIoJ0vDo0QF3bM/c1MwjvjOBdpcH/qNL4bWSbl
Ma8fS1QmCOOpvbJkNQodYQT9kqRg71oneTE+ppzIvrh7h+k1WKXCF++6OfBH9tC0kN+6/pu95BrF
+73hqTqs16Fj4Mppg6TgDyM7+5N0G7Rjn5lBT5TSGtClbSq5CsLXHCAS5kahQ5c0izkV5XUfBh6M
kPm5xE9HDn+TAixffwVU5FsIRMmc4W8vPNP4UBLJib4bdKPmNi+uYp2qjFKAHEoXDzodUW9qzIUI
pdUBDYYuD6QVyqUR1jZE9pIaCkCWPCyVyO2ix6yU2GlsdeCJ/2mkQq7adk8RonvA+aXRcf4bbNmA
LvHGk3mMuagzFE1GbyXZWMckH0RxqjrfV7DE3hbbPh8TDmxwoqa/lByXGzwJxFZr4Ibu/KXQml13
gsJlxa40X2CEqR7iIuXYtd6qfk3oU41Pwggl+RTXuSFbu9vTwEplRT0B+VT5H6/MWQ/FHNgjRyNu
UBGepwrlJechOjV0iL3Hp/8vWMXj8qXcSHiDJe77ZA3LaDx0N/eBFTRMI1JGSy1T65zQpfeM6cnq
pO2xIovZ4gNQz7nImr4TUlupEONaHXdDUH2hGS/lQBXrRd+GK1uFPWemRPlYUUQAMj2q+o89hpMD
5RzHafdgmpwmbQDq1+V8fGq+ornTfj2iOUG4jjUyz8W8DbYoM9RvWA8YxABog6aTnOqdqdpu+WA8
Ely8jYbNmTpntdrySda4rAOUpMClktdcLu/FjVRjRmUcu7z4ljyTBv5rEf0Haf0jZNPyntc/MESK
lxtjAnSBEPrq/657G1H989N6b23KHqcHWWYGNsdfsG+toEEUxuvhG6Z65IrsQgccMAJa3HnqKeed
V2RO2b6F8JLyN10DQjCMZR26ZJaHAGb3T+7V4X1IwpfYbJ9F6z3q253J2mIGHjGS5dHDCRCd3LjA
2Pmo4ep9ooshEZXd7vnoKJO1mIecmbmpostjbHu7loSaI/Ke2ybWEcI7VmgjHsTuSWnCukiMVPMR
MJ2Er6xYwrbt9y5XNenBjIQWMe6EEpUUHGoKPEAQU4BzX04jmCh+8hDDjD8qTHb4mH0hzaeNolKe
EumR+7sBwHyAZ6hUF9zdC75dNkx25f8P4G4zHUgaBQWp/ZHTPEluEE5YKPS9JO/YAwJxD2Lj0L5o
QVP3P0F3vfC2LLxCykkY4b9Qtm0AgbUgWbCT8ix5JjP3zP1d8DrAm7aa1WJ3wDwHo+Z6xJO+b74t
BctlcSbRDl4wItLbP3ffQXdc2+OtxE12vYJGlQoRAMv4comT2/D9ru8diwLfW0XoqyuqFUbb5JOX
Dhlt02rtzkJVkJLzh61nu1d34YM6MxlZ1eXm/8KO4GauKNC0MAxh1+K5a3U5U63j2rHy32+ModIh
t0blzEUEhOIM5BYxH6Ikj1q4POLcQJ9KSV2aaewgivozHDXKUL37CS5fatfli0ux30c4Pkyg3dia
l8z+F/Vwi8aOV5IMFqPUHFvOPmwEGhGrK3mbsNMicPbneHXsSRuRYBtb1NssAEZdKmrFwUmJA2ip
1Yn+JyeZoii/rSZG+lVt+YZ3y0K5AFN6gIUAuCRMdt+9j91jmzaTDHam/zTsNf0zbfzSxZobh01t
WV/UT3+iuM4qF9CxJC6QXCZkjVJPAEiYG4p1bBSYErsWDxLhbPKCpMQlXGFY5UhcJIaRHs9Qj1tF
Ru4JLWEyIU+DkEvphPs/7qgyJXnnquCXFORDnn1OV13onSgObgFvWetxIdO7QuftE+2r9H3ZWGxl
cKycpCrKCZTu/60ryuB+ngrmhbcaq3zWXb3jFafIwKw9M+BJD9pQxsOG8zP4aWMWw1A5I6uqeQQv
ISuB1y+1Ku9Y6D8+egnhZGwDvmqKvpawD5RRmviRyAQuHYrCPtvIkef+crA4VmHNkUxGAVpR7XRu
nH5GJ5zMweLTxbXqPCpJzBEVbfRPz4KiUnV+qxwm74mbcuIj1eK1AvYkIwtsbeesgs3ydik0ejxb
L0kS3sUubrXikYToDBehGV/mw3+43WNMzbfUbCRP9A5HhL+++Gw+RqmT8AgrdLycsvWE3NVUvSf9
xQiN/Shw2E1Clzd4dg1md0GArpwmrw3hgfdlBKqfIGYJylwrK4WgiCmJAC0uK0kspDQXFsNZTbGU
Wv7cIh0nYXeTafSIc2jDFBR9agZhztSUT6+syBYCrx4nB85HxAyeWA1IXv+ifNuHQOoGQcvomQd2
QI2Zuh3Wzvkf/OAJ5BRUpYTFQlybx3AHQvkJRqWe0gM211koOkmKbRH1JetIL2B4uUTIX6zjnr69
3ZBPukKBqu0LdlzEPBhxBCq3YruO8YWpF7YbtwsT3UBe3D4YZiJ1fIBZ7yxXGR3UqRhDH7uPngZs
r/gcgg1X0YpPEfeCaZRX08o+wF7ON2bWCTkG0oyXUAg0Ci54Hq8yUYWNHNuMlbK4dhpKxDoMRiZb
a3NTvAfxRw+Rlv6lrLBsOMEkirL/0rRCPDYJDTnhAd0W2aj9kC1qNMFvtXNoJoSSz7VvBKxOrk0k
mBludB7KC4Jom4uQZIcp5AqZJF8lhsdW30hCiKtVXDeLsZEUYn5TylOIFFEjFgDZ2hRcVcjQoQs2
g97fj2O++BsdHZrMLWuPoccalBwexEt36l5M7PBXBCkAWjqEdKID+wZd8XD5YOe0HnFHhIrreVjp
Edwi2rEvCG/UurnUUDbzeXGSw7vcoKKUTXoCugxaYum6dFgp4fFMd82nn7tiPOmn3rimZPx7xDzT
muoS7orY8L6BukHsXk8IIZHTJC0Nv5Bp0+YYedJ/+hhJ3wZ+Rwhb4L8HXv0Rd/eCh4RRNnyx4pqT
3yA4kHWFF4KUXBfLY//oQRiRuYr/ep30d7H0s11LnwOWgXjccW5jipuHMinPw8Pcqb1vVZdlJSft
xUe9A018n6aZpkzcz0ygS3TvLgDwx4xfNYSdfpbM6/CoPxrk+C9bBx2eOCewe0N8i1nwb4r0MhfG
HfprHd36Poklu3/ZJsPkaM+7je9SMxYUJ+0O4mmuuMkor9G1ybTpunJt2uI20f7AmiaC6BRM5dVG
2EyeK+VlEVPTcQbbaMQ+rvQk+bcSa5tElv03RMqNlskiTdLqh2Lov0TtWzlZVTGkwdISGI5QczC4
6ppWGETSYfw/kSBVeJnqq68EYRdAz7VrjXNhELtfWBpfxyyelZbHN82QezKQAkgCMrg4HWKq4uEN
PyQpxu/PpAW+gKuf/Bi0UmefHrWKLHKe8v81f/WiDgq8bih3ePog164I7YDXMjWeq9cnhRe9gaQ/
WUM8BB8w3lCTgiU4NhJI0fHoYjzjjOxX+GB0wAq7QNLieeOhBmH/dz5N5qo0tn1izT+hAxPohRRU
Y0nbX8IW0NSgXou/zT8Gb91DmYZDPa84VX3qylTJzMcI/KnDUn8Lefn3C/1KMyRCS2zt+rbGJ6pv
wsloqdwy/yycJrqPad4f7pnxKqJ55HLES7Y9kV4bgChjctQzFy+4ZYvR+XjTHBTawMlUBidUgXVA
owPlCGJu6w4dZJyPVZQKR7xFVQHE4i1btN7JOeisT6KuHNwJ35BTr5zaOBmjHt0e2Udf3J37+udR
5CZv1oa4rlMce8lTGsyclRv3q0LMu4ApCKYugd4X4QDwNu/puqOKmYLvKZCYSsV9BGZ1ggx+L7vX
dcDjVmHqVRuJ8E+TYY2c+NHgZPg1SMXSpF10dvk4N5g26DwlfFCs4Prkjx92ZxyDoHLBk4RdHLQ2
h08bCnUqKr+WiLkhh/Th3Q8JFGtCN3hMlONMxFi5dSXQ442p5QzKbJjohJwxt0ygJQK/eeIQEEsu
PThzAZM7yRnQuisCqlp52OAP6ldg+BT8n0cb62+vxwx3Wcy1GEUX7d87bb8OiroELYPC1iA1uZB+
3MVPsQnz3bRCslKMg7rxpwk/psfBogzPQF7T1elJBFWwbnZ+dIFiWKgwu3w6yIODNxIj99GBq3zD
cobVXg9aDtMwIDBJ0URaPRdCUKzPb6xTdcreW0d0G86ax+FuoNIw3DL2cr1ZsMHlJeCKKnkzcqnl
lB5AilTiTtPpVBG4JvqhmXQ5qWRcH5bdDaBYi8yZ4jem/6FMaEeDGtMJCilpo9JXMIygLLiL667c
3eim0m9CTqgVnv1zDhPXzzpE9ZgeZFPA3P2lDdOmv07huylNaKIZ/ubHaYzM0yg/AVsExTWIMl/u
Q8WR8ul7WiceDDavHbCPdO8lppcfdslk7uCIBDyGQHX1KNMnvFDzWl/tKH0FwwwwveAzcM/H8tvd
S9O+eo4z8pLgMaZN4Kxg/VtWYlMHBsk0miFdIZzPDQRRl6mOV2FAb5MVV5UYemv/mOOFbhEIJtaH
KYhONgWgR+mjQswH2ivwXYq6w1QlqFkIvEVMRUIZIDOdKt1ny6+XYBr7FPFzu1NT2yQQzlI85fG8
Dn2rz1/Ao6OqloR9YLsrOYOKE5aHhfBms0M4S6qEgFj3ikmjVRiJGTm3SxrevvhR+LPI8pkov+1B
Nz/Mjw/bc57kwWO7p8NjIlPiraQ3OqvIRKeYudEl8fPsxz/d8sR49QC71DrgdOxuDmR2ha86s3+l
EEm6IIFnJbwj9fgSRC3QpzMAtGViN6bXacbmwD7W1vSDTHQtmW9SnU4nbZ4MfSza2eO0EI3vCR7j
qYEn71scZAqek+wq/x3ADf4vwe6X5jx+01XWpViybkH9oOemZrIwsw3VaffmEDkHAxYmtsrV6im+
oJARxYApgRSFAgOe2R0cQY3bkbpYyIUli45/Zmnrt98Yg1Q4IYkVLzp1LP9WNUx+UYmkByuOEkwD
SLPdtCvZ7Ygq62oQJjv6d1uocUC1qo7KB+C4bnqByFzHFs4TkrwO4vRUwuwQX4/PhRF0NaMdVmpX
SiBDgo5HJuCXuBf/oqz0eAw3wEB7VVUkLgbj4yVfAxg8f3b7qXTUjogTDIP94GiiHTR9mC3Y+gWN
2uF9mPh2uePxvihwEYcCKs0mI3HUN9jeguUWohFxv/OIxEW5/lEF3YyGpsG7C3XTYH0UANpnD54s
gHEVH8AB64zy8OmBl3EOYedMmM0gFsOUN5qam7y67vNJttEuniw/gNHrL8JJSRmOuyP1lsbMoq62
ob14+8yyObHdirBrDkyLWVEG66V2dv/vbbMl8j5/SOllTmjsu0jeVKbG0U3jWryWmNTgXNd2Iipe
S4wyNfOWpr38H+85YhsbafcK9tlNETn2XasNg3vPC2hal82Y5t6V6uVJQyJkDyQfaODuTAmPHcQb
uGcf871sT317ORza5eKPFfWzizdYemByjFo7FNxt2Sys8lErk+xN3pwkD2SZ9sLtlLhHcI53HGlR
jOz3tNK1nTD/4nrTcW0uKzUEOFH8YxGJBcODv0lmtGGDyV/dAkGc2la4qKVtAJvrEMuk3dig34qE
bTqY4BGpAO2wWYZDGt0iGjWHKFQlqFts0ekQ417B0xFrQlnK9W5WkFIGbaW8rwDR+LUWSYUAOImI
7XOwx96d7UE5HSUqMBjq6V4BE47ZiY8xKKwYpi9r7G8XVauGYcd11HQhdoiikZUKcEr2CdqlRzYf
qvwTVU7Opg/UKfXJ4kElKOFHggFBVezfmiH4oZCBeVR6JS8CREf36L3/W9NuVjOvoCVGlAvgB9SA
pxkgxCRSwXCxb73cwe9o9m9V++kjM5CsoAQP8SQVHfY+9654SwJwGtyUldUXIv+PqMTAixx2+0s5
kMT4zAP8xHdaLXCJNb3x+Wae/SxTZThldejztwV6Fg01xfi7EVe5NhWJPQJuDVTZE0dyRDq9ZWVJ
r25PK0TiUs0pfUjN3xYx9lF/GxWKWes2v2tm7tW3bcCZetA9vi+ugGzNyBBS8F4lvx57tgwP7lGP
AqsaGMxx5LVPFrOtq64VytkbZxT0WdSY8eUbQS9g3veet5ZhCaZjpnE6uK5Q3BxADtem9JBBLWGZ
Usetwu2/2AKFgrvbUbNzEYF4jD0Ab7+BO2CYp6vyHaJfw/PIDthTyq5L11wR9qpx8TKzjWm2kMtS
a5JZHk/f0UwZk7psRLBd+JNh89ANj8WQzrlhoXBpg4+vwCzFINzz5PXh4rvmtvpVwgYQAzhWFeHD
H238mh+Br8sNPcykIQEXwuET22ovNTQegt/aq4XFwhdNWE4OFzL24ikeTJWp1XivT5EY8bnTMdc0
aCsi7Jb0xJruSHlP3/BtlD9qd/chn4Q6MSf8Y5lDZa6n9VhsW3bWSZXJ0C16dJrZJjIv83YT6JbY
e3iF64pmP1+ip07tEOx0TWfu/YDC5+Fg9TQsQHOVX68NskCNlPdbZnWBgbfv5slW7k7doreLzmOZ
uxT28NcouTV45wxN0EGXd6Mn5OVByJPgivtptFMJwp18jiJ6GDoH8mOlI1yHR/f8w8z5tMwISX/S
35di85kKoYdg57Tb81EA6xtseFx3gbxDV0ImBUvm5KQUiZEaps2HrA9nwHziEp0JrkWs/bXcPIUm
f5u7+SxqQ1reI1J7ipMb1eXGujCUfNmZh/6mjpdlmORJm0bW9Svmp9k2L5LIYrkGdjHEsJORkNJA
8Pdin1f8IiLjFAQwVj1Z+t9oBg6NN52RISACU2ivUNRj8ftbshCSRvIoW2oboAVoH/pha36IfLSP
OmSzBxLBKo6Pifful2QgukdLsY5GKdWxRAjoEN9clqe286bPAdyMIaZwxE5/I6/6s0qYVTomZivG
+Bj0RyXVUT8kyE9nEUVqOHNla9U6LDPYuwF829vkv5DcH0vtfZSftmuVaCvPiQ9YBKDaf1ASN3Bu
rg3pT1OdNlKRyCU7S6XQfiyI1fTn6zzIboKA5NbZahRfVK6kLsNarcXlxGjE8fv6CkQPMnuMqmZ8
W+xxtcLb3Gbkc9l/a8/XPJjOdsAQKAuR3rONtM1AmNmkGnpHzMpMjebuhRvOFLPIcgHpuZx5ZRFZ
cV1xxQFcKjypgUJBDIb8zGPo6YpzDqfnVnPsPnucq9QYgcTJKiE+v3WkSpQaZD+4Ekbo3h+Olhxy
DR8/q1SinosUVPPjgIKY7YgbblCfWzXLwiGnYul/5Vdm9ugGs0DK4xdMAY0u+/dMscpBgNHInYA4
ctiUxXYK8wv+R5/IKRkVnpLdmOgaBwjzOLSyIey+CYqpeaWz1yPGkN7mZ+/iWZY3HW07gglHmE8E
mqSJuAQlK2+fuM0gN9QrqAOGQcFKZOwoIJiDN6jMDIQ0YfYN+tLaJVvwpcLtAH8qEydwnPcSsS1h
MCCiw3UGKZy9usFX/P5q4H5kZBKl8sxd19KlprhoMrUELNOrVIe1GVYsx0Yg9I5/NrDG6lVF+uxG
pVx6vLKHVQ4w9zTXEV+doo0U391XVMK/SglIu23g9anjChBIBm9CspRc3RdU5y6zoVj3gvENsKFf
9RVkhE7lEBxvNANbX7k/7jFXi1h/REiU71+Doqb381CyL64ZBqvI99aO6c5Bo4sDSEnk5I1Y+F0b
/OTPT4HFGDIpNcc/DvDPxU7Bq6+F++e+FWUIP3m0eZpa3anJmLAdvDxkxZaC2aMThLPemT7tWF8U
8wwsEtthqq4fuE7e97Bv93fo7qzxrQ8cij9iZyRZP+64DkjznGmsRn6gynmle5NvXXIZ914MhrYV
SNOXiQRWqohZmj7llhmb3pq0ztpJl+YG/IsJJJsIlqk3/J3HOli0TU09PUIZ01QAQzrkBqdBEZH1
vCOl0KPtaRi4KcGe5tOyGw6GN1sHO/ubVNA9CNqiSi/HJUw2n5QbVl+jpavFXaQZ6N9Q7o1agIwp
HBNPdbvxvxzejXYhC+Dh1W5ufmlg4VpO8SgPPBpUnAKqlG2wG2xD6UA29OhnRPsqAZP9niIkA57E
Daq1za+uZZ2mshcpxrFNJHzO6hf4eoMOMKEbXN4V0063AsuNBmO1zOjthZmoH8oXVcvEMzclGN6z
WjoA2Y7YaI2+eHr6tCL2ea4ei23imkvWKqhQPxeOCYr5P3kmYFG9FcQCsflyofxAeFNlK0Z21H++
hCvVZokRtlicVSKb9Him5exmKf8xZzXGLO+Sey+gX7V3jY0EBaMvPkorknpv8uLvoz5W7RFGMqeC
WJkOEj8Q3Hu21MY8kwzJY2BVF2F7dPIgm5VTntCJBwfvg6rovSdVf5i1d1larDGSPix2l4W9L7g9
xwCuCfH70xULdtpeDCQopqWx7mfnu5Qp2cpcKzBmVC4t7Tl5rXWadd85tdordIKquUyPyK7MJmMe
xZSofJK04iJmQQiqSJ4GODcndvGZ/4SZxe4c8Pm2ZlfJ/48Jo3D1VnWhK9yPITixn3GlZIrCXQqr
+mtiumuLWbDwsDksAy0RcODIvvvLrEH9UcQzvah67GdQFk4JaiZjx1h3vVbrN5A7A4mos44CagDy
4PBv4mNavsK0PLyZMYT+bIxtUFXDesSNua0xHpyfMCMqoel7gj+bJIAfmZRdLKRphgjy8o01L/og
BBvlgytg2RjApHldhVehEpf7v0snLrn4BgCmqlnlggHhEKhyZQfmuNk3ZNoyx8Wxgjj62UIWqKdK
qTWvzIVFFcDCmRqpazxllKS0ZyETjspw9uImmUQlrjtBWK4Pkopy8HmKSL+FbOOawKNFsiylQYtH
kyQQpj+AZglevOT8506snZg7ZaIx2JjDcji1y1dtUYn5zTPGjhqPR8162KbUtjxQtK1M1KOYMdeT
WItMbY1NtAu7UlQtIi2INZi9Zlxgcw2KcJN10+rYlmJiaoxNrdnGxsWGtM3joaZKpQHs4rtKdk/Y
uydiyzSS/JiKQ+jw2gA6BUmUVkxAPveJfZ5+mSQz2UeMnFenNAkFvtCjXDJex3ZfjY6/hOURsRGr
SXYEHH4zfiwBn0q25vVsqFXlzxVU0iXwJLMSbTsGBuRBFFgb7Wky8dR14DE0hitGZoRLfBf+hlUQ
X3M+q9f4zI0z/kGRgi0Ec5ceUzs8s2EAFEvogL7uh4AIj6RNGeA6qu3Ks/wKEP3x94ebyRqDih+S
WJy3m0ljjO2F2dEF3+FCjqrVUxBTUP5N8p+mCx/7w2NbmgR4U/H18zJbk6VVaxCdGKXf5aHisTiz
7ZPFRC8wkRgq2WcizFE35jAb/GYXnYLz7bT8TlJKt6YQ7vdQb/kxqvCJgU6Ha+YNOR1Ufonag7WN
ymV8k1AWQKzfiFdRSfJjiQcHZJbGvdXr394AlXeyyCm9JsR7v6rKoJLzG8G1jO8YefFWQ3Ki3h01
cUZv7jkRTzpuLP/LjeDrxatK4tMNS7CZjOZG7vBavjaiUI1KC9JXjpQwOzeOnkKedImeS4+CmTSQ
iViN4Jk2s12zcsFmsxwkIAzRswtLTnCELYRhm0EAH6OuomJ6k5PlVreVYF+G4pXsbNhoIhHtFGTk
4XG391ZxbK/li44ZJz5OWtIOGB8HeQAr0WJGVD6b9dDazzIsGoUgZsxmMeE9NNJxC6FreZxHt8sc
9SwXZtPuzhhphdLUpD9sXLkfrZ1LsV+jHFw9j4dMhCZVpbA7u7XJVtD8orV3pSEQ1ZTNs0S/enFM
rsIBW2ofQUr/aKfOeamHn2LiBiYSK5W8mGxKxya6UpR1ohguiUNt0rXzeTy1OUbikWnbdRWPeE78
VqPhtK1gVfeiya4IbNJMkKnDRJdVMIF0tds5lQT3e+rDlr6KUVInkmeYIMASRELvP8V+SmhC09uV
RGL/Zq8DzBljsyWbRW1VmQ3aGGv3KZ271am5Dp+yRF1u8RljD2fJRtu/4bb3fUElWyyrGcFb9p/B
YgW/cxJ+YgMd8Wwry9IhgOr9lZIiH2+NAap+9PGsupk3VjrdG5WL2Pn7MgD6I28r3FJZkiBYoFf3
vlasbhPoDu17CVE+mBHeZiCki+e2oeF2Q92NRBonpauq6gmAgy5ZdpUJsCTKEvDXYinojGmCUgz6
rhw1JavnK2WG0kqJHCH1/6S2kwVNUQ2LbPUdBUn5ULdyAgQZoJQVJJJzVr/sLuVFma61QtbT9m/K
V3K57n41ViEGaYAxaTREBOjpMQX2yuL2r5dgFjVwjvbQ7b+9K67ZorH78VaImrSm6/M5ZJnKmiaV
L5y3eWb9rO42HmYKJwpBKLJtnteYAVdVs9pnT8pDLywXpF9y6g0tNNm1hv5VzxodlEZM97sffFns
P+QqXZ4Qlk3Vpb4pHhY94VzLtGXz+F3+uhYZ1MVlIOI7jH719ES0oizEJIKF9osXJcM0GEvs5ygc
cGA0Yrbzoxv8wWLB1fzo5JvY2TxjNyl53ZYnkKYZYJrk5LftkPRHOY9hfI/O0KpTgwP5Q63kUb3G
o18bNJNU54P35IU0rb+UQTU6eA5qjBijNcNApzehltANDEObMmjG1v6uborpsMYfdtZFOPCjUA2w
7LCByWRwniBnLn9jZy5RsmcxKR6IZpfAEIqXHHNiFMVtX9tqLXvKysBAfvqzO8KTCyT8m+VgKQN1
CCqAT+qjdECn7muDfiAzfk/bxpuZpMOPS43n/LyV9kMQqlifjOxvFVTTSGKiYXdFTtpDg2CWe/yR
n5DRArJ4/uzlftQqQ+3Ei0l3Ak19dCXiwF0ryFizDPLaMO9DBpfWxr8MV09C87VIId1LKGAv0AZx
bc3kRlFBOsimcvY1YSXeQJz2OkNa+B6MZNZmOHjS/CJXO/YEF3wjuSs/ELnc3DYcfZMVNVyhfd1I
Yb3V9peScDFyylkNdIP63sdmCDuAuXHbZRKC/701xGD0W/NmECJaC2MQaa6CvfoaQGKKtK6uYUGI
/Kv4kMDgISBY7A1tJAs5btMrNHnmh8mAB1+5SC1rbnkmyZ90gR2TgFtf63W9vRQ6/lmmyUGp6F+K
w/yYkr2aseXmT8zu80X+2lfj1k8XMeKitjisQPQjBBtqiIgPj3c919NowV0mVjy6NeHsxPTtEp7k
9xfC/7AQ66TmxAWzR0LWJWPBhkbCjJ8iGRmkw+EsVfDjPYTNkIM05zrTS8IL72wqLO4LoMxVsds/
vFcGpSC4vTW4qkR3EandF6OcQMOsZ+syBlWOOlGq6MPzS4b2XsOJx3PrD0JyDF+YHRyXBorvfVQo
BZtEwLZ87Hvqdhj+ToL4K+BRMX7Y2Ua3UTS3rQN8M3m/ta4lZZ2QRwwG6nwGp0NBya95blWLEfBW
Z4Yh340YDN/xokMpL12DG5DnQ6rlYBNiWBv6470Wz3hVOTlRQxaok2HWvJXnG4RZzHYehSAP2E46
ChNuqeEIoLT2M/TiVQ/nvsKSWGCJrzVT/wgmjlEa6MWQV7GL8o7kEcjURvndH1STNKidvckCOfnF
BiFs3jcYf5uKrOPkV2M0MeTmQoU5vCrRuQp1d9Yc9kPVcYp83tES6Hp7Cf6rh6ip9MhIlXRkx3do
91KgtLp1Uhdx0pu0JdTTnkqpsLn6eztMgv94/QhtOoOCfuA/j/XyBQiAzEBTr2qzDDqtODpilg/T
0dhY1dJZGzsC1+dix9D4ZFeokRwxhvGlnUFLIXairt9Tj1olutb6mGhp1+6xkFEdmRInTzNFvfl1
bbYEuiUzAVbb82zqJCti5TAO0lho3Vg7OFfE98PZWd/oUXuQvTCO1aGdosOBEI5GpK1mcMXNZG+L
Uing77ABx9rDeck8jQZQkbkKdVvpyDSUaABJuAxqENuVN6rglwmMe28nMegxjSY2jMO0e8aD2FaA
DwVMR3UrdMCIG3pq4YAuEix44M+uoQ4YoG3Q9lgcXKqq4l8/VPqqEbHfPNUbuc5Uo7Rne8XREkRG
3R/DqV39PscBOV4AzER3pwUNN7qQ+m1coCh5TySuayRQOd8xTrDnih6KoKpeNqsutT2CS0UlB7KE
zuSNOJVohNeIqconpw2nLRD0f/VHVWxI8wI/l+DHmnM6IM1yfb25sBi0DxYAc3GbqQ69Uzjbp488
BltVSZZOxLAbHZlJWuGVg3Aod/8ponAhv03y9u7RUnhFvVx1q2p/RsOHuQZxOa52pc6jZzroLq0O
jf3+DEA35TK1uOyuCPtzC24E2UAwGH09ys9QwO2Z7yP+nOIYKv+NrIcf8jK8oL3OJptYfoqJv5TS
7Dne4ekmf0MexdMpXLxdpAd1UA3vX403R5J47zIZqldex4BPp7Uk/tK3auFNquRfQ2rbEHZAckKi
DGLO5lAvMTrZ4GthMOp2M1DrbZb9Cdgz+Ia86i2sLI2kGjOTO2anltsbXnE4g1eYk0Fy5RiJFdYB
TQtS48KMl0D6TXo+rCrflfoaIj/eh2W8gW+sgdQ2+hv2KH2qiVuBCr1K3coGWiJKZ83BXJapSXjE
1M0h9IqPbYgbzSqFKlFPibRodT1YkmRDuimTqS4dTXm6WwtibaSIhuNmiXGpYYECoUbkyUDXkrH1
r3J3jhnYmIhYkk1jubz2YNgU9paJdPlCYY1b/u10LuAN2mlkQFVDTuNuVXY+j0XvF9V48cf8bk4v
lJRgJ3VEw9Yo6edR/4JdLz7N0iCFe0AcgeQMP2gCvUbQ5/nGuxx4QeBrUVTA2D0DToda6SCkzvlA
jgB7PXtfEZapq/G8VB7qfao+l1rIgftjXX2gg1i127VyyP1ifRobSQdrcYT9idnv44uIQZwG27bQ
E38iDAVAc6SHG0wJ7Xvyv3obBAD2ND5h7doCEwKgA0TLAK4kyKqDuwDSs/TmYJxdj2Ibu/5ijzch
Ktzgfuia7XOpoUP4b5UwYWIlnmhxgf9WV+agQDrHY+DP34aUPbHSK8MK68+pwgSCMld1TLdyBGvd
To7LCCqG+aMzlLOyNU/S+IWbGLD7aVhYjGoP+Gr71Vy5gdKAkHOq8TxY185oTvNrrd+emWKDAOAL
MN3CrXK/vHlNOdJrHveVcfeDO78NnbGGlwGBxP4VKse5FDdYnLrWdwMnHPX5TifCdB12HVzqRZm7
PyeHgi6kmjWvn9FCg5j58ObgGzohpTj+BZzgag1mq260P6ltxqATNQjdCfeudVgz9nY4XqL+I8Pf
VCv5/d0aBS4VPuWYpzPJlZYQtDcPaZOqMdKDAPNlOtm4PjJebWpqFFQzGBjnMHYvjuWGC1T+Xm94
ofrKElkhLacbTIaf80uAkYfGhG1kyVWLrcgLHH3/Wcj9ejcEIuyiTQ47/ay/OozHsogJyeYQzRgY
duFEABc4Wnf+CnufK5oCtWZEyxFmqT6LVRZ5NIiZlGK+1CKinpXzHl69wcokVSSfR1l1of15eX6Y
eC/q2HsdLIwXeU/AhH8zC6nB3jehsibG6aQrOgqS9UxbulFz81ARpNhAZXpGm99T+ZRGlOKiREdv
8q95ivd2QFF5fcIT/c9JnkiC9va0CU2b3WOAMofRnP+Iq+vJjK6ZIvfchJbp3nduGML5hMS0T6kC
8id80jiAPPh7DPELcGhLk55VngS8gf51cebmNcYKZUkni5M3+bTmDTdj91+Hs9wt5rOF2ER5UwKz
0FudJ67lz90Tn5+wzZIHIS9ZN8MFy27grJSfEeS2gRP0T6r7CWZxJiTTUVmu4ZHRJGv0j+llXkCP
YIuZRBcntTLBMwIhiOSWujgEXVNx3v5LtcOivJNZQGwJ0Ft6GHwC5sLJZS3RQ+XxXKle+jts3vow
ydTIHFSXJ24KLxqMHA4gu0YQ+FXT6Iz9Ytctca19uGSxlBKwjF5irUFCBK+I/0wg0mHc2XWW5Y5i
rE2oiwV9Udgm4UqjlaHTF4GBHTKFLpgyuqF0AOWbfqm/aae9HkBasjs3eDCuBmIptM+Qw63iKofH
pz3gYVe/2WfCpJ1P2gKWK19gYUlepLH5BaLsFnpHh9wW11J45oEkildjGF0IKPjofQ2bBv8LXVoo
gKa4AHP/i/ay0V3W856Tyak20K36aH+m2L7cwThETzw9OYbPDVwoUAkBdmG2AmD+Ir6dCh2TetYG
0Qs5jK8dGFwaGuyY1vv8/IFVcp/E7X58TNVyJi77/7X4zpmkZkdYYfp+0XJ2EMivXVcYRnhXzMaV
zbPpjnu92+OESIQIHWjNjWaqaOzLWQxWHJVAles6ZkIjdXsVbp4Ma14Fsb6JCy35gc1WlP+qP4sY
upIUZS1Q2SXzHJxBV61Q1zPt5Ij0adAdgLS0CXNyQZrOr+kd3DEY2+eDFezQturpcaG0pxzQiZtQ
oDTrdCnTKmdOjcFo3DvPlwODPq2ORGr1+U3vzJ5GVLi7AyHTDzAkzhKXqxNyaRoZ7gRFuWkprvjA
Hlvna6xjHtvEhqGN58QK6WlXQOA7lv6hk9P6MJL17b00eRdrxTtOzGUjPC280oikbZNNggpHsLae
tRywvxk9GSaPLSO464xuCyrb9FBH2GLzO0CoPbzZo26+U3gKLQ8d6Ua3idyT1M74KdukGhHhReGM
HEB16SSzKZjzo48AK3IlDTUihZD/BhZHrjQ4cTcjMCHPWroX059pNM+IeaBOBK/lMVRNjyn3BLEz
edRTwE40yzzXxadiKlRVtnINxnbdC67B3rCHyyrWMwPxCZhC3uhg1m4UyJB0JkOMjad2zY/35AXA
ddCbc5XsobdfOx6gyzhRlnyXKu4ncTBYqeUWFzIku7U+4hAmvwrP0QCmwew9WRiH0PL+XVxC5R24
m69LjSsIPpQOCk3fWuCc9QenrAmWsvBrlguy69aCDp+2FDsaPBcTgR8/5Svfrji1PDwJDIgl6JiB
Vdx/f0nSs9e+FAF6KtDbe23l/jLcFV2hE9Y+lDad3/iiJtZLnU50B+c8Ivg3Z3A/mAiOP+SUBS9V
re+N2vMW6nPBBfBSxqz0GmQYubyrFBkRKRpyIKdSOvtfABXEnx2e2zS2IWBwefkWH5tgadZgL9N1
6l5bbcQH8cQnHYjXcQ8IcLZq0qM7OuStP6O/dHxlmF0dsqMns2c90eOfVPnwptDBGlMvgdgIHhOm
x/V1kBOiJ+hVGDwg0NUsaNSggXa49uPYlwJdVowbpDoxIQmHlpr7WHWWCLNN8/DEXgOPoUpXDoGY
i7BQrPPyE0ThKmx67ykmW9X9rU7Wl1qnjbLS10T7xt91RP7aBiyX7KQ8D1lXj1IdE5qu0/O1L4bJ
OEUVBekjO61gmirP2QzHzeyjpPNe47lkx6ue8w/qb26jz3m57D1EvXyGQLuPhTd0rUO2O0Vvt5QH
vIFm3tdJnuvIanw6S1/lG9Vl0uPbMNBDgkut1cguSo0qXz1O0++UwtoB6lKLj+l3nhMH3POVnCnf
vBDHroWhU0WuNDom9PUBDgiDGkVze3Pi9ZXaE7qgWniSh2eaonB4mUm/msxOwRFVUDOMF4R0OkB3
x1PBj0T+iXsTrL9iNCZNjosE8CyqIw11JrO+YIoIinxls+obYDaghBrKIqbJUSpn/mBE1wBZl/98
SHfH6GxQNzkg/i0uxV5Yp5g/ts3na+EU7TnnSDsZzK1L7PTtS0dFL1TSUIDQZMkIaFrdCIYruBgh
Ao20AxA7VcML8lzpLMunI1X/amgQLIqJiEU93hqHTvtol1WZcwaS/aI0P8O//1IYXTqLQRaIDqpv
V1pM45fSNf0AfgV/eZQLjSs9wqLSkiEygDig7g80diR0FA1nLsNv0Lmp7DHV1lg3OOPWSGZH3rt7
ZpNr0neNJ3I5TTZ79pMvjRowG+DocOaPeEn61rCFDCXTDezTZDaB0tae/AbRPzFDHwDn/0xiVTbi
jGZjWlDE7fvV+n8Wm+BrZhYD6CBiC3fhTUcTt0VXgk+0iFOTyJrRDwBxKNu7Bzxs89BvqnvBtH//
SAR7tQAIYqwLscIiQqNwGdofL2SpWLkIrBOGhs83yFoLoBTthRDWEPHMGOdeJXb8ShUdLkrDLmqq
XkTyAfyryxMfbGn16rX0o2ZeyLHQksB75VX9Vuh2np5YcfRpObveTMx0azNW+oD44XOu9KKM0eww
hLLKp0nokEH8zW5v/RBUsakf1535CGZHDHuEMdooPjAJAkehTTNrKAYGp6n6ztHLBObRPtcovzuM
jOeL3QemWb2fSgsqx/3hk6DaJ3rYT7ZkRSy8fKXLoH8PWpI/6RjZQCLMmn315mk6KB13t5nUUA72
rA+v2z7loEfY/r5/C9Y5en1jWdv9uh8xX8hSiwodlTd5oTddGCrjygKz97ptRJFQZFAxFJeWG5zf
v4OO6inQcItTdLP0D6KA+CHh4VW6o8kp0hHjqnmLNEwrIw0du6PJbttgtO5+oU0rp8Avg9AOFHzX
9Ame25ssVWNjMCIKc6Ke4r7OiVqc5RSoXLDJAsgkDxRcXobicSdHzJrysDsuenfp37aAddSSEINX
MvrMuR4MRollzUHM18u+cTjsoa/pWs/NTiD5LE7X25fXp2c/tyTuwBNRX9xq4iw5xiGhYhECB/uo
aYaT7HJnXn/mZY8dX1ct/86b6Ze70lEPTKf+jUumBvRVeewMuYeZePnBsw9IBjx0zEo0wcVwdwQC
ItwCtWC3+t52RRDgNVOz/JjuDsfNMIUzHry1Q7iUsiNcS6ea8DA44SDcT5keUJwzcshW8zgR1XtK
exi9KyofrB+Lo1ry2A8NCORZJAmr/+xEcRsfRfxuYIfJrO6H/cR1EsGeCjj5n/VzTMvlAVr5Fcjt
aab77+p0jS8Ty1MCv9NYgYC1dc54msayc8MscVUwr2a3UzQe0KqbmvbM4X/3sFyIUeaQhdWy0CLJ
PyT/nfbzLxt8licUBnO1LAVVH3nbSQ4aB8uxVe6sKHjO6P2jMaIcS0c8DxIUZIfDTsuMXl7mL/88
TkKdRSVhJ1mJYJao5Bm9upeRIcztNUkj2imkYXgBz9AficB7YgtSy4oyJiBszWbgCm+qKxyN9Bj2
ZyreRizwlJ8kpeUq0DELDmTAwe4tMsLsn9E15/QxRa7OTZlUuTc232kUDvi2p66K6eVBZtdU5Pmw
rcLmoWqgog/viysrDDoWg5Y+pKXVwNJ/Bf26BRvueEqHXBHeMXJxxuNp+562QwXvW/420suhvl/d
OtEEy0E5JfzyDCng9SZDIVSPRh3PD6ur/E7Kr7FujpYO2XkIdTTSpGuj1eFSAkwXVrBYMt7WXll3
sx5t/nSQ1yQDzQe7PjN9vF8UOOG/RjWHqcz/ATQT0wN1y1yPWnRDFrF+H6a/StCetBKC/WB1h0Fp
ZnA385JsZYFqRITsyBYNpmZid/0h3zRPhcI5aKLcHAasgeCJ869R9W3JfVwN0+ejcUZgiRn1guMt
FAGEF7r0l4OitTo4xBg69xorht98//cXgZWFlW+jZPY1JCrh5+w2J5MdEgf95ox8UItgIyXjC8yv
uE8Z6P6EzpNPWRaiL9TeYpuCMI3b7b6YVOW2RhvjQiuvQ3FwvKesA58IBta0/mLvaJzOLNbKy6Zz
rBYCuZUfQExW0Rwq1ORffmrpYuzg0M/+tUuLGfZ2nSIpHoLyNMKm2t/yOC3qWlvK2vIN+L9P21wK
s4hXRLKxpg5HDPE4WGffwMd5GEg1fz8bfSfOsizCJ6+5sQw1JALW8SZCAS6wW7KiobxeVuS2pJ3t
+SKjM2Q67XK8YTaFbMElbq1scByW2P+/w/nh3fTWFx7R6PKn/tP4BaYjJedwGGMBMTvmVG6uCS7a
R64B6BMezUibKVVmeqS4QOU+vkdhMkUT5DLMR9DPV1CV8/bwTqxQHXrO6XDdxdnHiYrdhP5WKDxf
olQBcehxfmyR48Rmyq27XEl/UkowJoFeFLSkKcIWnbCRkT7XsLL9NV56DoHmCw1FWFh37/Pkockf
g1lfKhWmLA2LwrDrvK/DEGmpE6uNhPxNend2ghWVOG/AC3uZpYckAkY65aj5J4S6VvscKM9XLHoQ
xm48enfkTuAfd+DwuD+h7VvRb0XfvgFf8isCh9zhnNRyegwnyMro5HO0Qtmg59sdocte71c88xTI
FaIJbUgdZqibvqwzO7DC4kLRLdF4cEXNuYmSd5eiUJg8hKbeyiH+9U4tNCwRgV162LZSZvawj6Uc
HtWHwpO0hhNVsO1o+Z2ZUoQLxN+LrkwLvGKBGnikSbCD2ruc/w13WGaZLXZ+vwkXOe8TvXfVie/1
0QsBaSk7CLo/LFPhsg5RQGnD1aabPv0Xc8lz2cIcfVesYUmmUZI3Yt/0ddalw50bAY4Z/kl40oLf
VkdIM3HWSbSuAF+Tn0qLzA49ow21ibrXhw63DL9TVbpb5kkCRs0mQSqLUYFF4WKumHUROE/q/hz2
aiRjs12o+fnkop21M8XkZrlGGxd9klgzy4GP/1QvjvQijsCdnvrGGqeUBKjoGBPzUangZ0zWlPnI
H0qBSl/UnuiGJwq154Xkcb7B0LHdDhJ9MyigvVGSv/pB/zCrfh7zlDxyW6st0J5Hs9JCaufy9ZKN
wgqau1kh3Xsd+3gX7/9UfWnBl7nacs8SGnZ+AO4+mtl0yFrOBGrF06R0mhTD+S7OcXZ7d7erHr19
/ZCj7MTDSJa1Ey2LAaQUv1vgBKoo2jFWLG0IaRAfJOq1+NllZ87KADKbqTaMVQN0efgAc/sMaufs
s12cygMZ5lymS6RXsrE+Gf1gKPZOmgsfK+XJodhF2ZNJ2QyhiIeYJiAafZ4Fg2zqdmB5z2iIwqQi
DnAc6I9Y+AMmaFhvnNSfVU7zCM+Zd9YUAwmKXW3HpPAaqeO56eiJdasU4xia54RPUQmFE2AQKOlE
d55O4QW+F4SLuu6GZeTYFebXTdJf1FhLt2yywaqvrJ7eW3QJZ8zsDfxbNGUAf8FEBCGL7aBFFka1
h2MvtvXG8xHfj2Mh9Dz0j3Ai/8vx/ZHEwXAs2YsBlzjq9L5Y+UIaQJvZAevx+xg152r0+FFurzNY
AYSMb+mz+KlUi2XZT9M/6ujamhc0o2b3HsWhvgQdqz3AN5X7a+BREWzCMebQTUk8RaaZ4UZtsAWB
ZzeIRHgX+vGGRwdxFJ7nj6Vudlfq1OX+NKKE5vD30Y4jAaLY98n4KZeAUKOeAMZ0EaMNAWPdrTRI
Rvgji+J8CItCZJtkCJfJJdzwa+/IpyqcuQ5VvOkXLkFKwX6kyYr+Mv/FqCGhbRvrYAZJ45z1tPG/
f7YnGXyWLoZUPKlS73uOXSdISN0y9MtEaPUlNSOJs9i7oApPrrDMV4ypddlcvW4ZzdWTWg0uKCcN
m3f/lfLKVZBK5c3uqt+7LUGx5JX83bNIwwr/KNtKa8y5uH4GHoeNgxFGwEWfm2L4UODnG49ADN6o
kbfSuM6/yWAfPydcBPRSKyVnQA3eZjc6JEkWzz7kUZVO6ZcAtL7Z3/krbIOsT4EYgjJfOP4UVOPi
oXFgBZUZuRsxU3i0AJoPbafV4x/Ygf0hdpYN8kj91STr8lAmKA1PD9FlRWs/J/aR8qOgumvBCYL6
0W04t+HvZGxNfdltLA9QPgJLUvdyxhQrGMjuXRx5/PfDDrJcabCKy9r7FgHJlYQ4pEMWYcuXQzPM
9fUPYlAVt/fhX2B25ogZJeALOMc05A0Ra9xEFcWgAvPE12DytK1cfIf3JIRzHgEHHQOt30mtjIH2
j9+T6akYjwd+u25yoQVPXl1+D5Z4ETUS9z1D7a3ZoHwX/MlgIrjdp6aku7QHbiTnvXcZnFWoy5h3
EkiaTyEje2f4v25dPUK3VJGoss5c1IW346lZoQ5ZT0z/hRvpoQwPVE9m2dDD4/Xf0E9lesGlaVsG
TnJVzPbQuwR7OPpSq88zspOWCfJnpPmscvk7FjupPn0RRipNvnYpIExXEXO/OrsfwVw6J0n59rug
toWqbWf0b/reVYIwUWamt+raC7v5mqwPwZ3uVYbI+ReZhttoXHQ0ArVysGZ1LmJ00EaOITzAVhtz
s2VFscbIplmzWGWzvo411+1eCLrPK5v+iu04ZPS1FrQJH61bLa/CmaleyWqUrcjt32TTrntDpHJ/
zwmuRWNjbf8iV9V6KI9c5BQoHvZ6TMWV0R5n6VgdOPEjWH8V4kGFIAnfJpoMnD3JKzNcWpfXTqvK
T6B4bxwux9ffmbMXKdrIoNadW9h4cLTKWwaLXyjkWX26r4rA6Pqlm4xMHfK4JTT5K1kRZrNJAMdv
FoSvnAjuPlP+zzgdB5XKIYFqyTWlZEDxG++YnfyDjJZAfyBZ0FD1oP2FBsJVyDUACkrBuV2S4CF9
LtSwUACEeo/4Uk1fCYL/hm6Y+jotRxM1cAOKNKczwKPY8FTUiX66EHQ6IhESMuKGBZ5Ss1CT+iji
2d86fAY4xCwY0D1uR3xUb9jR2GfSl9z24SQiKVd2zoDgkPxYkA1L6n2UbWYLyrEfwElrO7lbhiNS
MY8Z8bbMfKraycTc68CuDks58CKA7dZ9/b1AEzHkuMISjaPdqAHYRttQ3h3xmXD6muR0T0z0DS4d
KqgIZKGHnq8U15v6OWANFGCMFYdSW9YOGlx6o0ao7Fw5JCXKl24kmKLQrPtjIuDRJCb7r110QKOo
1fQyaV5DMAgYJ5EE85MGQjpJwtWuPqZIeRm2SCmp2Z8LuagKpIXGuntiFnbHO9mJ8W2jSQwYe71R
ELxLMb/i0+r/u5doC4Jbp9BslvYIYIcz5i/oMU7DCGH1CRuDAQnR7pzhWw1NRr2xhdn4rsfpGncr
Z6slU3cenxZB7+akZpvCEUS274DzneVgQaisqjiyQ8VUNL/j0Y8P9lcgH7CIcfGQ8wydLu27cHyZ
HyoFeUfTEIeVMPm00PDx4nT8DnV0etS12UseEQdpMGs5U27Jd0q49inuCUHAyMH+tJafcdjn/v4g
m4I2XuCb43R0PEH+SeEJHRbhHoPZLQeWGXUnK5XvSTCqRn+zRsSl3jpxV417VUZrNqKDNpYLG1so
qULDRGFQXXtPn0LGvHA7pi69aI5c0HEHsIJPS9eK40/jlF5mcx2hdTjrst1eJNJiZ7q0CmrbIC6n
iPXRGWSYYA4SykLXC8EKvIJResIN1IODxia9eUMjqUKFvzG1CqCuYuCDmfao+sMcY5bleF2phb47
7WTPFmZs+dOuN4/+5sVxH1+KjFHdRgxIVCXTD5I/k76I6FFPsIZuGxAO/eSNWwL5+jKaEcAEybFU
FXc/pV0P+B6kiFu80heUaZ/nrp65ZgaEDjwq5gr0/gTFMdU5dol12i8q4QIYPUoLzT+K2crrKLYG
3uJ0YFNN0fstPnSzzd5BUuVVFVZtlM+r9jN9aU5ijOf4OY7EA1j0RJWyngtOvCRLaX5r4CvlDvPu
nnTooCMDZiewyQhrggMOHRbAAnihEjVZ8tQkqghG4LDFyUUCxXguVrRNCCOWw8yKt0NkJfT9Uxv1
MBQOP9x0LgxvBb2u66+pGtZZX2tdfd/NtNU69CSkxxW/UpnW+BFwJxNUseaUze428KGg12UTiMfG
C9Gwsh5xuKIo/GwEBuN2XJdcTYHt9kvJ4F7ViyefD174kJJl+7ognJrmlAsWx1mVdGUcfw2J7jjQ
1SVn10cRJKJUehEIkz8h4Kv6iuRQcAPgH++qja19GEM3oMmcEvm4Y1szUrp48v90Vi5jtXCbMZps
RvQ29nyeymQDTDpUTzyhApvqF0uBjbwuSaE6VWKpnFDokT5GyG5FFNrqIXpNdbzd5CVQgWhrR/cq
X52pAVwK6YfzRQN8ruPi2D63G3jzoWXGHV8oxTAqZ746WccjHteiozcQ4fEecO0TdATjRPCyJGE/
zs+FS+n5DJnnQuvW4uIAwogO3eYTg6/oRuRDi/SVFoK9j/obdf/gh34o1deHLWydcTpMYVA8zXm6
u2CawA5KncVYEIiyXAbiNZWcyZHv83A701RncN40J7cW+7zbbCyArPTUPT03nLcK1w3D8evtBNvy
wIbqkvtx0tE1bb+MLs1V8rwOWoxDEQWvJfX0gwyDWUHmMuCehV/wwU4v18Aq72Vvffmmho2tl9+1
ScjEAAU7GcBVt9+J96ffEcNDumwm6RaStm1D+1WNIH/EWk2Hy43zFy2zGR7P/eFkOINnMmAKUHac
5zfXSPGf099AvJe93wCMmt2c9z9jpSWkv4C89lDqsjT4maH78SSoBHXnbcielioBETfFNyipkuvy
jpGtzE9rcOPzqwJ/EfpxHjzRWfxO/OtsFYgUWjM6IDkUJtWrAI+HFYFlPvQCWVeCz/Oq3zR3cjJk
eBgqCPLjWwWgFY3QjXDQkyajWxlAjTswYsoeuXQXD2E8TN2ftaX6LZL7E346eVQi/z0TmYK9oedm
qjIfPZvxTexF+/v3k8VCCXrZdT74cy3efGdoIs1JmC893WHFlILnsLUrozt+u0K//fxppCHE7cBZ
PTTr9oKBcs3FplR9ld8DdcpXauBXQ5HrNaLlSafYDekojXqMpH/1f/8OFt8xMI7Dx5qtWDuiuDxW
yf8TU/NDuwSVVoh/LhcRK4gex6hkTdLj0onX45B3qFNVvoUwfgUK1Ir4S+CS+ZYyenSMKhGZHA+v
VYWLk8oyMDBANYH+fMeuweEzGZbyiHOWWkU4/k4kTyxFSs9Yb7Ap4brbbOAnGprlAW9mWwGtdJSy
uWISR6/SWx+XmIfs+NWgxZLbh4Mkz5p8aY6TNo+mR4/U0pyy95GT3ni6PnVTvslroKTrH+MRyV5n
uNJ5ZH3fwpveBZV6puRmB3/Z6IXH9gwcydJhE6byNMLSVEX8TtAd89DAetX2CAGNlEQiwvoGmXDr
XMVME9BfvS5BC00rsr3q41+W0OVP7nsrT+Q2qf6ToZez8WIR/0wvm9zKIlDPgbsvm7bQBUTbEI0b
fLp+VXEXgbebSpQHloQAO98gKHYXjypln3lJGgSg87nWgvry71kwpUWzC7Qvu2HwXxbGpoh5Tr9O
PmG2GWmyhCEp69sraFSVK1Hu+GMrGaGeqte03lb7qMy5CYHAF+TgUk8SePArgwLVXrFwVChjt0vP
AieG0AzqK3op7Lve6wtV2OgHd+w/YFoMzYTFuJaWp+ciV5FG2KFgfjfODF9pXEwW/T5xIFULEzEF
mlfnYhte2mWRt+RPuAP3IYpVAjB6IQiZQkDowZo7FXLbwvdD7h/QUg/ehD6zQiPn8QFF0o49xsjv
nljWHpa04iz6x0FXqz5Z5+SjziD3iOV09921Xh8qW+UGKw+nIUM40NqJfd1RJFOw+0z9vm7tjxU0
aMVVYt7UCYqfcdvDSWpaFblH6Fef6oc+oJ4x2aI0wlRWiWJnsraUQOkI21IgCb8kcHBDvneMcJo6
sqNSZMxZ8ouJpAoTrTghzIdPA9hwqBp030e+dOQUkC3NQ+XSsNX4lHILuQv+WZkm0QS/29wUIVtQ
uHacHFUAhmMq4TlK+olDPCpTfkRfrD1nqi9s1ps3GnatuYHS9ZTKr/wdR1p/lrP5QvpceQM7sT9L
kJEahG94amUB0lLRyq7cea2/WeoAGpWQUGs8gEqw+AWnAQici8zuY3cPsXwA/dsdj34cMxIUIGpk
UJvp5xVfP/o5lefenGjiibceYEul3x1PFN7BhA6xtcCivvGhmW4jOrjICYtILmmNfvauDGwHyzFm
LyHNiVNSAFuPVgc37wtyYFewPdjT9wqvc55+xjnR/zPNXh0K4z1tt9hHxam/XDU4KzBf/+wXginN
44ZILGXFXE7P3EXrPa1row/r0HbWr0nGXqjJ6VUfAVl8mhlBmGCzVglbN78TKOijhWNlAKDo5B3R
uSN6Pe6tLoXHhPlNM6+YaScN0VPykatemXEVgWKvMbIdyBH5IbyE7Z0vS9zPDwZ2itLc8Xud3Uqf
AfZj7QZIYBAP4YoaBKle63paJaVSKSpoxXe3W/CCewvN1EuH5tqzP+2vZP4Z1eb0TTWpau3e4eu3
vgvSErpvEGzy6UKqzHrm5XyAc+ScTD+tu1wlm6t3OrivMcjZXSbaEDP4HK7FhPqxfg49ZPhlz8aC
hiUHpR9UVPKKITRdV+jd/9peeoY+kP3eXzLTuGWPro61XpWMj4EZ+JEDFFPEsMGxkwXz3Vtwr+Oy
MO7aOwRr1qvb9s3zvQRKeL+juzCwDhPCGYgt08m3LwhwFZmM4wIz3YuVjLUEQoR/KfvZ3/R0n4Jk
vjyEbPvbJORrEg1Wh0PFqyDnaEkQCBh+RyTiSzLjD43ABuHjNGWi2BPzvmbSfEOBxhvG037n9EDF
hWb4iGork5L5uVZPiXlKtyxuusgH+FHOlwIxdxcPIxNyiDj+rd2kKXmjpauyz7/4Tbs+8fz8D+vE
bGnr+jydT6GRiQT8msnc5c2eDexUFlG9ljA1WmwZ2JggS4tM2zvsoZozELNJDXu7cP5vhmiHnNLi
W8//xdoruBO0WwzttW8rC6CY6nykSBIiWEEA6lRxEEy1E10FDy0OXkJ99SBvhocLlHUreKRCnz1K
ubiGQRwWKjRVgHtxg+sUBo5QflR6T2ETgj1DtnPy3b0Hpg7GBh5pVdzYermyVmMMa84wh7eBUnn3
sqaQBdXp5lJh6yVWpDpAeP2O4h2yNkm0eH6BTlTeJ9+qgpJRJi0hPEyQG4vUBXpio49lj/AsE2NS
mY1DAJHFbzi6zLsIwXTT6RjtWguMd7WmrrfObp817e2vxvaT55+BmWF4wfYkSmLuBKVxZVqbEuwu
k3AAYkeZy+pZ/8JPqgrdfvbHMSm+qSyaoBOxF5kHRHZQRj26AuIZJb3tllZdtCq61lWjJTLJRlrV
lCRrS6uuDIu+oLaOERMGZL68Cu87dB0KBEpQRtNhc1UgoGxJ6wz5iVfiIL3GnrtFvXvSIwxBydue
MJ43/o96MShAqfOXsltImaY2GjM5SCuZkTAk25sAamg36T/VSs8SKaLy4czh/2Ww2g6zfxZMSKQo
01ql55ItbviDDcaOY8H5zO9g6pF+xGWZJXR4i0TRxxs12uM9o5njoY6tLEfK+Dn1HnZIoJ+sWdXG
u5pz5X9l7k4eM4G6o4jByG56zQ5mnLUSR4Bq9guH4LNQPwRmREoCSXGPbx1OMd0cx6+kP7KY4qTs
CQBaDyDj/yX0GT/KU9x2rmPyLf5c+t08S/HZi6+LEqAgXS2clStlpK0FsSthOmkyc3BP9z6KLdWo
JxcyVGf8d1FnofpJD/JyKgoUjJ4dgJbeBFDyK1V7QhsuceArBOzoRfFprqjn8rqj80UCbiObP4bP
2D0vsfZKh7tsYbRPB9xeT7zk/qpF+jOxZFgphGCuupjilWPz5X+buReS6Qc9gC6t0Em8f0UKHCSm
V3d07Dap4kw5w87vn8cu0sNkT2ffS6blGgo+CSxBHmbGDMHILK6hWYz+9X2JMe/S+9SzskHHjqxU
gK51VrBb4kEtDNFFoXu7oP5fsyjJNgUVz36bkF8ZZj0ZZq1nk129mgTn1ne6SkqI6kgxMmb0UP+O
iNOoV3rabwvvOf11V343Bt0baGdh0v9APtY3riGP0pdQed61XeId4ih/NR9bvm/Lbw8fVkacugpk
iiwie0lSVRmXr1pC6eSfayvhyL5BerTaY2wzdBz57zlPhVm8Z3UWa5+h6/n7GLsPtwczJtUrArh9
1bnEVZfjkk4YQbyuf061W0lqvprQvN6nZ8Ju6XdrjtYF3t30UuaSpRQYQ/wHR4WOjT521b/4YY7g
uTfEFaQ+q8lr55zcqp/N9wyD72QNDSluT/U2Q/kRtdiWB0OYEqXGs7H6Q9/OGbUgmiQXycDcPQOf
TG4qDwHzCkaf5KuLxW2rieUs6CdY3ug9pG5ploAEEXJUxE4FXNXHuLogmvAyczSp4uF2dSomtWCB
lPxSBHQTmaOn1eLwRZv6da9iv2uJR6/Jqv7mYg6KlhZ2JUBIXvcIU5GQhiJheJprTKQRkjNU60WD
18UnMb83ECbIfmTGPPDeqXOsV425uDccx4p+0am9RHWRkXgNSN3PBSoofw0fwHof96T4VORfVjqC
9ei/DrHHkvf2xjqJoLG5UaPZL/RFpKS5jASUS0xz6BcCEaDeoLM/Z9cKS90LmCxVf+PQd11xzj5g
6NBNGnffIgr32WB3juVYQeLQGDtxNxdVtw4mWYpPh/LdClFZp8R3uWm3P+u9yEV8VLb/bJE=
`protect end_protected

