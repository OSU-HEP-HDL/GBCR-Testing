

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YWwSN+9l5ahBqN8tuQHA+pe+2Q7Fh9//dR3H5K2w3KRc2pla5S5ifvTi8Ak4V+dzPFwrZE+Uv4ZM
WqK4mWAaDw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WcjiphsvP4YifX33L+r4vrauIXRkGno8B+olsJNjoqAxagaZzNDAFnvGiJsIWLTLoEkntxsgRnIo
WVce53gFCvnJJkmdaYhg6W308/4ThcXkZ2dT7Q+TUTpvKAEe2vDwO0foHspYl4iLWX2KqDyY9jge
moxvN6KH420mg96l6zY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wvng0RPku5m5MHpJv9WwJDWJ8F5PUKDSPU7V99zR5erdP7PcyDhypTKxqOMHkizg+gEusr/QYxdH
b3OK1yRKUZ44xzg4dZxpsvitjqx51I8wGaS5oiuyKX8hGtgTVrbfoHo6u9pcLQZn9XK2J/iSrjf5
dyOg2xTIXw233HzwIrCKg5RT8dfxa+iICMhoGVZIGJ68DJPwrJbT6Swg5gWMje7MS+Ppwgv0Jxqb
7HSKZuEIyqOKVjWI9mOWG9o9+LBatVHO9cQqYlFkeCwc3YeZbVHELaty1PZ3GYbJhCtr7obXWCNH
f42iQcUXnPWhD7j92uOOj9mnGCfQwEtmFpOg0A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mnRNLVCxq+sgQJhai+B5fZRsJzZ93rdvyaCrmwTY5fIgoqSgRC5N+TQCYgevu6oU/nSzurf6krRP
lHQ0Ztrjgg2Tj4+uhFcaWXWp3gef6Qsz8XcVJ4aB4xMaBhgkUeweDC7vzOKD05WXxyBd0/qZdLtt
lS8j7xW/2WXeJFqpGaMZ30TpyNYKEPbTG0s7zfxCOI79Vadm9yVGLdGkntvGV8guzxeaRo2Qkmsm
e1+jXsDbdOr2euBE7JiOnNqartejTWUhtjRbkQnS4YCtUcNrW9+ObOoPjivEDKhArV2d5T5dFhZd
vZIU/RR6j3BExhd071LKzolsdnCqR62C9tEZ5A==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E6549NUXinEnqZcngO+xA/zs1xe2Bus1VEuxweH9iD+10PgNtRJtsG9EF7ZdZas4DjOhgJh7DHf8
ndbSlKTeJx/4QdIH6iyjSx9xrJbjCC8TeQlSsBzTcSKNDMh3HuElLUknuM+x5+UC+hkdrw0waGjh
tjj70YkP+K8Te1Nhfp5PHo+OirttOLZY7Bnhq7x3KDxVSyWnLuCBlLcRqRosb6oaQVAF5dnEKVG3
DDqNFX/V0KONWbfs5QSo5gM8f237iV+nwxPmst+L5casdH0vfnMagphcYI2Gs12f9zJ/qipttgTQ
46Pj/rGC5IRv5Z5f3c9wnJBWRVPQ0uHojBicwg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ogp/UkagRFxN6D0Tvatf3PJ+RNRc6aGWLVAuekDtCdp1urxgWDpgdUpLAqv4gVFTloxR/WYTIPAy
tqnoQwfvxF8+1H1sANWUqIMweNpcUZzEYS0M2VRPa5yH9GDRSd+LmMbbrq6RbwvXiR0tPlJ+qF//
xXzjGxQQlbn5MtTPwO8=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WS3NnUM3tGvHLrK1+gyTpPfI4oWwTOYDJPYfQBcc9ol/GaO7Z5AyMRqRkk+WEY00WrbCfviFYMzU
pGl2IHT4VRRzqqLR91kr2OFbN6OGXGirK/a2SoQqoRH7NbdhMzwc2r2DD8mzssXGs2HnjNYorDiE
Vs1axIRZ0Xwgll0Xql9UnW3+H+bZdCSjNWd63t2LxcoNPpatkn50Aa0uZrOTFNGicGTTryERIIjE
tD/W23CkHq3rM2LwJimtfOkZfT6H17TZIlmdf4GzYYEZqzxs/jkYFtiD89KMP+/WhCVPGWSzHT/R
ZumbUYGnUPG9wSLIU2c4b/c9CXNngT5yj0uIjA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
of5vMGwv3KZw4NIytIvgNKCXm920VXPicMue1c44JJzZuv8ST/ZZb0lgDktB0M8qEwCiGhF/dYrD
U+5ofKHjXydnY4lnoYPK43lMwrtoQ/UXeT80W+2FUyJ+WW5DI4a8LpLPX4EwG+iVTk8Fdcr8SAfy
wJ4fgf6HwoTQQ1vinh6PI/C9XQYs8wpPNoY/z+EnhH2WwvKNl4pGnlyy979fDxyexgnVQoPhhpFI
cnSsYGanfhHPoYMJ0qSo5m5sC0lbhvFFT5EQNFGfwNRtXvGO4wyDuzccvD6skSp0SKG50g6sfmcf
MUTdcrfyRDs1nEl4Q1140ynz67OeUEu6iqfEQ0qifNblNr2fUqRt7wAITr3u9vCjNWEkW974dIHM
QYsSglcq0y1Xw2BAsDJU0swyisK6t2U86sRugQNwnzFl9EE0SQ0/vRx4/eAzEZ24PVKLEKeGfseX
/K0OTMWUzXnYf55yUyDX+zHc6HABAqq+orhgVFa9arx1nb+Ie+GYG5gkMzlybg7XJkwGx+48NxVC
cvb9xQOnKlj71YME/ejyOOaL38Z75m2VqAnFGZw6EI14DGmLikLbZaoRw9KkierkBIWsxjnQUk38
k8s5THSUhTQ9z9VpvVeLxeWn9VkR96mVs9wytgtIGr5dEzCYbzRvBEE0Muc+6Tn6u+GH2oeMJbhL
yrzma4V8fEiKknAsYIFKiWKJa+FJXd7ewMJ/gM09bifuDzaPmyydJlL31pIoPs/feb+emINQvjw/
WxI0T0lTqONkpgXyn5bJfFZEUv+FdXcCgEtYEJ9FsaEYa+nqyr88/HVOvRmaY/GVPSlnGagdS2T0
WHGsts9vurUe2tYiF0jw104A8UT0vcx3/+vwEQi7tNMl4GGGLZijtTzqcRHnR6cBjyV/+VD3X5Av
xaVGNJn+SpHQlyTm53e55r9QTrEFlozGq0I7w+7lqaG5pdRTsTMPO0qjSvcRBQbnIwKg9f4DjYOp
k3jPe9FbSPMpxHRypMIz5JrtVuqxXGFrxFuYy0QRz7ACEv+JRmYXxUAvgB5WuUPrS2ReLqePGNq7
HzijCHORFOjRfy5BEM0LSqh2QmMu/hOeTlOCRFvteOXVwQ8b+4wT8jHOmkk49ffwLmRRdI0jYYgU
whq/ZM33eduH/H1F8KZQBWh4v0vrOp+9EnM11qMX+u8AVGCFrce1kUFgO58lszLm6AA/xScGMrvp
ksq989+zvZFvBrCoDTbc5FJsLVAMeS1pD3jSoj6GMS/FM7DQ3p9vgVcWAJ1XwfTTuqDLS8pHEqkw
y5DYk1LVBAOPM0j3yzMoaJapqVmIWl8WfsGNNJHs28Czds6eCzjmhFGWivBUX6mR9SKryctHYn5m
jtGI1euk6YdoU56BPCAejfYJUUIcIDIrWHxWni6Du/NyGtHPCrPsydWfd3ijZnAl4nFXhzX02I1a
hi31gtQQsN6soGYSqAo/n0LrfSKgjWiQNPPHNSh07+p9DRDMUwGHUK1rCnwUogcpu8VKhSSS/Hio
y+KdihIbmesH8SPTXWkggOXTR+dbPTzuonBjjEt5Of+M1y79Rktgw7PN82FTs6dKACrfV/pDCg6j
23QBd3H2xY1/9Z3J7Et0d/sgXuYwA4WDS+THjU06vcXjY1pOU+SWRVZ46APJi+8rwTqGXC/OlFnj
KboP26IkN0I643XWvIV4s9+IwLy3uC3SaL5/0mFx5nAXJoS+7sDwXIWt+/1Wo14dQFmQIfxefLzR
/mVVvxfQ8BttecxieL+FRsz0DfpS1uvD89J3b4sE6MA3wop2PXIfMxwAhVNB06NI7gDlTTcupD1v
LIg+M6LSPzyUcEKCu+Eg9VzxjjP8lYCJdO9bacFdvsyBYP60N0RxADgihGoel/kdMLLDe3Wg3E8q
lR62kBEsnzZmeFDE4GsxKhigsoYGYYSrk3hSqGaHkjeW+/9PMattwpKOeSJPHmc5MVK63staIncn
jpW7splr9o/DJiARXXjVXKgU2GseyBsJd5OYCHNKIFnAsBStFjklrqvLiLXBzhyaUx30iTv49Upl
0k753lT5HQnttOk6zWoImME5wPJ+FKBfNajrPRrXZDSPdycsKE/eDUCeunfzFWo1W7ThKb42J98N
QAPRkyD/4DvIsnL1icziad6e0jJVqB74ABJSq+Sjq+U5PR70mMOAhukevZSaj+kZEXXwOhMEHxB/
OUAKdsP0eCsMmsAtvYdr2iVEAmwwX1U6dlGEQX0BVVURZnZLCqd2ktx36Y7HmvKGCNR+f89ulXmr
fx3Ye4hP8D4+qbYHXiSiujKIYV8JVZudch2i1Dy2BY67RBCyNuJooopovetMWbeDm3OUH/FzrbHK
Fwze8YwwtLgsTQqJPoH7sTB3OFO0VdolpfNIzojYqZT749uTNgFoQ6AnUt2bMt7DptbfhmcIUli1
qiQ0nUkIkUQLe6u5LPzY4pqOl620jI+sdK2nvBTB84iOmXjoXpX7jFGq5uywAQgEFKXHigwEiBXs
bnziBWRzhC0vDg0YkO7/TwYqwPmJjHrYrEY7EGn9oZlQj5TB0AQKMohi7ibEZYgPM6Z32fqMQtHN
QRuCmALoPHYiaiZSg2DU7kSk1GLZjOW3OpVnAoXWSdVDFcYpMYh665rZRJK/0ETsGYJXINaCtxhN
UMyuWz3RjoKup7ONP/LtKeeuv6P5ply6FQHiZFuytybBsvrDqPVrikp4NBOhkWneAbhvDAyvv5vr
8H66+LJZB1+Eq7MV2MwXGajpPbSCtBqWloksnJNomhBBBZw7g9hG1ItG0+dqUanwzVBvk9unJj6V
3bOyXSeLgft6q1k/XjHooKQsC3/y1FF/574YSSBKRxNO5vWeS/eRB4IdX5kYhFUgN5BUdrKQZH9b
Gfj4MrVKsTjy9IQKbI3Udlzy1LCIYWWK1Xb+Ly0YnPpSS9pUBmmjuxcNH+hG7jvwAIVHr9s4u76R
4tXR9DfhFC/M/JxzlytewVMMkCoYNHxMbR+wXsNITZKvGx/WRXMlAwdZiDtpBd+1nXerACLxrhaJ
qcET0XA3nO+xi+Ct0jBNg2tN1j1MBpCLWc88y4FcacGqSVLnSvEei/oG4vs+Mu04x8tChwP1M/DW
ScFSyZSPlyy3W9hf1/5GD1oD06svVypHI09Qbc9ftkUcc8ywzfI7JzXVWjiF8xTrzUlGYm1YbwRJ
8xfy+yLwxGRoc5JuaYUh4dAk8J1kTtKv1zQ0nZ2nq9ldLFXg65soqjBobuxldxrfy6933Wi5DZKt
iN67pypb5dap40rE34EQdgNfiiuaiOq4Ga2E4qJI35EtP9Y0Jeuyx5/ycO0u4N0DuzbqUk7pfitr
r1ZvY9o12j1ViVq89tP6dpHS4M83rWEUOwi1wuE1x+TH+PtPcVFJztkFHoKKcudvSu7vWO8WFqli
B8qox7MiwpgtGF4rDY6a7YilKwA1Kvb4YDyV2U+KzFr1htG+ZsTA6Z0wPbY1pSq5dO7Vp+/8YOeV
NWA2SICB/g5t3XGe/5kR5uwwmBkAfZJ6mX1hzQXJLyFWxZjoN9pm3Gt4V00Q3Rsww79Oj5CwMaSF
TiHrCLQnPInLW+p0gRYOCqcgFqCKmCtCRUrV+WYYdUULHReV+vw6mraxSW1uAeEQ57xVJ1iMUHzY
MsOW4YJg+PiBl09a6s3U8cpzhzywaJyBVXPftg4T621WYn3PT1T8/X0SSM+j7r0JHBYZVhK5R/tq
myf9ziZZsBAEpNrraO7c6RzPwWM0C2IhxTeDjPOFnY4PWOI/UsD+QbIECAuammW0eYKeaDTa/X0y
yMZTsCOncKF1DaDAwINu+JErJjbCVCFQvDYYXRcwEV+2CdSPu4zUjLAR7SrcQeJdt/vTv7+uTlGv
sM1dMSL24ZIEYdNxIkSxIGH/OivTmqZs+YaawshcR0NEvQI+l2aBN1lsjW9Leg5L/BdpN3AvVFxM
JskKefa7uLGFkhLLaNKQUggTlBi+nTZhejpCsmLtrfDy5enWnxiGfYFJnjuxqRuxViTnEU2tZjb4
SQ7JbylJ5lYJpcA1lxXNX3GaE83uAeUvWOB7u4xHgoT1eJ41sMoWVH+fAWfGp6Gos7yzxX+Rt2U3
g1G6HtC/LOZjCoEOZ5Um/iw5RiKBSNEzmT1MBjAoWTLTHmUxm6hDnxfJRjs6SJCbqcmWT105ew/5
sOYKxtqmmTe1r8S8s9h51+4mfdxh0I1rdGSmZALX102UD+idYjXcfpuyp/GI7wZenf6JMe+BDxu5
KOGS79DNNSWlVU7d6FUTSF1EyYkpIt2bilxKbJcvo8eb9tSJ93dbTbSUVK/Abpvp/+0tjsxUS26H
bww/kV+saVuMl3eADc8aXBnmdT4X4860YdzYP5QBZPLV7zghfQoxcHGhdvBqlqL1ZUX+B4q9K/94
ftSdFWLOqwKcNTpfZ9kdkG+6MpEm6FUyB4dVxeHWiktEqyHwiOZvwmFfyQqfQK7uQ1W6azn63Lvf
5u/U4hXjfnuv3D0xPZ7l2PrpYkrNnFMI8/HU7mGLhS+1bfBDQjf4PVQYTtxH9njA4e515TR3cbih
cB8OhAylxbJeSsXC6/uGDckohZn8OYhAT69/ArJKrhcZsRJChDcMXbRoctmKb4ptGjaYKR8f8h+w
Dj1krVVNMwsdFgRbyHbpByr/wt22CWX71Py3M47AqxgaHCFWbpSUWe/hC1pKKml652uypJQjGUij
LyixQTb8FbGuqE79qcukQuppR4bByOpJK0C9jTl8CDKdH22jb5Rvz2cRlR8H6TlfH4qaiin1HmyJ
cpyqjoQC4nuoaHcK8CYn47VW7KCxrAoOF1GL9nt5HKUxAlI814/9eX6H0LUrgFpon/Rw++61+ZBa
Ecv5MPKj5MMrqTibhlrHmEL4F5ccynWL3Xd1Wb6h1TAu4C8VHE53Zwyu0z/S269lZVRXmLlg2OVL
F3UrmUMPzi4XboALcm7R1haFw0JzW3sRmPeqsdSS+vE/+FD92Fa/zX1cQa77q+4Z5FzlRaBNjPzU
J3vWbvKravlc274PvIntVPN1NFceb4FO1s3sG0KncLlTv8MJsBdWHHcRWsT+YGtBYXJbkYUDssqm
XBulHOXvYj+tVhpvHciq+SKvZXzW+7zBQ/TJ3lV7w/TH4Zb7QXbQ1D11TjGQRPs/AxSHyeEuxf3t
E+5yBwMCEOCEYnxGVL/PNcP93Zp4Tx7cf9r5FF6UZSjppUvxhUS0rumYsW7GdhuPoIWYrTVELQ8D
aSAYdaOdmu80sTRUPDLoPao0QeIce/3U5V7ZZSousydGOyXxm68lL252v4HJV9d6vo7oXD49z3Gu
MxZ1OsR9+v+xIL/LiXHCNh8F0DZovyKtCNTesfcwX7SI5Dc/nQamZ4GXLNxG3xkxuhFdAtYUVkos
4FfATYlYLKrsLVxHh5uNXfvJcscYWUn9dEfOuq4ua265uHfb7OH6t5g4ctJK5M7o72ghDs9mGqe3
itXCBwgFN0e52GI4pHn1aUD2feFM17NTuT6ZpeGjwQODdSJTkli1EBGa9Rn9U68jd7WfYObEFBE/
eqM2AGGiYDgftnKna/1aYc5rVR/syeEmgkdXbY/5X+dAEuDBfjN3Suron2amJjM81z67V8tn3o1m
dx7LlcNNZ+4YnmLnoRr1CVuxu3xss2EkSXiLS8eH8S3oyHedWKsth5/KwUNCO3TZ6TWawxxXdLfa
ZzCEdkTLgRo7JyoKR/fHNl2BbWz0KX5FYQJv9u4g52YglD6cmQqUfTKbNrosJlWxqJADgiwQQY5c
22muNMbcDwhf6nZU+aR0uTK5wEGKM3wpLWKDTrhZGjWCAbM0NYzRNrFrO4bQbH94esuD5pcVxaMx
Pc/moKg1NHx2zlvzOJiKlmvWCaJW+TaxJrVacFmYlxLoea2qzFjUPhEaRmi0QWBCchQrfhVVAFYA
Spp04cP++75X9DG6Dj22/T0j8kHwQ/iDFPWODyNUzjBj4jELqS1hiwlYfB9dQH/0TkEQ3NNdJVfK
jTCk3yHySXnjm8t3T2cQAakm20EkhyAIghBsofPyqJtPE9TWaGSdF8cqqhxvvlwxUzD4fkL3HFXL
bcyxN+jLiV30ERLtWUUM+ZgdljexqSpqBnlRtBRimyBeRHX4s7zKq9tW9/Y2iUouXGKX40e6ySwY
9oEbUKH0SJbPAJMy48R1U4xvm/OCZZM1NdrYyiOFKzr3dbC360EyK8p6qJkwsOUIJ6biAtCiASVe
DioV2lHZMLujurBOcOSca3lO2VA6iptcwE+G7nz+zKG/YH8pdH0xZS6IdS1Id+l5aL2qVe5SuIK1
P2y2vnsZO1tpfwnHWzGFcvfHRTFqIbDeuVFzdLTaK9LFD/sfOTT38AIdaNtwpcakmppbq6Gk+Ttf
DqTUFTvtp8SO1bkPNQ7F+8j8pNpE11jrVOKAKaDGJ9hPKWVh7GD69aUTP/mG+RUfxBtu6Qie02T9
5WYe3y84yMIGbt+EiQ6UXcu0581oON5tTHrcCmw7JQLt99UcacYGy60Eoji+JBLHFCe+t2819Cc6
9NfjzGGcNUfgdcl8/A5464B82u/3BcKDxxue4md6+hMIC31zi7fXmC9W0RzHEHrp5n4PVAyZVP3R
EH5LN6JWEkjnQmZtN0ogUUguGyuRttFAH/KQ3bWigc64NygPWk67ro3qF7I9F12rLkCbluvnbYcz
obajAETCQe4NPpGZaY1FQleonkfK7TKQIzu4BktKcTk+Y1qxXLoyA7WD7ym7XHA69x9j3mYc05zi
/kzjDZP6GjrKV7UJyCcy15RdXKMNXjjbnev1cdyk06cL95d8neGAPytK6vU7onUNyxwcx0ku/bFF
IjwEuiPzuucKmGCMNaQ394zmrm5x4dj1AiJHG0K/cfm+AcxcGqHRkUf5d5LD5VGs1i5RFOY34/dF
MooGriTHGwMv0Lhui6sd6z5mo+w1iwPocZ1W5h3k/SLhMCCdtOq41/DlUDmYvJc7E356mTmAKMEZ
PX6KMEM2AYNFIhq3KCaRIi6mDPouufn7rYa3ABxJtOPT8fprjHOf8P3Ylj077sl/9XcUxnBWtvps
v4sEQlf8ZiLcBrtaERpawpc9FkvqitOnpmvE1eyGu+K+AtZmon8cVVKxqR4meWa+cwuvcekkIqBS
TfDCcpY17cI6+Gf8LEt9Vnh7e3d2qf9Vzv2pS/c+PNtzmxqq2WOMuDtf0s0c3sbKHNkyPZ5E62Rz
Q0IOH0FL0qT/3oBgq9LCsKKF/JwEQ5uaX7TnQG0LTubMEtqcQ3t66PdlPQf8oBTwbQjeQ/c9AgrK
GTlnGecwVJKEXThnjFPAmUDsQk4FLmdoef629lhHqRDFhfArFHGhg33m3Ujopl7hj0rm6aW0Xif6
hHMQEoyMAIvG3Dqd3e+/RitTZirHp0DYnXvYgJo/NwIzKF6D5PVCr2D1eX9+xO6CFncdwPfsuiUx
cGmJz4KSNiET7EPKabmuLsfMeiPTkHY1ttrQMSI06l1YSrDjZg+IfEvDyrHpfnvxNR45ODx6kQip
TxGCB039oP9/GQ9noqHUBqOR/KgpUvj0EqLjro+Nrz7jX1Zx8iIadqZYFQuoTA6CN0NWnPfWixB+
XQvK8JO971f2F6Yf87biO9307mHfOiY312nJEnsU/4ApQG8RmPj/B8i41kkuaDEvAcnRdCnz0w5i
Yje3rKEV9iqou6e6bx33qDwC1DGFfsAS70IFvD2rL0T7dbN1F+Oqi8Scucmdh+uogvxQpSjggrFd
mBeMM2kuB1sXhlZnhrMnQ5pka591VZzDghGBPQOPkwdXVs2EqUBuwFLUecL3NGUZnvbs0EHmwod3
WfN7AbW+AdECwr4hqVYNlojTzTfbm1dVnPCadEEREot9kXBlJOz5zdewovQR02qy2JAqgZnU1uMZ
MsipeZqt9Ea9xZShWEkF7HjRg9740YDpx6exW2oeWcAO5pPIWNz6irVadou+yb+WtUZyH2lu6LhJ
j+PTSbg3bw7RkhDdI44id7tyGrbv+Qx0Jph8AYjaKrPrLtcKPWMPvy+AhwM1VH5N7RXyFoIrkfoa
z7blbt1QapmV9MSl9p4bqhjven4g5uwAWtYWa+KH7+USKc5GdiZP/hI4zbMj9aKxyNvCY/Nz/3t7
uMbTpooZsP0xLFlIX754j9yhqgehrk+2mBtMlGadAh8Iub91VC3DHjgCKMueLoQLQ7G+haTERrSO
+upBMwzlRGQnbbvWIUv2CWqkKwoAF31r300HsOWrQmBBgV6IbOacbSAW/lGmHA1rpaNKRkz+hgMp
/vBEwLgmjE6oYqUVfBS3v2pbUGr4yyU4u2ssozacXCIWm2jQiyowhT1d5A3pPp7fMNjfIPLBSDCG
Fuq2fni8GB98OcbQuyxZBR4/fiD/d/9f7WXX50inbk2jDiCvTlHX17S2FgHqpDfwygzHk/m0Z7s6
oTVRh1Gz79jES04GwY9uqoyXSbgYV4eSjEnd+4uFtqol5yf0zcWC/y2/BXg3FTwZZHfs95iBZgEP
xZykjbvPR8WlVIF2olfIQJR9YdTUPDS09Fnmuu3n/iLZU1FljxiykO0hS5rf8bYpfvzZgeyl9yCM
xyAVZd9L9JC6gxvEfOxg611tcrt+mylGpP53YBJnMNt2eTMHTYVUIA187Nklsimt0O1IhfkFwFwT
S2hABkKGue+EWemn1Y5UJAPFyFNsibxoCjup/7pem68bu+yiYL+wmJCR+CI7QD68iDaBQJj8llB2
GE9FhnZyvdVChDYtkjdncuQ+HUx38vo5p/nUbpD2ahW8BKibkfw02Q/irwDn9ZMHBelaRlAAMGm3
RPaBIL+Y1js5sbpLxu4qyNnylk4Iub5KBH4lyRhrjq1YAwfGxdAjKVbWRA9DX7wkbXxreyacc8kP
njVQzshFgeHNBXgKvoqVhN7Xmako8Zh7thhZubRVZhS3uzA1P31jLUE8CacbxEyVt9togWJ4AXK4
y2moIqXRhoEzKL9Hmfodw/kLCs5fiTMa8cZpo8Hg08IuEeSrZihnVK694UHwmP9kLNiOJNIoN4Cw
2O978xPqINZcXcSsT0kl1Rn6n/j8iRMEODxcSJJGxilGs9bg4+CDXWu4ci5pHNFWWOwxektPKmlG
Q0YZbPcoiGX7LyT6TxwzQxL6eO5sPxwBfCXEh+bBb3QXT+Er00kmK3M9sMrpMeWRte1jupKR1ys+
A3v1MoenGTsX/3kyRDWUIYOPxVQqfY6Y1K2jmmnFMzb/8E1UKYjO1dmEKSjbrqeozBp56ju4bXLA
wZ/ORnEAfPw8mSOwLy6gM3saGA1AMzLXffT/JqooCDj3J7AsPQoY4iGHcHLrJh4lpT7pPlOGtMBG
yodBvJjJQ/0gN1csOzjso/QvXrp4jRIebnzWONMw59KI6Cq4IX1iP2reETO4GCsz8z9K35QJj1N9
MxB/bDc1Pho2LRo/NLVNyP37xwaFEFyNSZ9WZ1J1Yzfiy/9jZHyHUWC77087d4RY0f2E4jj8ynK9
trbdoNLTQbyTOVgxxHzKo3Uzl/27Yazx1bFVp7mHOpXVmkdGxNtrRtyF8xIOGZXzRiVLX0sGfGqY
i+7MJ67F9u61rLM1mVoRCzhk9Rb5GW67qqw3y6km85SMO57dFoT6Cxfoy9Qk9i9CSxWJl+HYvbWK
7SJNqxBeOyRmayghL6my4AD7mXnlp+i/tBGh3MJOKiW+3Y5ZOzPpUG69gaInP2+bqwkspS0pBCek
o6S6WZLQ4fcTTWH/L+XthZN+fEL8pcBrlR/vHVhv8iFu2VSVkcWZKyz9hvYUnT8aMMQm02JiOAec
1GyY/+93WVlFEMrlUfRjQHwDO7pX+SBjZmHiSxjuBjlmfkm2uzqZNvDSUXDUX8jOUR4TERQb2eSM
hQP5XKmICFatbgHZb2E9L5yFIi6aI2jI1B/AdpeAmYbi5tax3Rc26FqNtdZ5iNZMf4fy+iN5dxfi
e7h+glNe8UrU2zqIZLm6KC/Wn1P77SQIMfuiphRf0u+/xLth4fk+m4uAVUkKEcoM+M2J6BrR0Ryo
uHb2WCSlPPhbzklpErgnKzHnpWsqekhF6KXK5p03ST+2NjGusLnOMVnVEj+EhM2ho9aAbmaWkCUd
WVroVSS0NxfIUrvAytluxxiGu8VQ41l0Ljf1jH5j/PK0DfHxw+G3eBBvNIp75eve4wRj24HXkr0h
rVQaUCW8XgyuJ86EPz8GG5saIlAB1hDekYWDDQeSkUrlv69vNGvR14MZNZ7kU12ehXT6kRANRlI0
R9wFWUB9X4tDD0OOh16jPaVAiNpNWZTjAM15sNcNNEGwLxKK7SgLdUnPg6ClCT6wXl72OxKAkTo8
kfCg1CPpafiDzHi+Tm6mtk8040siOrdIrKQNi322TT8CnoKRyumrHgTmiFo0w5JsjSiOq+OdeP3p
b6qx5BE7MgUaAfiDXdYBVIdngCAJXS+H23/FgqZYcSYSKhCR8kxkq2RvPPaGah+4oFhNuMmu3vza
mwsLMB6HeZz9bm6J7nv5DDkIPqqrh1bzKcT8Q4DtBBqlnzoqhfGPM9F+sHLF7pXqEYuwRjGTIadf
/rj1ZnVnwp4e+IpoL37iMDMfbtKLAWRq6E/doQyCe9hlQI5+mNfou77hEc55NMox0kSddbR2l5Bq
I7iHLCjNGNiJ2nlkkmskBfL5finRj1cZ7dIj8va3+wQpki+3AJ+b/YqJ+YRxJljM7i4gtKoj6Rth
n/18S+Ud0NelCKQaxQ9xLxizojddKuXtK7R7pVhbm+qn2X/iMLoJLlazoFCP8re9uW10Afw78Tcp
6KS14IAJozOItdJj+wCch9Np3O/eEMjDi2AyPFV1rNw97x9qXt4EvnUbuw8kEbSxijNSvZ5m7LFI
igXr1fUSw7LuHgvJR2cmaSBbogKyHg4NjMNWwLwpZhVVyaA5j8vLxuLaO0eKVExpTlej818TPffK
yfAsRQE2rhQmCIuI5XNGYfmGfSFUqDgK5rM5gUr0UUr0Uolp1J09fDd0CVI9gXOyaz1qOjF1xyUE
icfgb+9s+KqTOFyGeU1kTdtjXtmRH73hw7EqVA7FoS2C0T34xjKrkIagcmDd5NPTcMprWu6tO81Q
tfrmrHbk2Q21Gy6p8HZuhXei7HbXXpSO7N2yxF416ybo3J1b4VgmnfnZsknUkTlUGvBL6dgbZ7ne
oYSAATdGRJxDp2atN65rO3nOHuYB3k/BbgBRSZzSmVqAv4JzQCIy43ft8muaPDG2UZ6O4MbUNKVt
L9YifzWwPSQm4glsEnFiVGDB9IUKTvs0p5uZwPmi9HWmNODlal2PTVW2wtpkOAA/N7XCdK0lQp6f
sbqfVEuONnMkusWQazy63zdkgP7Ihi+MkY3gBJjVKwIGMVTUMnddu5iigClLeaaHi1VItCK5vJ17
tGjF9CfznBJbfXu2e7sj4C+xLfJlWaasOtUuvpT9yEiPQnZyJlLrTN1elVw3pb+YVu4jDG1p6Jd2
b1gIpDY9TzqhYXBNUChNQFsxc8wNtRtPmJWbJxn5huRqtxK+hE7PMv5MYHurr1Ol7rQVCTbvP/Io
v1WBL0u3GZ6lBF737+aXyYJf9R/TcuKMLVSaGS9xxWKK7ZEYc976BilW8meRpzpyJ6hrKhhiMCrK
PID1o0A/OESElZg/pNoH4cBZLlnMh8YnpDTwBz+8wgdePiAazU3JyRXhsB/FFQLMJcSMaD2fa7IP
TNgkJnvzHWxPN6uf23S3p3bEW1ZI9VFcAUjULt/UXpjmWOWYs7IKJO5TMOrqYJwEdjtocbprQM9P
QsPlf2A7ry5ZYeDrjCPN6D5y9t2gccaGulCNE1z7Q8uY1aoCoJraqjBkE8TorVAoRXyHF28uFtnt
ThEIDRLMhWCpyMcbaohHgeOV++gUBiicnO3CQXnkGyWYdBgZRkmqJq/wLe5NPdCVbFGlxd32gWjL
NBchIv2KYkpF4CDoqKeHo9TmBsMnTBsbw4s9WJ6A/R4F76mM7m7vjnjricnQiUpwNcdu5ydxgtAd
2wJq0vr9T9xupzBh2zGh2Swh1UFfnVW+NMmjvQARpxGrw2Bt+9cj1rgDOn2ZvdMTZyzvQwpdPMHK
kCvF3QPybQaVKVkPg0iLALQrGBPXCTfQeMgz0whN+FhqqcGCPVdJTgBcPNfAmLRkiLx/aNWLi2x6
U3iPIZkd09lepM1LOP80i2fYtjGKCB4r83+D8hFOhN6YEjUFJcwMd4eTNBg3KjEppm+b8W/9foPG
FAbXRnp0iPEqqH4aHYa1lWGBpNpBWuFwfEYRYejV5p7qkB5r5xin6n5RrxX3wa5MMCBx4WHoShV/
5NVcYiuy8+tAq1SGFCkk9U1XsrcNTrw/adQSPRnA2s4YAIhoMUTcue043ZyVbeTmTK1bvxf6JAuJ
Af4xFW9AsbsojjCzDnkgAU2xCl2oTY/Is4F/umDqyuOeAAY7JLdqVLmxd4mgGOU5WX/mh6bQX8FB
gVEQorFICzFlkRftEqs7QmGdx1U0jJpuQ05Wh52Q/tJ+gWRirLa/BiZ4U4+m6A8KB6G0heUTG9uP
88N9KVlbdNO7Oi+9cxIZc9n1imrFHK+LgJPMoR04hvpv9rU2/FGRjfIHM7KBDOwixtXcQmy4nme0
hMNkcasqBxj63EHPpnezm7bVRU9U8kyr0emxurL+faKn52BtLF2YUmyoSz+9U20KRbo09w4Xt28H
mTgdsBpKe6KSOZ+1QfWOv/BK8ue0aP5oTLLw4A720ZgtzB0GGHEA3KbfubeffqkKqAz2M0IEZbFB
359tK4Rq5mGqBtPedigvCJJDGk2Gj/WW/XFBpppVMIUMe2rCYQCvNtaF5OzjeLDn3mP02RmUnFua
zU2ubpez8CMYt7xyM6IHD1gDJmOpf8pkV5uWpZ/GRx3KwcMpBVGfL6jAUOKpGtvFMHg+kxJmWBrK
u7w3ydkNvumaGL0mEm7Scg/xIoqswpXZX4p3nZjhAajzll/LxQ0dCSIL60sdBY3MT0hTnaUGTRE8
u2T5ULh/BuzL6qT9OCqD2sZ17RQlPc6K7D5rthks5OXq6fzzF7D0Vl55zpkOlrtlvRGLZQ2JobnA
1dpudzfj64dc7oWLudfrVdEPwKOclO9ESEX6B4If1QqkqrnVbHxHewh7ACoYX6FdRw83v6Am1hjd
PHP8VB20nlQcNF5hWCKHPNDY8j3WMgro4pm08KBMwPks29jUva9CNdU1t3Rp9k5kygBtxpAOxQ2v
QSUePfQPsWhN/jgSCetHvlV/Y7sQdgn1PDfmtgbXubbGpA9NvCPRwbAMqn6m3j7ePh8xLx16hJQv
TDKslHgkeOR/LCx34pdne9ykCgPLXnNfmrDsviSUA1axEOQ1X/8HMieN4kJQKbriuds5puB2PLQB
tiQo53Cf9PGPQZGdHS4HMobElKTmITkKml7xv8f1KCrOn0M6TDHVEp0ZQNeF8JzTMuDrT07ciJBg
eKfFON9wRbBbaBga80+SraiK93r3NRj0Ultt0hiw0U29HsSsW/VI7+DqyURw5O+8GhTpRT1p7PBf
CXrtqx0w1G7JllP9e4WMSCqYWmHwcVqCmclHfIUwrvASDZnF3OE5M2o3OsDAJ9CsmLqDB6ZnAYVb
sC8FOP51zXeNbzEhwcg3kPryQPvasQYoufoVO7FGFQjwd/BX6EHJTUrXdVdwvKd7ayiVzZ080pPm
qu0vwP6iaDQAghb937r1SFrZfYuLBn+uKWMeAGymg0fKThiPqk4z6aGsH20ITlwkkqqgrbc060Ux
xG9dX2ZEu7jaUyH9vzqmRg5oge6nTm51/+21uMzYZthFg3kUpWhVOCB88xIve5chnF+vgJQK2le7
N/LZrTUBYkndRD7imVL6Qb6/0fmFEKVupb2qtESjxoMXe3AGthJaLI93RErPKzk7FlY+K4Y9aslZ
Or9CX8E5wI/GsDG1KnFM2Vob6RxuOIW03A35Tj5Zh7+V1QBVZsxAFi+FE3IH2dnPJtofLk0B+rdV
zVcX3rivkTpEzbQRNkaGfJ0gosBzmaHukQjmMTn6aH1tO23UrKTH/3kY7VR9MUoSzQyd81bQfLPl
s1GKuL+1bIgU2S2NTRUwaw2QrZu/i17I6+ykixXWqlJ4G7H/I4ubbKe9Sp39GuA4F8kEv5XFZWgm
tMYYvxVUqwVepnkCl/XMQ6VzFnjuyusjrp+M5qCNC24/1fhscXwvD+69U02TelW80H7yLQUYuRvn
tmoUUzRh4Lzi4BtAE72pZGSA0PXgaqKvtZh/3RAvE7Wm++5ihJ7kinRS0XYDVVWll6hVpn5L06R8
N1EEvNZbRRZAVqvU5aXKW7kUnuilS8lNkebUoQqq4mJgC/BiOJAqNORCywYdw05/fR5W8EeZw1y6
hZp6vdaqlG5n6IcFj3AdTMcDGBKpIdJq7OLUEtpYoZwFOR9xNFbK/FCkekiXzTMG0xsNkdys94wA
S5d8IxfWVJPQJaaoLLYAIDqNDDIWo92Wk5MCPikr1THMQjCZ2Ep+9sQbW2mcdl+Kd2G0m7nMrJ+Q
I9himwcTXOfr0/1KvKBod7d5n9s24YHLQbe0snuKSzqajJKRkwm7C9JKiwzDr0HkKbHiydkkYoEH
SE43cGWBZXZrEcs8E3n34HSIx7exkZq7VTu1FfYQyv8rwYlmjOIPc7s8UGrL6f/UtYrgs3GPSPBn
imKghlLVe9SxhdRtr30x+RGdR48qVvjNDjhvDzkOJikYYoesj6bXeeCtEhgHwTdhKLtalYDxl966
8hBiHXuZZ83zMsA+qFgmHub151HSp8n23kBq1DiUmkvKV1sCDug9pXiEu3r6UxAGQGbG8Haioj1y
OE5CvqUIf7s6cU1WJ3rulJGWl0euVb5gSLXkCst5QskJ8GRiWgEBLpjclr/Wt2Ik8ei7dZOl763H
vQ23ySk1DgZL8tp48ebmorKtXdQW9hTrvLArhvOyXVaTNYbwWGHNO8gNJPAUdQQlSahQaTqC+GSF
+f0EeY6ofpYE8RrZV+mztzCISKhgoY2bXDPhxBo8UUkPkSrvYFAomfwfusxgk4t441vm5vLi1XuI
bxsVrYnFev+GSkCiowpPjOuC7UrcL/u3sYU9p+iutJKAQiUS1ezJDoPhhKa/fse3e4oSrt8OXvXQ
Lp96R9Q2JV/nb1IsJwLZPlnzWh4GL+UXHK2ZZ/F/bkCeEUoWsT2IN78YJ168TAqB+27ExvT08Ezi
N4MD0TSSzAyUN2GYDt5c5RX14vNHsvi64OKdFi+fm3LR/pgX/1sFfCJRKyOLZAO/tXGnzXe2tFXS
INtiVINpVupZdvE2RNjys2pYnUAezpPdwEYHNabuWj3U2+wZtYwJn8WKSq+3/78dkDQE/6UjrhCI
Md5/dNXLCrB7G6NVppocDNnRZz3k6MXSAzLZLy55tnVAQFo2xPtNF6mR2DGqIM/yHL8PhUbPlGfX
hrRUX7LUWPV2XZ8MNo3OWDBZTS5Yc0HEwT9vAC0UOiRE+3pxecgRPnsc2AvWbCstnsmXKv3xRLFZ
mHklK7bQHdg6NQdOUZZcR8NwZkBHpKAarkpY7wsy5M9EIZPBG6H7vU2rsTLyTczQNwhx4NnUoloc
ZHIcO0DSWEmL6VbGyst0ZhCgRchhauygbiWQQejM6W56hA1I9WMHkYdzv+UnH5SCuxMw3cXazBcC
gJ2IOPsLJf4az+YDo8QlDx6v206pDq5NtSOxqFdkVqkzjv3bZNAWG17jhUS9dsJ16Vv7QxhSBRl3
9lr+kLIVP0RQPalwcwsXqALl0IJTQq9AUFQFJE9bThwfXKesZ1DMXVEY8vRxPW4RBUuUzIRuH+TO
7s9etiW6foldmcMU/XfksXacY/9XeDsde2YsBTGLXFv7RQUUtDM0AOQB6CWnsGZY8i3fsE5JTfkZ
bIzs7izblJ8DtQUn+I5HcnL2Zarbsk9Vt9Mhyfl09usKGcNQ80PO1JJ4yw8avAxOyjlqP5wqzTc8
vX/6C4bF++6kppOG0zgnBnJBqwYuVN1PUd0DShgUEy8j6lKf+oj5027kqZZPyGRS+t5UU48yUiog
hx023lbobAQJ1sxMTsRAxwllKPY/UMB0MQ8mhMGfFIkn4MC0Il/NlM7HWg5MNVg9OiZyi+zTERNg
KSVDfdY1GFOtGRmyZ2y8+upP11Dh8oczm7H3wnYcT6cJBSkwwqJNXWgBcgTNcTznUrTsXTpkhIyj
+avaYBIcKRHlg+LwjVe8nklxqvKHxpbLI+/ip1VgIENoExxphqQI+/44fYD0G+v2CMPStUEVOOUH
A+vr3LO7eFM3WQylKGdzyY4N92zHoloLgSufyRF5ciLFGKa6qLJ+4lHfNU+ulwOvcPU8kzZkSNdT
kRj+qXE1MeLBkf+DWEpSjGxmE7BMrR+yprMhLGAIQCfUXkEEe0h5pG+6TtAmB3RHktboF8MMGcPM
391X00joyUGLYGgYUm6rATuSpU5HGDm9MVwsq775dXXcr8tonwVpLo9/mi3F8j/czPGO1EtgUUwV
MQaVSrRorCMz6yu5+WB53CP+a9GJbvE49XWhE+FViv4Q5CUfCPcWCkWFG8f3IVQ2siKHzOmfv42S
Oilod5Nnyr8BOcKfy8UKXCNjMP2YmDZ44jbTjSZ1+pkNQXRJVQ+R8KcQwVHvw2nOJmCQLRP2qpGb
MrAlrxpUHV0s2oG+53yyKqMRizDcO+Gz72ka/pSuY2zU1jbXHo35xKY/pGeB0w2y8dJUVlUBA4Tg
dpF2MREmC5/eMO0utNCH4r2VZuaLwz3/BUU/IrPCSMkxKntvVzrfZ+rayiY4UsGGAYyDEx0nTbwj
lv9LNubCad7kEHl79MfQ/+ZQvdtUE23+EaqJ8pJL6ahHRNIzbhd7P7hfy7y3iiuJ2JGvYY9A1ySr
nDQvRwxb/QTvtFoXevSq2J5hknYwaS+aH//qrpzdJd3JPFDSa0hRysl+6GVqpqYUwt3xxU3yLz+B
G7K+n6AdiZYTtoazzv2I7o4LY9VcoTbVqhJ9v9NQjJ95hGdgf0lpBMSHaI0EImbfXEejQmClrxMX
JIRYFD9Ptau/FM35Gei/IhyzSo0fReUyoaMpkSasLO5vAGE6vGSIU5C0l1jO7NBBqRrgrtKUfahe
jqiyya6hNb3RDj4JBs2D+B06eltQrT9xVa9K+VSerJsboZ1VXVkUixaWcnRCKlKt1VHTBc8kPb+r
zbbOyXmQUU4UJ0LbxWUrTNa3McFZfyv2B2YNJezpvbB/Yf1ODzXWAKDinChqwxYA/E5rHOTEDnfF
c5RCWCNZSjpamCLUcsqWvYdO4N5bqS5SNPlLyuEfU8kLpttGBhP5R20VgK288ymUOfVFyxS8cIOC
4nGboPmCKg7lxnk4Fqeroxrpd6VnTF/vFJQG9ZDbTk2G9zWULNS2/bBAnyXkQl5HrQlGPP5yye1U
9x1A3yCqykm15R443Iub+txb8FW2wWrxKAdHzc39XhTCWiaLWpMuXHyxVfackmStG4xGL4gsjTBD
ihL7KsupLDnu3FQqLM96V1ORnuiWBeH0BxELf5W1DL/ZRvn3axINhkp3XwplZ0KQN70OIRTRklIr
8osanZd0zUD07iZIwC6zPV5wA70virhSCxVuMpH5MF0zrh7Mrh4bcLczMm1De2J29wkCnPM3stkH
jc3b94TosL5kVN62a3aM1QrZVvCRFPpd9Q+MQ+gVCKfYYgUPIjOSUuMrWACoA/5+M2S9YJOIf5vq
JNOkCdq1Ac9UlHkX2JXl9US9YVMi8Qx3fbK590tGJIhmnX3REypuYKoaicGj3Fu2BQU8AZa9/EQK
HG5axeezyCTlG0YpXPPhtbHeBdT0LX1DrksxMnasNf36SzKVGvd7L4piRxr3DISF6oBXXHflmRXe
BmGLgm8X/L5x3w2x0UGkR7TzVW396OxoSpMOvARkQJM95xlLuojiWlQU951EVLRB500QQWQv/vKZ
k/TdZDYL7hXHgIoEt11J0nvHKJenjFBUNzONne2KMDpajxK78xH16K3jsq7S46dekIMULFcsluJo
A0sVfMWQzEGEr35Tb4RYdcFhhDHpSYo0ckyLWv3sL66MBGHxnOEjSAQqC2FYrwv3b45H34fvARGs
mZNHzJ9EzdprpEiwPr/pErBdKA6RaYYRvJyCjTUDv/+K/J1TWNL9BxUMVjbuO/oufwkUOxoN1Ry+
5OrJ0oUAdQ285CB6mznvYsvDTYPWUIS9U5+bCxZQhFeMfZ9LnWy51wOC0Fx0u8aKf2rjcbrSK7Vu
GjdiTY8atqo+UX5P1D4rKHBIbKmt6QxWlkatMk5ppiSlG3wR3X60DjoEDyAm+b0EfskRZuuqB2yL
qMM7Qi6ucC2j84D/ToovTgHLFGzFYOEpc81kKKcnj61wOqfmwXfoFwvvApBD0j6wmM5BrYfzXgfV
CBD0lmoObUzfgwwmKLL3p319l0D+SXWs2+wwtU/+EYghH9SkFadjoZ980OR4Ac4E77e08r2kKoED
sBvW97aSYCAKQXpDlNhw7vDqCN0VC0DJwhSgf7yh4lvDbvoW7YGExnF1DjQwDXNXEL455hW9Knzn
cpTW8Msy9+qnDxUNIJA29NjsoJAdLdJcvjDCgsWsEjXoMXOel9TH2cJC7w42KAgfg6lfM57pL/eb
VIuJycOvG+q5LVRpy+GYn/QFlIy9o+D0cos6tZf1jNBQg5t4m2q0O8i/Y24CHbwkp3Nk8jnYDa3I
+dI3v+o+vdSqkbgjz7yXSXziz6bn4c8+JfkUOjJnpzNlIrkwT33+hOuiqMngIukTQ4W7/XtllVMS
56mT8vwp5PJBexX92bSqGjRE53k2FCG8VZMW0n77DY4zb5lr4e6QGKvl6VDFOiA1E1wfUWrdtrPb
3mhq8WO0fxPy0oWKIZqkKj+xrPjRFp4NWGfpGnsHTxcSKaXZAIkhc2KWqATnBNg6fzmgeFxNlpRH
mH03HcsC/eelowmfeXfmahncSsJxgCExWbBf0KB+BWm6wF4r6pUC4EF0Hkf+TCG2vmVodlOjRsH7
9irHd92dPIz5l71aMA7e1m+JDE8PuKFJ8F9BsdCZcvMQIMQxR63JXtf8P00GaeiNUuhQ051YXEkc
lV1y72Rlxlc2ghxnVrkJK75+f7liCHnOuuW5x3JA7NQ78Qt6IF4dWqFQGTyzPUO4fjoSdgXKWxmZ
ZzwgZOnnnBP9ZnieSBj5zt6UOCnNdZQJCXWEShviW47ka2sT4c7n4yu/W8ZErj4ac3Ci1MLcdOUr
LtkHYhH0TpeH6xiyaYLQoYhkKJ73marXKdWTKpYiv+PaVuLwLbf6/pRNcB7IIwXIfrAvJOGVfEWY
V47lzujKZSiqJqcA7M+gcLUKDQTNxVhGw+o06t0szyUsG2ruyqI/0F4VCvtKJYZTnaDH5/rOn/m9
tgH12XtaIIxKlvAZk5oFkyLW1MN4Vj+wiSitlyFDz3sepfNg8IyjTLRYT9sxKTXEloSiWEbDP+lt
7BIkC1IF+GeXGYMleXFSIxxPmesylesJl1Ff2IMtEtGwf+fzr768Z8KmzYUf+BpnYagBLGGmnFSt
bWSbMWlDxcLGSFSaxLyJRPRsyinvoUVZlWW6o+yCaFghiU+moQDmd1d/L1W3Zusynqbsgyv62gSP
t3+rNeYkqlNq0XaBBY4v91RoU5iLAEWnilG9BChEU8Nd/9r7/U2r2ViZSnzS6Enz+JZL/kpzLzkm
ZiJ+nt4WKGxpFqMM3OmdqMc6K5wHPCJViP9+rKdQ+tpfW5Holnx5UuBrkG5KnE+kLdR4BAs1+Hfe
kEJsSkBg8ZoIWKvf3B1wMus7dYoV8ab2oelDhX8mLWsMSvLtLKwuMh9nX0+Ie7BO0ZX8/WuQq0tb
ieWMJgl24zazY/7pc85Hf2sbz9XlZOBp3Rb4EWXRfKur7J+MRD2q0jd9WPaeHZlbUn4bT3bSsE8I
lOf0iIJ22LqsLIGaz0eh2JP5cvqERTqe+woDbyLHh6W/X3J0hsVjcv0UXHvWpxK1b9hXyyHA8sdu
vUQ/jIsEh5ya++ca+5IoqRoTp7caGaNS4OjJ+/5ohJ6hnixddxB8EqrJeZqPFh9vztbA4vvljZXn
+4r420a7UGBNQaxBSA2UZjY9ck3S32Kmcp9aQAbtrgxrISns1FF05Cae9F3kV/wRtVkISVxcr+bc
rJnYrJay0+/9w1G76lMTQcpGbkdQE26vKFCGWtvSpgiz0Jl+gWngbGAuAAxeCbY+yO+Om1iQgCNX
2rDXx+NPzJNIkbAJKaGOZ5rrfE3DGEfNnb2N8anXqDekGZuLiyQqrLvUy772Bes0zjA673o93N9n
RBzXR8TnZWV+JlmGfsk7pSojEPvUzMJxU/Z+rC3IP7Wvev0kTOmX+Nckp0BY0V1riwo9jR75kMUm
KgBo7hisnxUTFbV4qd4Dzt+RKIngbRexkMLmU6lpJgvMNAvSmrWRv+d3DBN4i6kB11Wop9EW7x71
CJLKkRAnOYWQEkOpbu+EW5SeFRFVJjrCeoq9d2pnvgq5mJOc2G0Vwk0mLGzBo8uqOjfgcoQZgCWh
D+vL4GAHJPzTqWR8S83uoNybGU1hgyFVdpiLy/Xlsnz+ETkJa8M6brPGT5RJyohrvtny4gCX0OyW
Y43JjDpz4vAKIs/l+OqeJuXWfSM2xWq02akPs/NV/DMO9wdXZ3V0NmIEwI0djLzLISpZKPSqoakm
lBcrVxwRsZFmLB8ekwbZvvHlWzVqlDeuUmkzUt7i9lIqwy0trlHubD4S7uxNDr+/5d2EA4wKFdhB
71yIrtyJld84ZYveaaBBfZD2lYSQ/7Yk2Mow7fPJC125WjnivquTljzQsCRrOy5JeMyIgLczXWxQ
y/RHC1jS0ETQr9ehHlRwln2nX97xW/DJNry9XLyHn8kAD7KozlPrLSzIYQbZAaSqA0s4MO2X9KE9
4MdyVZrJ5KNc6BQzJA8vg8P3OtmaoBThyw60OXs3Iw1NEAtnsFRfG4BHQMpbynFgaCeecj5qsx6t
iMWrYj9X5lUqJi5YtMEQVFrtow5yeGE0+GBIeFuQHiyVl6TO0TjPzweo2q7A0F6degziLhZ7Qgw6
qrNR14sKN2CihODBtt4nFQnLQJoRc9j6m2RJLOo82xX3kZ7Vqkotsqp3grVo/gkbV8k8fZNK9cPs
tBajQFE6DqdLeirVB9AcdDHrFW2lXmO1Id++xaEwnIfWEanJz+zdUIBvRSWht+aHO4wpislcaqeJ
+pXyPQtvphurFm7DxpGmmx78tSijXpqeMby1Ta8vt1w/xekNf4Ww3AO56MML3XcKKrSwvajEktZ2
qoTM8N0vdZ5H0e+XJaYa1dvtZVZW3aAOS03A+M8Wsse9HS+5fyJZnIchzzbUVXI8+uZZlkaRYNd/
0VtjDqi6HDpOSqT9yYm5aLOZp8yg0Tg8Rl59roXlOTgU9ZHKmXyi7OSmxjK7O0PNKem1DoZkNiK4
FomODFiQK0pQwOXQxP7N7Y0lg8rAndZfEfI6fPu9t/2881bISchVhol+TihWjnYuKutcg92GaY3E
IsXwwgdJGJ0v4JHgIwRT7+E7cav7nrikJLp6pU9jWWnG9FpSYsGsRhphsD+ek9XVK4Ha2sBqYmUm
4iep/f/pLshAgrMHtML60LzBQc8ZOk7ysgSoLksspu5KlXVXf1wPWlcZNhlOEiRPw0ScdfkZtaXr
1p0gQFoG0YF+xjiyEi4pGKARdCQJAVkV6gg3X77xz8BF6z4o7juaRv+CcZ0eqyiceiNj9V3+fAoP
HgDcrEl1l8JnEvj3mymmU7m+t2oSVaDNj8Xz9vJzSddyFH5Et7+gXajCYlL506yLwbwaNHwAp/2O
q+NDiUsXMLs5AAwOc9+nVBRDSIS1UZHAmCNdipsFlIGMQSvM/wImB3DZSDf0yFCH078rBT6lxZM1
LC/gDWg5tjjtqDj75Xj1ay5HS8cFUE2My2XitB7CSlMI85dO5CD1oIxYh0FBX+/+hpK7pIWFSL25
rISkEX29X8Lm4mx01pUasBFhNJBB4OXRga4SpCPgUTojfH2p/ZklNkx4NZVyx5fbDqqRGeVdwtuJ
iHFpnfTKXmpvKLZMzQScrvGLWpLg8rlBBAb/Gk0sNBi6o60gIJyne2zw5dz2Koz+I5XunR0VJDUf
ocFpFZ53lA81idOR2xw9Hfk0snBKU0hJh2rak7d+bLnRoK0cmDmWlHBvmHjwrUeRcKRdF1bJeXBL
Rb5srR9ePnFaIlPe3il7NEga12hmcHFWubBBzzz5QFWz36LU41q72J0q9yXkvwdXUGlX103VLMDO
hVFWvrQsJIH+/0g3t40CtBwiv/oGmFEXEMmzo15NZEFgmvNo8R6irDUgj+0dFM4ySGFz0XLONAvh
kJQa4xeqbk93tAvgSHAbfCAYNvJfoil7vBxByyAegGipFUhUS2q7HbXty4uNsUZ87Tyd9L8HJC70
0qs3KsBuQP2l4MEZZbB2I629YV0zXRm/XP3hsyK3BJnA1KZGQBeBo2tAOS7nvH2NVIZdKjh7cqCh
ChqfBXbHZ5C581ZKh5Yxft55v7Amep9ETdRSS+3tJa4wqACLT+7fgGg7xPTsV42peN0RSF8WpJtP
TG0wX4R+q5c/hmw29RBtDU8PDdRhdB5dVO4GQHT+7iMj+Pa1iNgxdRiuVu52QIGgKjMrOUDqPXuo
Aea3jh/C7KsANrvCypn3ohEPm0m87SmP4lSpCHr+lzbfaK7mFzfzzdFBmmjPJRYiipgOdNEfyDFq
vcbQnx82UJ8f+yjNPbpAaZE8wpOSDqmo5yIihPkrl1bjezDU1AYMic2Zp27JdpqP5JtbEyZ4HFn7
nmWl0rQT9ewXMzOmyqQreQLMu+tFBdK6itmiP8/oWCRfBQTepvGU/dNypEd5oT8oqqWoF/l2p937
H46lW1+B0ARuh7Sg7+m3gyEAvEEmaZxAyl6jxq7TT0cX1RkBRIwDSugo7RL1XHyloXqzVwHtjJMe
KUI4zLf1LdhfzykcD4N0PKNDv1mg0pR2Uz6GD7wZNpD/D3K4eIFArH6YW4VCJBSDqbCzwI6oJGn0
9u0j0/oKpn0InuEwVbNGi/pITyVv6jYoJTjM6NsUrMjJZ3QH/oQ+eXkzwxLmAzmnk8MkjSPv7aEj
PmudVONDp7ZnRiWHTzJj2t8R6mGulMjBVlHa86Nc0hG8RGB7gFilVe8bs9R68ST9PJw0B7P+lohA
wAus2UenOTKVUoifM17utELCTa6VVuUmlMU34SqbgmlyRmIOF24VD6Y0zqoT1/ZGjwI324RsS4ge
tt878KQDwkyUUlC1aOYQh0i9bcS+KF+TMZISgAnCl12z5vtvzVGIdhnz+CsDANKpG4MIXVoH2Btc
wmfVH61Omk1Wiw5LPPcTUQDpg8WFZAPko92Mze6HR+TEpYUi//XGVsy2yJgbl1obCAPOmO7qXeJZ
ctzugpsYXwo4RSnp/IMLewv6FsCncBTxXVJ9tFxjACbcPQaP7ptrdGDzL7VQvWgXoEaMZfWi5fu0
VN5RL+AM3nHco/0BgeB0QTB1DEoiSB2CAv5LdvH3LRhe8eO/CtNAut6jcHYYhIHq9wNhJUJBd5v3
AIV1ebKmoKlerP4GpAlZFc+u9vEoHkj0h3JskAm5Mkv8mDwCzrS5lclZIotU+afmTaEeHfNs4nbB
flNIovMKoLe8Co5PT27HbFjlpmm7rZNxiCd2yumtV28yi0xjenYy0QVv1hE58auPgb/nd7WzOImk
U2cvSFeci4gQTk9k0BJS2EsSxUf7cclpBnskS89OZHzTPj2JwUu9St1CxNX/5qaioPn1HQflBJ0V
Ugh9fc+spdtb98oO0c1JZabTlLQPthhLDM/zAlyDT494qUH15EK163Q3EZ9hLEul9iwQp3xMHluK
/pH5TZdv6GkwkFur1zodyrC85sSCUGLKBaqoLJ7NOXoryr1g58Qa7b9KFRvuJOmP1OgQcPIfzCWu
jMxcMSlGm/Xd0ZjrN5YVHgQPQxFvQPvvrlykuNIe+RGwnKt4czSqBJYPgJ8XFMrD4QG+6HxLVlnr
mnClRzll9QX2ZIm751BACUQEHCzcnN5/fyb+cuZhop11IHcFWnEGCWCkTG7ZcWry9Db1RlpJyNR0
slHbu1cI/ki63xpnY7ZdT92/n90St5JVb9d92wV+eLrgu/vgw53mqy+xR9DLRYYwfg1f+naXBAEa
aYs3xIkyWUHSgXcgu/NGL3z4i/avW44KIxBWwQNdV6a5mRPW/qnA2dcqrRosgZKIEP1nRBJDT45a
dLqXTKMaNsbyQt6yjftEtWqqp6spb/pOHCgRbBw1VGaG53YzFp41h4IkCnZWAWlexFPtyqy++/V1
maQSd9HMd70Asow5hGVhkzrq2hNXPl0B9aJ9cwuA4HgynB1RU7dE/G3znHverivXkddTrhFtbqtg
kVgLnjZoS6rbHAncQ5eWfXNh6lKSKozc+mcZVUA3FDhG92VlNWLC3wsyle/4xlgv7IFSb160Ls57
JD0sE+weAUXd2YblS7qHMK79k8BTwWJ2qVedY20OdMNHWPV8h2V3AMJdwRcV+64HKKo2Fi3atuwy
p7uySG2ugB6wq2lXxtKbTwoN1nE9n0Voqi2xrLkPC3Hav9XCxr29DdZtcYb3MM0joJeTDncumcbk
NboZ/zQTmoJBlRbmomHg/kKswcMb3NckNCTZU7+UGjIIvzmUnbmbR9dcFOLwxXO0fxAmjYchDQ8I
GjMhg/1jg/TDkxdmGwU/NUVjC+6suMkKL21TyGjG/G2CDs5t6x6DAvM3xDDD0oQJKwiFfXN3Y/nb
EpZBHZrVCkoANv6sZGujwMjkazawF/Tc7J0r/+sVUFw8kMCinnxDsP/SlXnNSz/1nU/XTBf0T9Yz
7D+zO/yGTzwOozZtPcsHdXR7pYWDHINdXWlpMtS2a9t22H5EuTBzDqf4yGGHNdwRpemFC4NqFLnx
0zap/yaaXFPhZfACoUmtDcYuJCJXOlEIS3ULBTrIcBmBwjJ2FJHTfrOzU5OfwtwoMaL1bhxoo5FW
9ntxBn45W+t823WHmu4fM5qmNjyKettQeNILeSy+G9Iz7LNBoO8Xk4tL44UTgnlIyOgsPPm/M30w
WUE8TUvtrlEBDdKPt/H26Q46IGPicfjp3TmENz9l8+OLcCb3Y4WNYrbVtOAjWD2BuNXQinA7s87I
H1XrroVD830OXYOMTPEzVRDlk6jnMezscZ855HF6xPa9i2LVfiRH846/eBrDwibJxqipkppgyMOi
1WQLoPBXAymgQzQUSSH6eYVMhk7rP6hpY3n5vw0fF+Qze6uQs8KAlJrLUNnICCvGVD00roiuOe1N
ZnxLPzmfMKxfrRSIeOGh4nsiLIgz/DGqRgsVP17AxQKguu5yYbCfuiqJz3GmD6jsf0UlNvCIrn5b
pLcZh+ox7vFhx70dvm+/2a7/axUI/iN9yGwAHs0Iqrt6Zs6hcwJ+X2+Eq/S3hDsnjarIxVke7tNJ
oqUrRRHEJMUJM2vA5P2IZwtx4Nl/oI2FbWQCruOVmTo6XACKWuX1fwQ9j+n7iEysWmfQjgX8AIkP
7SQ1xd3VTbuUosUiWsM6rASGdJk3YTtsnSmr0pe4BWW2ag0sJk7yFG2t/SP1CoRJL/RgwuiQ5zsz
ea9gbm9Tq3fIAOBILCKtpnWxRCmoljwDuEse2MUfdbJogcW4nrztwUAKinNl3fTpzFvhD8ELBuKE
9eH14n6uO4EQYFDJS9ha8SFV4EkzbubqlY3HRF2XqzD97BLGH8v/kfiGAf/45PYLHZ3YMMW0z3ep
N9xM6C5bCvAYNy+wV3x0o2I/1xQkpnlOLrNhO8FOJ0UOlS7I/0apaTK4Z3C3pFluDRNlG6LVmd7p
pjH2kA8E1cuVFHBiDPEZPQ3FjPVVP1O+yXwmdph2sKEhxmy8jxrIYSUd4Dwf/zMW4I6DC2tpXV7D
B9SvV153QJ0bQsmpcdNwaA/IcN03fNVHwdM2VV6BlCjkueP7xukRQ1W/8RG588Sli1JxpLgnjQlm
Wq6TthpIQxwkAip6f+1WtXp2O6DqMu5rCSY5hpqfdOBxXGsBCYIceMi9kvlgPDrwdAySVnwvjAnL
ta3/lgShv3g58rv7y/WddLFQFLfqlCFlrDSbB2QG4dItBCv/C+DQzYD7lZ4Vpw8Bv2Q6cGqKWzva
dnY/pTAo14TfK3eDZplPzmqFosOjgSemJ+Ns4g8YKCbfOJL9AECxP32z4TZ+cLR9WAjvENm79Etx
pcbH3Dl5p/WU3k/f/XWkOy9I1UIAdJlkoq1eVQ7mZj4BUm70O0bue5BRQlaevAS8zYS1mo8Eg5Ru
AtIl1UxA7111Ck9XYKx13TW4FOPdojCETq3y65UeuPLYsOBGjhAOKNxcSnU943ZMlwizJnvRERIh
yTxQpEmN6XEWq04IJBCdsQy9AGTmn6g2JS7Zds4veD9YERfoNZefdCIKTLhX3fGOCLrn36pW5UT2
//bGPD5LIaVqveMbWdJ4y9w7h+QK2NCIvJCsiHgS4XGRb8wydO99dS0LGxK+BKbbR3qBKPxeQxuQ
LaathxzRHTM7oBqz+yTu2AHEQAsRiPFr7pOqL+KjeKdEfd67nGWuvgazRzaHD/4wXAdXlFPEgR6y
AXo8oNf83CG3xbtJ1uOE7fQ6bvX17xrJ6nnCsW5KJXYB6pBpxFqGp1FRNlssiMTe6b5K2fJ8f5Fu
2KpmhlP97gbaSPSpq4hy5k0OpSDhmUfYXoTlTUXwHnjzBoVx9j0W0LWt9TsuH5edIdUEDVNRHifx
nW0v1cvq34twGlIiEzDlccCpUbWYHRjNRBs7oZZ3nQHdmWgHK4DCC0fhNdfOtDjiAULzf7BChd8n
P4JQ6B/cAg0pFG/NoCTCRFLuPWPVNhP4zbSFJM1elHt+WIVWauuYsmviMTHDRleym632du+P1wF9
vL2n/JDG/RyAps/z7bxLnce1hiQFYTlieCQhkkKLJ2GANwhOPUxNO4FL0WqJu29MUz+z4Gt8EeTt
azvOdvbtlwCxNAG/FfhDsTvpl9hJpBuJCYHEkK+XG5xPNk4XGGzIHAvKJ5YVmJYMVZKDy0OuHWit
cVxOOfX9MlORN64bPikbEr+noYbtQSsOL3uxlCPPudgFsBkyMtLI5ykzPWVUtZhr+MCw6mSlNPvO
RCla1Cc9MVYtHh/4pUqHFqvqMjsGk19wL6GgwkaBSLhvsONLn3NoHougJMLVjmnExiha+Lzry9MJ
RZiLaM250YHTFW36MfPvmjO40PQ9KPoGikrJA/RjRBR53oLNxdACaghNOLxVoPkX29tMpvh3DLVh
aY3I+yw8UHq69EjQaIOKRxo8ed194RiKN31x7dwZPuJMqGuD9u2Yy2/jd4IV4nb/ODPtPtghY62s
3qNVtswDswcF0AKCNhprOYtc6VMIvsu6Kh1hsU5L4JniFnmHf3nHxotqDw617eS6eB63r0OuFaHh
A8VWhFHKYisiWOe3qVsIfQ4TObdAot9AZxjNsF5EY254mJiGLCxKadYzZNnmhXL2d26KwY8dG8jo
2DSqof7AdKP9mqpJnHjNRz2ZTxmwDHg5U/u9Q/ksnKw6I6S3bsh1rm/7SRjKpZL8baXnlwHnPckL
fXHzZc7qD8pMsGWtXoKMr5YVbuHHcqWNEkSQzsvu819MmuUWw0NDAn7UALfdLW2su7j6ucaL2VXH
OOvoroalMiLIpVcv4M3KfdvPe6Op7cU6f8ofK1U1ZuUtA7sKIWVhl86T3RaJBtujaf7PXwvuMvFF
DZMdFYPRqwZ19E1PmAxFKE6prsUz0PS8vrpcxTLi5YmMU88B8alZR0q+F2rRO9Euw5fsBgKq5470
fRRlp6OeTZ988uws6x0GcgnQeutPKsl99DZOymEHL3KXVfYVc4nfxikAb0mTpEXQQlAVwdqJIPnF
L8Xc04TvG1c8gdTMOGFl0//JgWXSCevAh/c36G6fVb0Daj07kzZtQIy+v7UZlVKG2La5l2mgpOqq
KYopdQML+nbxFdyf2GGHzttTnXuaavrb+Z4RUX7t8uzMWBDoDk2n6svK6uWvoOGbr8C+xij6HUlo
aL3GfhK2rvtTUHCb5/MCdcwgodpJLDpxQbOi95s8G4dqsLHrV8piAENv51AwnyY5UoEnfnKDL/M9
ibtap9vFUUtKJCm0XeA7vNajducLjlidGSyyC4znMIruIaP3txZQgYPo6tV10ZQuLa1LbK7XR92n
tfLCgQjIJkjkYNOnni8DlS8lKIcz78T7FaK5jlCBsDsEQI7OhMoIsv6Xomnw9XxnR90GdykSnL/6
8RDBexSZYOgKcdpgeK0HNxJCr4gsjXMjIEHu4l1th/Uf1QyDORiuLB+AUtoLVdmi0nCxhA9lgkQd
HYFDaLJTyV0mzzPx+wSOUTwNA/ROtp0cgWDVmhvInZtFA2BeniZ/9NO3VvUC5w5D0mNcizx1Xxkj
7EU7JWSG2QCuxaMsynegSVzP4QGdkqU9iUNKpcNTDj5QGUq94uXmrLq55STh7R5Vf9B95OLs07jv
0ai3OMIjLcMpnfMc8dvPkVovLHSjJ/tkeJdrPXG+kCzHx0VnUs1/hxcuhFJMHGMJA/Qbf0fOC/p4
/PW8J28XNr4bsFdFXTsFvp4+1PNXw+GtX8dVmPzGrMsAmlp0p+/hyroL9c5Xcf+UUqBMbsuuFLG5
l4OA5T5BeYAfk7uPZWJfz8GmPp0sVGNSDgUFi2/xKPQqgkI6vtmYhgN+ySlhRs3glXeFXcDA1Fr8
7myAGHkRg1VgF+VoA9qi4QNIepPXcWr6hwux5uwOs3QGQx3zvXxOU7lbRe9u7NTBHUkbmkwsqmBn
6Gy5P21VLKON2W2yIY8CiLZibOTDA9cgYqJEbVagKKzy7mdhSGuCBbomMEf2zBPGcpjYEKmGt8OP
VB2O0JsoSofHCwILRUvSVBXmWHfpCZk95rJaDlEIlA9ai99sj0EjQ4M8GAWDMwTG2Z1icZwuJe51
q7Eg3vEpkXQ4ijEOBoErbx7jD0nE6vcTO06cEJ79MqmxLSau7nU53xyAl7K/lEia6Mkvepgzu/Mg
+YlcAOMhIt5nfxoH5r3n5tmlSL7BtCyXZJonfbK5FI6PZIzyxhcn5I7F5yL5GkG2/sh93S+yMHxF
NDq4+fFnEcL4PShpO2UXVlM/3lmwHiTBdVahPSarMDEpxpgvV5hJsCnYWCE5w17fWOVodyI5Y13D
15Fo1UCBvpOoPB5Hggv+Ugkt/ufyl6I/gYOhn4Lj+yyLdCX939F34kqMBAO6yQS1V4PjwUO/Q6xN
KMnXSZGTKG+EZ5inVC90Aw/LlaV2vRpcP63jPqcYMnOrICyGj4xN8eRl4KeOIslMwiimd+FZG0Gw
dPm/6E8xH5fQ6tlbCENePeGa0vCCazfTINwLF6dhg2keujfDGPcN7FPGipddbHI7HabmMEHS6o/X
5iadMS8pQG/v+WWUVEyAbpKgI5B7OgJC9E2wH2W5IDkZzy2ZQN9+6luwd9jVQC0M92ALz1lmCJUJ
+tJWAe5Yfqyvr+IF2bLsNH6s1o3QHP4qVB2QKzl0evtxiaAYwGjrLXH4eEyFf9KqK6MzwvQ/zaOo
XA8erggdcdNuCOlqHLZrYLGTDfF90f7r7ABajjNNAJXCeTFNH1Bl2dO9GWTmONeBrPMqtDsIqIq1
nve4Jm3s+xfhQN5Q7hKadiV1mbpva7oLBU8gkvtD5/+rClJuOm6TPwr0IF5esBAcPK5YfK9zRfCe
Fz848owPua17PHH4QW+5PDh+CFREJLJ96lloBBgfM7Q1dFeY1zSnhj55q9MU2ooHovwc8id6jHrE
EHEhfdOIXfoCNZoMRXQyEbazpBVRfrzvqc8lZTOmLrWEB8Glt8oTKc2QWxPg3Qlb+nXvgM0Mi/To
bBc6/imENqhiQETuDDqH4gPsCieijB2Ps+Z0n+7gOFfZaIdY6mA+XgdrNYEBmDqFppslEKiG1s5F
6eT4Ne4BgusMYZVcCqu8nqqGmDi+MbSbcXquiHpCxuua21lNwWMB/EXYZfjv+bJ/LTsQ69akuOP8
xTBeTiyx7lFCIN42GgFA1dVXs4XGkDBHL3XNeGlB4EgSLJ1pHeybIkLXHwTCYCj6rvumcHHufhfl
LAY5Vpw7P5TcQb7wEGI6g3AxIaknInDG/FU6Tn9BEUa1lBoeHewERZIIzVDdTZRwZSDguwKtbJQt
eH933wpZUYdUhtCVkXufdO1iKsMru6t02WoEUsOta3gwca0VW2i9L0pHK+IxIq9kWWZV+hddX6yE
P0xpSHSXpiLyaSep10RW2KDXJvd6wEmwfbZM7LHDfvXnIRDg/I+hDnZT+CrJ30uUHs4RFfP6tmzB
tY/xJf8i3tYaD7Q91OlG5tH4QQ2/VOfgWzBgnU4Umt+xojsVKD1GUoMnjLqOsuUpsaWj9dkf5iv9
OoqPuhLJ4AurEXOa9ndW6sKZe4sMYlSxmzdKtxAOPXKJg/N6Z1jxoh8AeASOhyx0/I03iRhq+2qv
f3mQEFooWnznfasWC26JiuWBwdR72hqRxNsEe6b0/1hIkfuOdfKNJ/5gio7a/awSALflFEdtpCr0
2eY0JhtO93bYooG8z+IPh507pHtmVPR0XNAjnfVM8axOxOZ3Nd20CEVZx3VK/s8q+nJK0xlggxpT
TnldH16BFnWnWhMnt3pCem//5hqkpH4phLtCOUfY1PXIfKHladuSv+JNLGXtzN7P3gOirAxg4gbi
mno6x3ynqSc/MuCrvlVpBuuMM8AP7/Lvdaa79O7ay+RMI7shm0lhRGTFXk1Rrxr93a0A3XylCLgR
Lo4tZu8BcDeHtDnpfSKHI8bPhcTEbfP+M7XnOjGDB2M60j4NG0G03LY7ucCBLC3gxni5SH4cznk1
4vCLEIch4ajwWRlKhJZrIM7+hoh4rUDn5D/JP2oE03BuGxK4qWrOI8dUh8KSlo4Zj1ASeGOdkjq3
vj4IC+6tgYkJRAqNshZYFNnZdT711bJ7NJaL+HsedWWom0qiu+Wtem6WoB2qw6ign5NcrmylB/Xu
E5XHH/OkbmgS1NWyz21R3jynvr0pEa1b7qlzF3I1ah8oR666STj8wq/JPrIuTMOC6HewFUcTCnPN
3/TQb7d783A9ZjLa7JERgMj4qhfcqKooETcYMxahWMSI1v49GIQ3qjcylbfjtHtQHai409EsqjNH
UCUserHaoT413tEqMJ4TPFiJ/Flud87lXrjBat9KBWx55m/+XZGD3cH011rJX9wKkdAjJMSua1DL
AvsAzKvV7NkdKdAdiwkTNwwUFJlhraSjiISEgy/smHRLEXAePekL6ohh3wwAQUmJV66iJ2WXghxQ
l+m4HKZET8PmrZSnSf5M4OsjWrx1h95fBwCleMik3G+rtRCCmpw80p/mpn0yPMyX14oNsOS+Whfn
7h2r5PRKGFaqHo49RT+zGyhOlD5+jS+cc82rCjO3l+thGchucSYNo+1lqVeslFDAaVMFubTrij6Q
Dma+ehMgWOWbDMNiMo3YDShBenslsPt8IDt7BfkW9GPmfrtddzGPrizpAiT0/c8KiZapH62WwH5l
O2HjIS2RnP/wPbES3Qo83VoIY3n9j+MbMCwWyMaoMD2pr+gFsYra2fnH1d5cF/SAPEfRnasvG7Go
VRgqeww/yx8I0mi+gCL8D9FtRZ5MIV0QS/WqNZNZuqXSmfTJXZwpZlc2JtEBxFApvvWRE7mF1kns
tPX/UUZvdci60yEpnotnReIHqQ+fkFaxwUFZiIHrKKnT7xTR1cGF+MN1DmVQVDu9+l9j40O7Sjgp
w53Oj4yPsHQh63IdQ+SA0MbTyml0qOCJun2NV2KhfEVoUphjEiwohOVSu0HZpEy5AJgACn1XoXcu
4plOBoRQn1Ra8Anj8WqSFljNMQ1vZa5kCBQaGiUjvSWoaNJ0G6lTKfpaIo1sVD7RzBxZBEzNthS+
0r60gSfvaVXCaQjR+H0ktWB35Imd0iEw1ypxfBJCNn7+C8OEmTrUED8GdxyoeXl/rOgF+vJedPJk
3DOxMaWJXb3+QvGOgasK0lbtEd7RxT9iHGfI4RYl86CYpAhv7WPYCp6feJfCnylFryaH4z8Qttay
9wL/D0UvlRwCHJlJmHtiRv3UwdYw0kGcfJ19/l95B68pDWPQIlc4bTS0dLc0dYOlNpSnY0odDqeN
3PSDwLfAhG0PkXhmEQKfVn8rMGOoaP8mOrBxH7n17Ay2ddZz1tuSSvvkPUuORqg3gucxNGidRXjf
9AabSrvIypi/90REVDUVwZLIG111CQZ3zBSorRzrTpiYtV/90xD/g+5rf9pG1G/eDCvo6aL4XEc6
SAYuOBVwZp+k53X5zNB1meg3Ef0CNBHo4dQwyGhPgbjFeAk8SJACZEvyJQP8ysCvuGMzGUfLzmqP
xfKE/+GD7K5lHZb1ei1KwnmBjQ7aF6SlrMWqQ7QG/WZztg/nSlOBqqXRzJ6Qq5ADLAYczXiCkkOU
RjgbE3po7zdo/3WLPa+vFS4clgfFpgR+TEoG6MMr/7GSt04Gs7D+0ZLSc1G/k4gWyIlbZwo3qG6A
IuAnd3gJnnxcWq0nWa2D+nJYx+Fbl2Kb2B6VOwuWJQ0IezN3UZNwPVe5Hk107BqK6Td6OIKKtyTk
Uv2zalQf2/vLBD/YlTPZ/ecSfnxXw7ot2bKG+hKv0vH9GznbROzV99aBo20ICveMHUwMw/1MkDOy
KF2jl22nDTzOgcHVUglHNVxYS8yBiWVbi6uOkl2Ctu886Ao68zEqBh7FTqOD8nw/tJuOtNb4cqwb
RulS8iSxs2j7e/jWLhFveHfP7tuiSnoNW62mv74+eihobuT9ox5iz8wG9dDpAJALUvE1pcoZFJ/k
EjIkHwV+8dqy1mykSYbOc2c58Kam4Mm+ORAqrsELtws2Nl+zK4ai9m/aH7fuydX+0HpkSvkNjK0U
zi4pVPT77BJVjc2Qc4HQtD19QbUjgOrWePwnozJhQ324ey7eC4QhRW8MkM6p3fUuDf8UhXMIkGhE
ogYovt4WvlMIP2xaAz+Ii7xWBgPh6WRosOQJ7r518NZd53tKa6nQVV2Q/b7n96RVv4RLsXMNeaoS
MUVMKANlKlwMaIJhRQTl+yod3ktHAb3gLpu4Em59+JKm+VxrwSPwzivyF1FB3PEXqL5SzjTJOgTj
Q3D1tzBj8SVgSQylOxxNrH1m1e4e5ZkY/dBvBgfGB+tPQes7NbdU4lG/mZIczG8puMcRojCblvm7
pLgkBDbcl+kS6Ubxj1ZPKG0HY0JM7OBbUiUBMsNt1ESrz2QmnpDsoEyz3BAy25IUe2ts3KDPVV/F
lrgVLfJkoadrxpBsRRmoY9FBe1ZrNed3Ck1RWSCtC3fBXejq1yTBrFV7cAx8/McIAIi16yHm2B0g
oSjIOjOejJv9Cp9A6r5UN1mwz5mos1/txJ688QMkQGeig58YxTSgJi2JrKJMP8pLpEWz13rBpDZw
iIGi31Hsd/0be3J4HPAOEGiAPDigyQt7cUVYByAwlmBvVABzvKcMcug2l0US7BU7aMg+ZD7BVZGI
B0GbUjkg4FQhntPKe/rzMtpz1e15UEt4ZUa4wsdqIzszidgjV+qqeIrOPTDj1hpo25XSKsxc5o46
pO7mLjhSY0mI6IY6PFBgfCbFH+A6u5yjnhixuSnN/LHxDLwld+/GJ59z31jZjKu9GpU/lwRgGZR2
RIKEhzKTrbsVjLsBRclfqIMoe/8BuI7GFLy5s59SrtYJNtOcXnzxAjkRXvqDgTKXHU9HwC1NTVSS
K9XzYk0rYPqBS680G+ikc4OkCQL22cT4UPpFwszRGgW5BCT1bXAAtDefjviP2zFOw5kCYFQSzCuC
1YYueT8EnxCcLIv52RZG/4v2WK1/JveKrx2MUKbjd7k4Ilf1YMuTDyGyH1U6UTWd7iZV794ZXVlP
f/JXg59MaK4Lmj58GF2+BTMTXw29fNh6EMloQzHXJyAiz+GOfoL3f7IwymENWsALdnu2U7Mb80xF
2zh6sfKpU4yfN2+v3hv6tfXCdbulRw3pQF9a5oWhFQwOB6xd0h7ppwedym2m6q3ZCNEoOorLemIo
YN00lvfGG3/E4eWuMZeNohMfhdOLKpZmVrIrr8K82BZvTVgNYed19akFKUEoyVrudwqd4QHt4F5D
tlk5+3SMZN7SS+KlhqzlQMqj1cgfJ5GeDt+AlreeZpS0MC9aQ9gi/eYZUkuwmKJWMdPv8+iVaSmb
tv9ffC/YOD7Q33cdZpIopcWn5n74C3gkwvROmu7s/igNVH5YBfZtUcLNn1Gwo7tQswiL34/7wZhE
zfIUvISDDbtpVHYI7hjC/4KNVkm2ohFsTzULcZHv/gbL0CT0x9btkHK7+K+N1kwaI0Yg/29V+RAP
6vLfEQke+trWcPZJejeLkPskTGAdmglmP+tjgbVXcckscHh6WPvP4sC5/QFVyndITrJgej7k3YLq
wWhogaDzJQPdAeeTVqXti6aPHJnQUZGV7zR3LIpqp3pIIoZD+J1MjOMS5IUk/6xUNjUSlEZE23db
7ZMEI860/WxpCU2P6BOsHjJv2cMX1nlWLAE3GyI2XajKR+tNNNIQFVwvmi8vdlEWS9hcT6g5uQIA
o44ZHwGJCLIci5w8QeKWlzv7S6Qsh+wcuZgcWQ00VPegZW/W+hzaaO9zjZXumWfSjoxHt2P5CDtz
bdaKfNN9kRyvG9jIujyjvF3Hy0xKoBURZPR15HR08U+RP0uexrnVyiopErFKUAoXwjPKfj3WPlM4
3EvBDDdp47AMWqBX76WEH5gOTO1eKoFolQoDxpg+CH06bGrs0+Xyw00hF57yWdyFpSzWn0rEBcP8
1ormAx476Mb6V10+QcNW2a9IEFjCMsZP4jGqfG5GnxR/P9UfcCd5hg5zEcLj4HMpKnvSM0vG280J
KQ/ANvmWgwfL2Zh3BwTRKabakSv+cEg+oiySmR/SJuWth5zDeMR4HHLFQZGdj++e5LYRDJAfnKJT
A7Rpg11DSg6kLuKDyo/1mOFR/Up79+xgWBRxkxB3KsFZUbDC21x10kZxV9B/0b9H3t7Z3Pce0bQ2
Q5kdz2TaiWUF2qDeNiIneP9sbuJmA1j6CJ+tVSJI0AqRNEM/8snqqBXA04iMdkkJuireP7BFJzyQ
2INS6QRrgbPOTC8LqsHwm3ZIp1kvdrFWIuPO/Rsilt9Sz6yBIFPQ1l7qsqog6zMLLcJbJ2TFLiq+
7u0VwHsjJuzzokZb9mB8HyjadS9qqIbtsYdLWzPY4UGWCJyInl5k6Mb8Z/rMnkszhO9E98Kuu3oV
9jd66ZAu7KlCj9FkBRvYDPO6zGtGuGHviIQ8cYvnVRJIL1r6RALtHj6EFvuSkV8PnqTuckmaVMYp
q30paJ6UtrRd23zL1wi5yf73eSsmA0ULUDzt6DcpA4NZ/S/nd4VxFye4puevsyTVlD4+zVXqJ6BP
UuKFX5tRsDsg0McaE+F/qbS+jr6CvJ+9k/1VeCKjo66GTDKK8yuowMRxz+Bz5UVb/i0n+pFFh7Ph
IcjMNhMQJ7pnhydU0eil5sD1fke6S1wuenqohDcn6nCGhW6owitWWH9RRamULSUZNOAeKQXZ/8IN
8bXFRf4cT6GssFm4vJ2jHva4G0RVeIHvZBsNCJzvwB7S9fQlHoNfZtR9KHB+CjYdyw50CD50xVZD
rhQRtEHoOz7LkP+Ta4/WARmY1Dpjc2rqLQnrnV/MxM8U2aByLXFM8WlGijT3wloi8S1Zh9GajMkH
aL+eWp40mcDYxRDTM49zijMM0Ivr/zab4+kyRpLURVBNjsih8V4oZMvcnTTKDe8LYLGvEO3kOsCL
l1SGt9c3uZFiMFuXRbRp5AoR71Z8pDLFOtD330sqV+T1BeEEdXKD9dn0LVj3a32NCqQ1JNo20DiG
vEMzeMb/4Y+0vXfLCVjkQRsqwXafuTSiqeau1F9TuiuOm9x57ri/tCRCiNORMS26gxHBXrCjqnkw
m9fSA0xsJYSkoZD//mS+IBj/eB/rkrEa4fr39C18Dv8qT8Taic+/hXbRxamXeYZuVHmRtardFOG9
fsRhCU5t3MyCA4Cb/+AMtDTlxQ3v2ZyPkKI6uwEyjD13PiKZhI/0FtlC/6gfTyOwW2tDzyldPO9P
VptkHLmPmDNWuEHHLu8plbY03DRfGo6uDFytHHBwvACnNxg9xiEKhRhSiibxB4MGvPORq2kpvSDu
SOTwBUA7TttcSM8Ck75GegIE8TlfqrLJGjV363hNW0TP6JNbkH3/dAQ8s7Gm8kw3uuKucSVC5Kjt
Jl8HERTFzoCIMYWLV56f4ngj4cM2AKevMGKLIGKnZeBU7ZbiTDwdOap7qJMwbtf28gfd5L4lSPqG
LyhMdofsqfyVDzNkelNH/3TJ5odyL/nyPE/9GP4ovTQ6merLYEql/qaxm9Wfjrpqsb0mbt3N/UZN
ifUA65BYa+WH0CBPHqdICmB9faVJKNni1eP5rWNQznWTmXIQMTx3W58csg+op4etCIit+dSBe2h3
gqPEh5os/9tEHIo4HsbH2DB2YXdFQ5Kb2Btg7Jc3A7rQLuau1PYwLYMuKWOtiqWiXFA6c++eMwk8
8StT4B21Dr/oAqcdaCsIyPUJKUmK3ug0yC+U2G1H0MI3am133SISz+q/fxBTGsxf/k/3jhCUN05i
FNXAue1YRGnSZD6jE1Kdyojw4aIhGrO1EuNoJqgsGIkGznYI2U0YZ9DkwFFGYtDlGp9tM7NaI00X
15IUbXNGpdBEx7oyVA2WP0Wd8zD+0ty2/XZHTDYprKuzzEPZ+mnip5eF90FZQLR425u5KJfipVG8
Ie2p6vttJO0YrHwnFhyODOgH78qxeDxwMnlP5y7cYTqPHRknxKXqCp3C1eyZx2zXk4DEW65CREln
pZKbEFNv1goV3vvJ//8pMgtsAGQMvOTxb8gx+Bv8Alaellw0M/xlyOH3t0VCIVmKRuyggt3wYG/3
tPW2rzSwYOoKwzCJQ1oyRC1rYuuiRdCWY7kco80HFnuBxlZm8tlPWkImNN4Pa8dJVU+93ZYWUL6o
FKwlQ5snd05212BqOiuPf1fMKdOH2R3VA2e+G9EMRwpH063PK9V++TYvRgSI2zgi1kHNgdCMnp2L
Nkp/sIbG3s5TTAFRmQU/Xv55P3yZWL5lhVPYPmAvzLCUoWU2Lajw7VwAUXTUK0qNwD29mofL8aSh
seiUW5kpzCKPuFCZtU2q9qOeRluRWQK0b1IoiaaZ4amEb8U/bkgIfRux0xkWJraiQC/jO2wS2s9K
NGq3DxHkpfpJ+cMo2r5jYlJlNckm2YnUIOoh4ItM6MpUIJHl0NkQMsHGDuR5Ycqi9POnLnlL4g5O
jp8d3uPolR65c9SDEzA9yZJso4vKIDlg33NIJ1GZyPiRInJD4FZSyNAU57xQ+Ho7oHsWZdGNjUAp
7woKvhvLKUTxdiOtkdy0y5YSWmB5ettLvifASrhRpSz7hOg73cLKCCBKzm8N9wXm9P1XoN4EXSee
Pc/684ZAl/j/8GJ8DAS+K/3fPO8tx3MBMNH/sgEPu07OargsaxZ/RBcgYSpOb5zzzDuD0C7WHDpU
SJzDufJ6whwxWSteKP65KZ/M/P7bFmsEBrMfcBMdHPSn2ReI+iGBhigeiPoFbfxEu9JQEfrxVYVJ
UUIjfQBppTkkQ93o3Y3iSQ7dFS3Z9uPEn0ei+G0JXvq3gzUEkkkvv+zFs9bxt7eIwno09gV6EpX9
8P6gP6LTLEaGo5jEc87IBq1YqsFIZjqtKYyf5DINJSYKM5PxWIckFjYPL0hMOZMtiaUyH8p2Y/1X
7vOW1aRroZ435+GSrAh8sy1cDy6r2ruTsQ7mDf/cReJqGIGDlnS/y17krFvcUrReycR8Xzp6Mupw
jd63zMPeBJtSNTUq53HVShk0ezjQjfziESgw0dAavv5JtIpRqXy2Yh4bzO9wFXO19qpSBVkTzAzo
3XqMnNUf8WlCQHd7HJgXN8lH0jpQszRQp0MjYJkHA2wrbzfkMzMMhBhTAwlzj8csYXDsm5qIvhr0
AkVcARPwYd1kH9/kYbQOM0ooU4TiHoujB5tyYLm2HlNBVhFe9bs5BSFAeOaot11/KT7v/etIFpiq
7o1ttkZPfgnu70rHmRQDgoa3nwWISagkzMjpgAPgqp4Mtcebr5Ym2Vy8DzEGqZnruV9FmKdH23Kh
UwFMrAFsZFX16W1nPByWc71YQwELfnMjbXLDECzAXS/swsAUEg9mlKQi1wog4XVQU9MfRfzjJFSZ
k2re+VL4OjEpauYp1bxFOdPJEGu7ljg77qWzf44hZHdWFmLcQeKQKx/PahgzvRE4YKGlvGLxvMfd
jBk8oby/HqeqAZo6rWT7O4QhmEMglWRSy8OCCivSTnWlixyFvHCmZWMnEmjGpDmNh5+WPIwUMUA2
+mhCKP+x18svtrSPPGhQ35NtNKXLDP25+lvld4i1MH2D3ShVR6W9klbkfaT038yE2fPeHB88UKeH
7CRZcW0Ex+tgaaRM27YrT1xho9YTZj4zhcrZHo56HGYqesLwVLsy16/jTQuH6SlyM69UdOQhR0BD
KDFXEh11sYK2VRkA7rXuiDmT6l3YV1OlbCr8pKX/rPb8lbhLP0Gl/fYb5a9jNyd2z6ekpxWXt/5C
zpW+iqriy4dv91baxBl48N4Dx0yDu1b12TBuP8iwfbz+I5bXOjnCgzLNPApUCuiKdysLHpX5Fw8E
GK7LHX1RIAp2DzOl8EFuRFZrgAyIxq+c0zBLsbB1mwLf0cSU+54/7udJVOvqrWjwA5ZMpB7XQP58
xlDc0cI7yy0g02X2H9XRNyVB4JgTyOP5USeiGu6ClbhFM0iZTSp3pZowzwMm7Ivcwi73DtcRxOIy
3JAjH8A56+nBg0TmGOsqdc03wUDaAnbwTuVsWP0bVyXYL+bd+ENLrZS8tEujl3k+aukgFPBQy5ub
jphut4foRDOh+9eEQpP0m9n7pkiCToCPsVsdKvThQU3qKjAOwFHWT/jibTIB13liy/HjlgBrajMz
T670XahsvsH7o5YdcoAekHkOaVRIpidWZQ6sNXBZLGYJXJNg+h/tsHM5Unnt7ON+aUV1ZTmww3b5
v8O3fi91fziWYcNjx1cytK6aNkz2DxYFJbdZajBA/nmST0XeBMeS/tDPhzdi8cbAL6QNLyyTom37
D+6qvReiOrK3FoVBs3XhIn/ihaEqXMQUwgVhUxNiwXh5FcydNiQEiWFSdyHrVd2cTcQ0NEddyl8R
2wp4i+d2SwQSomhQEulMkP9AKT2Yi1VV5qX6UduNSIXHqM2E7WyxW9ChYPyhBEMZSIdrBj3b9Sv8
Q4FAnijLWA747wl5wVU3jhFAkY9hbyYcmsCGwUn0y4oQQ9UXiGiZo1QF1antS5T/EXsJgOfun7jU
6hlvkak8bEHxf/ZPt8e+yUNFP8aBEr3frMiSD+WZzoViz9sq75A4iWRP2hpIPc6zCjzDWrQCBZ7j
Kp+hFUU1zsgoXtu6KW/MgsTO6U9vfocRbAcV3pTZcgJOVw4a8J8LRuQqp4q8CD0S1r1GThBew0BQ
Djh7VQIOkZh213frXsXLKD3SPLay6mYlgD4rSpf8nEhiLLBBB3wzk/Nidv6EjA9GWiS4HzxY3b5l
MMrZd7j+Et7qTi38s/L2AjCjqG0HdVMtzC6yeScVNNgSoPSURvkH561yW3zVYmqdiJV3pQm2qRKM
EHgdcchpdH2jAsju+uTCxsosJG+dCOyLO783EByaDvbvZioWwJp24r8eB5P6Vgh3ZE1alpxqF4AS
mA3Baj4kFz9tfBMD3KJ9mHfPZndtrBXLBhiUPaHvyoxurSTJC2/oP2dDaZaMxJ2jYmBfNtUyXSf+
avtGbN8G0Kn3ML8nknMEPLyJJNvgutDow5lK2yOy9eYOx4kU17nbU5GUq3QTLVdtmMsuEMkQfmN1
jBp2G6CLNLI1gNyPYNGLeH3LelaclfB1jbMeUr26IatmXVFWfrqk7Y9dsBe/yp7z16yC0Eo+9Ozv
QEEN3zH7mFpOYSef//HHGBMylK2utlYzqpTu0XXYpP5VVnzSyeviUTRXheNaxE/rTMUg/xM2Izy9
Yb4Y+37X4WQ9RKxnp0dPs9zCih7mxxHal5y5G3ksdtNaq+O/DZ9gx88SyMhOdPFS6rF8VV7IXM5C
laYbzrq3Kk+6SnZoiZZPf+V+qlzeyisoFUmeZfvWQEMKChnX5Uc+vIdkWoZkmo7qVoNT3W+28rG5
1Yjj3PMafODI5y6mv5xbEserwMDPHzoEjnLLnsQIsLGtRr0V8vAiNzV1L/02yL88pxdU/qyfWZxf
3WAdaTD+tYjobO080Nd8c0cvvLmxafqwda39RvHayGCoEZUi3pIegaYNF89UDDwKoc2UIZwLhMZj
vOLcFFCUHOnDWl3TIBzc6BHdSAfqoK5JEpmT2ZhAlVVeHj1vlwXwl3PMqegKeIEKGTsUIfkyNseX
SaECHX0VP1S3HN9CzOx2DLTTfj0m4jLhd6VPiG3OEqtAn1Rz6XHX+MgrPrgf5Ao4LaMcHzQDlWyU
vNf/3a6MNAeSkp2ZslBUh/4Vd4SA4cqN6V4/Mn4tb/Mc9roFQJnGjPYtL4qxYfZZKS/HWonh1egy
XgTyF4uYnGoXgougVc3DiTfW/ULToqeQHIKqfr4uBSyuHZIpNbPOH+ngzOgJo54S/do+3e4jbqjn
ifu1YRg+WrH8vlFqTDKVJ3tgcLRXcn7xBdHasxFULy4IJDqtn9VrUBAPb+bfxp644HxYnQpRQ3B2
kftCV+MbLzBEyv6ZaEUNGMbcV5Q25jIUeQUkfSKwzC2wLjuOGKozPn5M4s1eH5ZRGbJ7boFZ6lwb
qWAQyJcR7y2bwJDRjCAEFjCRCciAjD7TsGy9fSFkVEAP9QiV59ylhMUUHMR28+CqaZfN1vAVPmSL
hSWtVc8M4T6teMaYMb+hwdm5l0lyLinjAMHNB1YHECMvS9BRH1Qbo9JOnTYNZpsNj8/ndZruUuSF
Hfb+l47cyruBqwBcBrWyYsncBwKAWOdip+8uBhuWH5a00B3BTyoG3uHlm6QFdIHs0DEzh4FJntS2
m5YBkgw4qpYLYKdOWkzAwir8NYxa1TYNz+gHMGfktbcNT/CEfrSrEbqvfbIRscu+bb6I/ZSEOnX/
2f5CVLMMxd4doqOagn1KGDq/cbNcdlNRI29RQ2wvUVzyrQL6q+ztCPvgS5ctrpsjnJO2pdp+XBIH
rK0VK79N1Eo/Xb+exT2Zn2E8s62aZMQmHMkhpvCIuBAGVq8qdgFLI63PYf4qRGlP+l31TvoPD/US
1MkRnHk0JgZjEF2N3qENGxQ/mLri5c1eO5tQyrx6iaP1pqC4YUBj7vXeOtXY9VZxzChN7msukt5/
x+rnTGLqbiGS/tb9YqZCruLuxsTohxuubykxwv9WYLok0q6t4FHGBYOSEFd+9kJAN/OibQl5IbLW
4lmSwkb3EPMRd6hIg2E9KIQJSjLChlCs6W7Apn9jsoOFbWU54Sqw57f9+uZnio06VqryNA/DQfwW
X8TldYPmszwzF5lbF4MgZFqc/xAymxyCCFvPTHVTDgS0U5qW5Oobjo+aGAp2p/Rcbm5T8+cLrbv/
1NfUv5MfyP46urE8U5n3d8HPcHdknKpuTAWzeaN8coDMx+acyas3mrofrPh5h58z/+/LsaNGY4Q/
rsUVfXA86gRpaCThBn4bqawl2TK3pweP9W1VzsL+GKiM9J84r/BW++ZzvcocdBHGh1pAyiJSnOFe
G1CIs4rB/tK4cpeSMiwHilTRA1ZKERR10tuxJ91I3Zym5mfHTTkEQaUisiXzl0VF3C/Pmy9+0gBS
/PWIRa8rxJbgHVlNTQf+ZXNkFWKAjy1jtzDcNbRCwVgkb/+FsPOR5AMYshgZKHm5GYIQOGsboTrR
ZNyWNw0WjSSMYPnss7az5R8XyExcErgvezaSmBDEgh9/CbEjeVg57U0JyJj5kDrdJ94FyCW3uIw3
21qR4Hv1i9Ox3kX5M6TAGWlqCf5B28kpoRFjXWdfA+5cDVdb4LknCMVOPdj/A+2crDyWieCT6Gyf
ysb5whJexOLKz4lktd+XhyGl2QQnvSx3jFG/LhcVLzfWfDcMcIC4s6rfhVelHSOmRZ6kGXR728Ua
PEXpsZlK+Fdka+NYnv3uDMtHv2NfUrWXw/AiJrS3gfoxB2LXAzsrFDoxJDvpa4GUa3Cj+9MkdJDu
c+K/jnrfGD9RUQJaA/fiCvygYHLz6Wa+v17HzmsAUACUoTdcHOuXxd1rSIHXNm5+t4PSVH7TA1mM
PUCk8Q3X3gmwlZCpAOFnlAvct6uIzRLMPkBWDVqX0VPMSC/J7utSS15M9ReSM4rfS5+CdIdTJN8V
z+JoIdIKEQ8WmDJyYxVkMZv+0cuz1RGrjVRQQ6+Fl5dZ/BtAOzzD2NQLqYVZKb4sUjHFyHz8RC0a
Fvet8CbqIgasWlecy+c/aLCkHORFpDnhzeDgxHp+WNHfxoI00nH5lAet0l1/X6iLgdcPkMmZnTnA
NfSvDWzWLDzoZcf13F/qriQZV0/m8INADHvjXchczWhJp2NLxthOjvRZRaCCoVTYLp2s2M+A4Gwg
a5YM2SFpToJtlo0UyKsgXXIV2NzP7bUL3bKSMf82QbKC8OmCQ5+nUyoviaoCS/oPczAXzape2nuT
6nDmXrhRm+YI+fWuXZ5Uve7hIbjvjdYPnM5REVhkGUzNU3YbLwT7X6FnMF2UnvIQ6GAh/8XMbXTu
oonX2PE5fGBCwmfCYAvGcFUVG3KVloj6QpeIuaNDiWMAtODhpXcV8az6zTS/O51PKotG+3RJwAcm
bfPdATZWXv2/JdkBiYlgfinHa1p2eiVw6dziRCGm1kb/7aNuHuajXhDUcQLk1ZohIyxROF9nR4lU
VyUpnE8JIC1XzAfHSGlrRX3iMqe6jFOzjU+st+Ssi2787BNLXSVSiRoGeXYWPpsgXp6zA4rTEvDW
Yes+fOF5slxCEWIf+4ScD4OmJHGgaT/5k/8aAwjhYvLGyHE+imfNCFvhdj/5x2ArLowq5/t0suuT
A225NPRrgUyx3AjHpv9fiqRa5o2TAfMc1p4pOvMyuA3RVd4P7fAjKH29/E8U8I/d0V/dQPAbpnCg
tH/r+NHRiCZ0CzODOZ0JZrhCjzam0VV15gJIZQFZgnVIkbOoQ3lhaflr/EOuEokyk/Vh1TnI0oAM
+CK0N6Bx9AVGN3K3olHPL7Ll7OkNCJtybPihG4bu7s1o21r1Dr+XxtyeAxZbEZbvpY8OG84hKZAw
Z7p9sepB5ajt2PwZlgLw0gLhmh8EkuaDerHFmxrynMGZVX7/VxByE/+C/Sq6WIoO87SN7CXBOnDF
u+d/WmuPDYWMAZcRXSOdtdrtrMHTWKlQmo00tqXn2H3/IjRYq3Ob6UygFOd+s0F7x02UvdsI+kBL
Pk/y6R5sOvK61Y7NrSIcQqDHHzv3nwqqwuO9RxnSdVafu1/7FcCwufzHnRebECLOXKsqJgPSVIns
xFTnLX0TfWIUehXaO6BHeQC0RMBcMhmz4ivL+NjHdU/wwtrblNIKGuufmKmkH930+OsUpsWbiRaO
9Zo2JnB03HOQB0iZQBJfkC0gIcDlaGfilF5PSbJLCTDh7WtZVqq34MZiZL0owqeWmnJXN1dbGVDq
xV4z8bO0yxET8VcnNUi2cLVUI3gl68bUaIGcENYAsYEdpIDRt/QzSEeMV4Dhnxk6dWUP2PrnzWDW
qREiRGYJdDVVaIwJ/GMnTOgaDw2QbmOhhq0LiW7yXLowk8jk52HZ9ti6nroq5UYGNN+9DbM1V16U
2CWP1kAVYlJUITr9mSxQERJyNRgZAOpqavDIW5iv+RwvoAVKNA2Z0t2eU9iEFugZumLr5LVBqrJk
uSrlvnE0EOwQcPjJi/afdHGWjyL5WwdKXxdwcoSzbbjid3iuAcMRCLHWxTuGcLyc4RPztZaiz1eq
EiVWcMWnXwb30MnX5+01lYet1VNZ9DfSxMcG7hiKyAwDCAmTAWtzlpgcb16SLfMN42vrZ1u9Lk4O
aoKx7BqqcYfmfhc9Qn1cj9TyuikETOggAl+UO84I+Wrhn+KhJUa70vjyM8IPDSi4+mPn6Ehiv5rW
vRwUuchfCzunNCf/UKsAV7FyjyQyt3ixQP4a+5JUeFut1N8ojvhmMi1OCpZvm3PWqyrekDyVddwo
JMuLpUppdzrenWd1U7+GIxDMh1p2IFibEE+5JAtnYtSYmb9R5awdC8fby3gqRafwlDlHkxXMG0C6
pVbzbyqdN12uuxWcsQSyk6KgbEwSiTSdDroFLiRmo0/Ia9I9SP0lQWH3MUaqRKJp8WihKCBWZDhH
pV0hRayeSWYMD/jQBNTALs1sx/at8zTQXIUjrzeLAQg5y3IIgz3ls8KReO3dAhUkOrMAYy9eDOJq
MJaC1e+jBc/M+U4piWd6vx0md0oJ8sJDMOqeoX41rtR8JuHQiznNDiJPMeVoigtHzCoaz6p5ELmW
z6+5SYP73XelxMqmWjjtwya7LVgD+eBH+BTKpnGy351XaiJFQ1rPq0AzbsAwTXgBhv8jHUUfOlag
4VdsjIBcj1Dc23NXcXQIyYYgeHuBxHAM2jLE2HUemCfqLPYdhP/OgM0QfD3aBKwRlMGFQph+5Aay
yHKDPQbvCXValdE7upvhpaQGG6pCoXUQm25ivJPzebqfw9luYuZEj0FdL1gSdINw6UnmAq5eno74
wjZ/gNNc05VRZRMxI2xZPQ9K0yFTwx0DyhPJusCLa6EgX1BCgx3CeeWu3MH3t2Vl3L8mElD0gRPA
6duFI++kukkg+Arnye9hvWbRt/tcXP24UcZMgnEIeUUyzIf1lMgy3ALEYKy9XL8UzesS5wGC6nUL
ea4H7ICFvF+Gav3iwQIjkxL/dd3TPVogbdwwavBK/idM31jYP79juVuFTSjdV6YmSND1gS/STQTo
5H6ERV4MX7xObseWY5XG6jUrRplhq1JbFeetqslhOYQyZ7z9UzzuoaAJyjDLJV4MCQra4SMDQieF
B0U2DzPiWXdlBwuAtRBXy4OYHCruzZtL5gM1+NfunkUo7qMXwxVySM0q2mAczbsWbwdVAkQ6bfLI
x3HOy6bku5XsziMdI8eltvqsAWQhrk++gxlJKLc5+8AG1d/pV10Pu+vaAGIZmhjnf1Ap4GTQQPWr
H8sMyyFPbkNhRRiR4BjUg+c8ccHR8O9E1v+Az16MLff9toLvke45zAd2eq4ptzQd77NW+FpAYdKt
QLy5jIJ22iw8r1+a4xv4v8NU81LRmIjUMAHr9UUMI7EqMemrQuro6+m3MfOk1b2GQ94zQWU1sx5Y
rTyRYNre4edJD4D8OYU8+CPz7yTuZwdv3u0BJrrDbbUS/9I7Q7SWT8vAKitGeQWlGw8YmATS6nI1
J5SMTRJfvIoPVnvwY3CZ67yOP6TVFxFgCX1yfQ5ovbvVsisRPsMtnC7r19oKVrvU1r3VVds4OKyT
xlyqH5bXSmDi0kiR6oYTvYyBekRmroZqMhwUgY7vNTG9gTMCLkV5fcaaLXFCtsOcI1PtSckMbkfU
8hxSdPYPsXSRt5O2d6A1QpqTrs1y45G636XkWhcsDg5mhuOFGv+ttsFKPzdYung8gApe84EUZh9w
69AM7X8zRfcGNcfzbipSS7jBVqpk4lgDKUlVol7MfQuAJumxdlXO2JJ8nv9r87LJltlOhu+FKJTp
BBkTo1Ddg/NT65TEPdYAndsrXmYtNBUS6tE8KjO4hZg02y7ihe+G+YLbiFsydjpasJxUQHiBgktW
tR1c2Ga9RqIQZQwVjD6iZmi2MhV6/3zRQ25B9Ho2b5Ikor7pP72uAk6Z4RsbLkTFB2S8TT5spd9S
gFYStKLgx2oD/d36Z0qeOcKaAXr8SaSr/IlAuInFqUSpovlgQwku+4Qn0qXL/1nzhJxB7KKmJS/S
ROjB24DIHsTuruzQaGr047LwHImkJZIBOFTeniVbv1bzgAnfnwQUTzfmBlNeYV8ow2WaodOCZFuV
wd8lIoI4v2znIfN5ye8WzaCLzXn5L/iIrB7kuEfc5Hvfcc2FEvx+1T+1o1C+zkwiWr7cMqpA5Uh/
DlhY9iEgQ7aX3mGpHcfZA1OsZ++O2ilYX07c/WcOfbZb3V4RwXclBej29h7YjgziCYxiYr7Xvav1
jLw3Fwab8Fceo7y9VMBxLoc9PRWTlNfvxs3JAcbnYHZd87iGTqlOiqfpDFdnXT2L0ZGXxsMK5tpe
dLV/ZSm/4m9Qe9BbtFvci31z6PZTYOUEhAmNckYkHYFYEYXJKLHXEwXe2Pe6DHbdW/XEC+cdYvIW
FZUib3EislI7J29gExUEW6IlydhdB66rCaM7lg3q/cxmGvxYd8ukGvE7W//BuCk9i6vGiLS3Ssn8
4l3/dV/J1GbhkCcOoCTV3WCqgYmXBCPMdcB1xaNsWJUxh7VB90nnVsL+vP/9mYObwpRzyi0eVOMa
RYhWY2zRur3WHI5Jmh6sMEAJqIuEfLMo6YJGxn9qkBT2NchP+KSJ6il0KGTw1PyNqfc0Z1HsRH/E
YFG2DB/vAGe3mcFxF72C7x7vDG1TtrmQQqor6xfbIXdP09FubER710N5YHkadm/AbTpcbtQvY+l8
MHPsNIOYOJkXVmeD+Aq4n83IlSOfxqdUBv2DAVNKOm1BC/gx88Zeht2N/2RzNtpQwajsWt0WgL7L
/lKKD5pV0kmGsn/dNQG6qu33l/oUYq6lWGzwVUl7ze6Gm/CGkvEwL+1QXjVXplYGvdVFmLYzfgQt
eGiH+Xbaqragx9mAXBEf0yQuH5Si3HyKKBkADUhbjaXLRTnfQ/zlkoCJdRoIMlSrsvGHue9VYvLi
+0t45+FggWjAEoCWFxl/W2PFW2KRcgzx8wSrMlOEal8DyoE+pWWEtJWvk+zhuZdTYoTZBXPfC9eA
tYzgwGHw/JP0Msmk8lbMqGFq4JFTu+xe6vuX188CvNVLaMsCs4CKWnXodwUbMkFQ9LdaQ9IV/9Dg
dmlYo71TdgaY/pLi/ZfB9aECQ38NQpWOtTlqkzBy6pggLsiSsYTuMy02UWp+NglM9xBuaduwdmEj
4vyxWiZrMEZ6t8r8uqJ3wEvwwSaSSSgbVvJmZ5t1fS2qN5myvuq0xgnScXWda1aLI22DYJqdd3Jq
zRaM6stTryHGpBNlFagqO/BNmsYQzXJaxtQBv+ofa1Jdxr9TUgepW+JqoYMuTF9KIy4P993h4Ln8
zrXEPVMYnq8/14G5Kv4eG8AC3pzt8ej8KPhsUrS4NhDL6IsmR+vxK0cAj8kNXN1KRKcCncwfDgwT
eBjMjzAtqaXL5ikQNwnGzAcS9wJJsRyPC2Gdp7KcvAQHKXchu4pKv27LrF/F7nfH4fiA3OudAua2
nZVIeQTqv3uMZjcz5WhVb8Db7dj03lKxqk2ZLUPEVr6NUXM6ZT/ujba6Mzg6nR3ELoXxSE2HbvH3
ZQk5JPPza/DlgZo+mXWqwP53KeBLcvggvhEyo4sRaA/2l09Z8zC3wxylgK3jvAE8ppbf7D9u0qJs
f1PSWvqap3GW7K1NLpSL48/dwDdWHzg6PHsgRAv4T75TMz8VWwWAkgQmL7YVOHx2P9C7w5BqyHW6
M49ACwBsDkYuZmQ6J+3od2s/HjShAnsslydX2OJ8z5qo4xtA62DRUwQfKCrk2YGTkswaHghSmQBR
taKr8SiNwov9qYhd3MgRW5orLln8tq6ZvwQzU1TFdM/fwOf09DfD1ItsS3gSSG8hDjuUrOjLn85V
uN+8Eyv/9GODnH4Bft1LPtKrQycG1PXpNBG+kIBjhak+svQ47jQPHL7Rh7L8pE3ftljh3MOwuCgN
D5GzgRMkqn3zMUzXMWss1L0AkaLwvwtiBBvr4Ywjc5AXqulcdtvoaL+mG1LLgRVWdWvDNdHOylc0
KHBvrfOpGxFtdAZc9kEUs1DGVJrS+ii0usFUdxqeLRnKlxRe2WRbqOjkeGm+5x6Bkc+ZF4TMNrGl
UhbuNEAQAlW+G1fptuS3/QTGSyi1og8qLJqzc5/XhrgSMzbH10Nsqcqcq84GxMcHJEBD7x8xyiEj
M5A0hu1oGrqBR0TALzPDwOWC1c/bMX8hOl/9q8Qa1b9NSr6JMiSM4byK5ozfn+ET78wUE4CQ71ho
VcxjF82x9819nuhZw3ZIwags3QKzwfA9nOyqRCos4tJeF5ALErw+CuuFQWyrkTUti3PrpC/Pvns8
qq0jRFpPe7WVj9M3KcZ5J9VVVphooympS12S9JCAhWOA190Ta63mmw5ppbyH7EgTx+O8Z4oj0BRm
hX3R6rOEmK5xp/s+xpwiD6RE7MAZ5fW5kiGAjjzhqmg+znhEOKZXpbKOTtQVaOmQjv1JH5akOr51
D9xkGmkPft0O/C0HsJ0JMrMToVfDkPoFl8ymiZSxDEtgB3C5WIMf+Cg13MOM2od69up9mkEaxgMW
cLZMaFM/cpA77KbjzVA1mfxeOVzjvMiUivkMvOBwQvMSAeLmHk3SzS2R7eTbtankeEa8O6dDeC6X
2t4qabHCsOOwRyfxPqvCU7mWzxxETEgi6yBU46xUH2kh+/co/ZtYQuAxPqQWWKZGQzjI38+Fh26e
7xD0CgFvMN/6KTJjsQQWU4DOLUQyCxMnu7DB1SAti33jQRtUrYpXUM57EFqhh2H6xLH8UYTfkntG
GKUWZZ4y1LsS6PoC0QS7aJ5Q9s1NCJvPZLIRADzy4mf94Kq85QXbAAJbGGkYE93v87w1cuu0puEz
77o7KUqd3pKBAeD09W7wzwUV+GtWOyAMdxOcTqGyEm8U2R6rNjmOJSZobsdZkFBYp1QlvfxCYh3U
MwG8dQU8+VVNiTPnJENAi0OmPyWyHWd3JZpDA6LK3aCfOJHwzZz7AOp61h71266rBJVa6gKcjN7e
zv17iSXROoj3Ub9bP5kzLL49kv02XuGuRHUN2vDzAINYEJO6DYjr0/FjpghDKk70udIR3pv9ybYC
DcihfXommAAazrKPc0IW472hx+cvWkN/ApdqcY+hgsg4P2TFFsnk1lKzu0j1D5tywII1ZjMaOCr5
x+WG+C22+KT17heQ5NFoiNM6jKqyf6dDrhi+tDaCirHQElxtLKK3dRTEeU6L/sY+3fWFanSb2WRN
c2B8XY5xlaQT/hH3wyWbgWJxjnkX7X5E7ebnOjO5h7KS6eSr1yQwkQATDk7JWbjhKFFHO32SSRtR
icE2h54ICVk0jr/fnVVvxpl5vBCwQlVFTWiX5upAY4Q8uWz7kY1csQMqS5vmM9XRM0m969FhQQxp
qRmhkClzj1DSAIDODxTob/MBkeRVf0qgXkFEcGACax8f0+WC8oHLfCuvFvoWD2ZyEX7CLd3WdIPo
bbm94ijjz5yZ86S+EgOiqWrPqJOODWNbMjJek/efm4efFyt4apZCK9wpD/UF+ES0nk8/l664jIGu
5SnogkLptfU9IP+s7Qc0CnPACdmlCqdar3Hok0dL71ZZiIb/M65M5Iy6gbAyb0NcMgbq9KQMZ/Qr
pkJKrVCmyvOyXmKZcr7SEcPPZz/tARvbERL9m06gTsxzrVNYDVqkKqipLexCEniXpVi+6pdsmJ/E
aFOf6uDmN0s6NRtUEHu3srAYf5Ggr7JT3LIlENxqvvHpvwNMXMizdBnSZNlzmqEUN05BvcPooOQS
G4tUIDC5THJVgr8pDhQM5ebaN9Vjq/CIcXFoZT+7UXPFcUBRu58SQPBlxj5Bt/SnvxpR8cgjfooL
WWkCn1kR/7Rq611WwQVi+YuxX8B/PND4NKQ2SsSecXZITu9nkuCg/Suo4/5yvhkgtTEC0foG8F+q
KlxkC1EOtz+QwD+2RuR/NyMGJLfBCllmUIbMbRYBAR8XdeoNKOnJ0qgVif/tv+bF+XncmgoasYn8
jQl3o1tB1Ykpu5FPG0VjamzJ+dhfCn17FiAy7L4NvpcQKFfb+TX1iVvcWF2z8pGvISh/vXyrX9W9
SqXuwJtWyXX34bUxtQSGcM3i+W11njs/NIlfvq0O4C1q07bIGF2PzjZfeIbGxydDCnoiya4VdlSo
X4dR2tkRkRyd8AJDlZ67H9JnOktU+VyhozLaDstqX7nnJPTxb2OhVR9gMRxA77wwTiScE2xv3GKL
OZMG64S2y1u6ouE+32KahnNaKj7rs0kOUZfa9Tfpz74EIEXnfpXOgiDOttu9I1YkOUo3S/g/Aef0
lmb3BnSghlCVndJmOGRm7biOlqXSVBEhOFfDP+4J1t1Qw4OBKhBoZz4KGvWaxMHGg/Uqz7EgYaI8
G0nqLZNgNgQWe1vgYUWFaXkvjidd6f7J9VrUtEZzkTt5d+7T5zOBILkfDPNGmDYyydLTr62JgDBS
vUmTdEv4ayoYeJzycx6wgHe4O/T6aYirbJohWQ0EUdJqqsqgWXBtWnTIqDGjT8yabE41LDMBaZhy
poCT/N0cJxRFXuoTLDb19jTHiFOLJfchr9RrJS+SfhY9/4f6tkkeI+/KFa5PwgwWky+hcb8yfPzy
AhJEgtp9unaGTK4mEfvGAevLXe80inSvekVftPSDrY60gYX2M+NPnreqUEWvBIYb/FSO7Ii5gIEO
tg5JS5+dGt9Q0PKHmFDVBcjO+R1agL/Fsg68m1CZ5V2al71ztS6G2zXDATx+De2o4dccpE3almCg
mdf7UGQYJwgqZLWm/BPpR+GSRTFVIQfXeLfAjNHqnsiRBWEyjtB/MApebik4bVvRbYKXJ5EyMCxf
fSnH4lh9nOgu7887RDLqivayYZK7IIJM3P7ayKfiBXSWlpjxAISsfPCSgWVdEZE1Y7/cIwn0leW1
tH8+PlkFbtBPJU0tAAhLOhw5ro+6k5z/iONyPvjDmG/9R2XYKzcsHNSEVdwTXo8zzxU0Glb26S6G
XN7Nq/r6vHc57ADEC6ZPkn+IR8A9KUPr6PTMgoffO7+E3l04RWq5aKDlFT7mp0R6IAtRxVWT6JQQ
VmUeHJ2tdjrojcx+f7Ab5qyzXlJUNUWuWTiOBw8IqodnnrAssFdUepyBVHPVR1PikPiN7n5dCNyi
3XP2iM7QIn6g18tvdi+qiqmq3jvN3Z7Vj8cTpctvyKkyrHqbhLXDGWgztkPZOg65j0li4xNqa/ob
+G98rXVP4DbWkoqeMYRrOOsL5lr9XV8XWDoIVcUICR0WE2xp47djc8mcxQZ3Ln5PU9o9nekThcQj
h3j670rYH0CQPEC8BYO7Umh58Livq1u0COkoPWvYg3zb9pv3dHN5Cdz0EJjUHsBpB/FRLAdDuAjJ
Crfj1w+FsailA/gbJqFk73EoRhcp25tzJKpjxSwI4TMsI07aC42ncd62RaSmNGq7ui/zJDMk02u0
pBPiYvvxnBobqQlZQCp80izh5NGbrlNiUjTgEskbQCORE2zmv1DP32ptjfRWJx7sSdHDeQOG8Yn1
uO+bXHJnNq/Ut1WhP9hAWcSxQ4X4GmnYgJ3hHyu6gqgh6ifN2UT0nb12KSmdYLY9N3uwkqQfgtL2
+r1QvwZ/CIyjoHAW8UpV7y0Oc+OxL5OS8DvqJxVQ8bQPaAtUbOJc+AGppveSfwAVy7304gNR12OK
p2z3N6Yp4RT1TiAyaXBqSc2wadSDNE8k3rYzO+bLIXBPvxhxt68F0QtzKK7ROTrgwd3ATzaDcB7j
i27jPEuCKqWzN4DkyqABDuq2/zaxHzp+NRkqsmrZlYP0o0AjnWP2RZuA7EUPHJ9rqlZC1e1yvT6h
lRJnLD4OaMX22t68KaMYXoJ6CR49SsBFj3jV61AQUiRRg1VfYZG0wQXeUSYrO5yuUWe7awrxRJmS
yB30AlqIsgI+VgIpa1vcdzuAsbbSlp1c/jLMTteYiEYHcBCDJDs0OcXmLTj2La4Pwn4W4x4vC7bi
LGBr+J3Os5LnDYWRTV0mmthPcTKW0W/LiF/X3yYQo6+MHioH7oEgc5m4YfTSJTeYkcJs1q/lf8dS
5lm77wqG1yY1XRAe7l51owJzxRW+mPFJVdtHzQPhd52d5SUli+T6UH4xMKNU8A72ajewumCkKJqn
jxfohO9zcouOze7D9plSxBahZXVfgAQHlV/TjBPZmU2iUMfR4Crrtlu0vnw+MI4kxQLncPv3RiAE
N0tlUm+ajx+ymQKa7t493jsA8r/zqitXuMX1KHfgLNL6kGkVROlTvZEnemXSaDBQxifvEKdsNDOS
wRICxdNjWfTudEpc1PGK1vs59J9647YJp4t2Y56fnilWwia/FuM/9VhD2EbnkV/CnOAfcwyYmarV
88wHJeHy4AlhDt04Iur6Mqm2aiBp9rFPmojzZEBbM5xZ180IBZhARBdnvfEUM9+ZGSFCT3N8tj/Q
QwQRyPeeaHbOdYSUkGX7h3u+g3SKv0u4+qwGDZr2FhJQM9q2yEA1DM8xHqLKVOMtcsYQDOyJt0FB
HR8lPaAX2PRM36j9HUCLjb+nqCE9P5evfVlQUuehjYpj1R4JDTHAhfWJm/y8On0BD8ze6Qaf+Po3
w+EzpffnooDfEVdKKn1wAPmxtHGN+Jz9mXFjFWwqe3hnMdNYViWNssFSVFh5445KcfH5yXv6EVNS
WqAMg3IXdS5+zHDLdh33MNic/NHQFkPZn4su+q06EUlYnDTPsXEPMiDmzifPU2TEmbOblJDRBfJl
qOydGvaey44+lcq2kUIzTfxWOtt99CAYdrR9Tcg4NzIokeBG2FtCwmCSdTtbXTXkZVwz0/LAYy9s
8YfZNPe7sikh61wSESRKuEkJiDVYNob0hUYKLPOeBy/4QM/5HBxgbfkpVSNC8J5yBgC8hfPe9nX9
clesuNUH/zy5WQ/kRBy2kKNIDFgGrytjJEiBW7zGuMbR20DQKZlS9uT2V8ix6NC40zekogsyHIxZ
aTDWQ4p0cujO/tMjPK9/9kJ4Txm3OoWmqA9eoLxu8+hNqmzlZKZscMnCXuUJAa2tkOhG8DW3VSWp
Its4rzL6t1jQ+Qcu/PVbv70CEY98I6RHwSc3gnsQXR3xzxbwmqx38DHNsT0SPSBTMIBTOonGRueb
ajfNucgXg9sEgdMmlK/phtIdPGtpJpobUJDjq7Q8VE9zVvF6YpM0CmIV0/NE2Rih6sMkxtQzAEVP
GYf7Blv426felNEB9UENGUxZWvdlAzX/v3DerATu6ERWbYyAlia84D+1Gm3jqLxY4f1oZrYnlT5p
K0Umktg8gxWVfGP7DrX3Uqt0mddax/ZfaXueJN8sExx0ed8U0E7G5AJ/gIrLIGDWjMIFXVwvUdGG
gYKn6PaQCw3KS2QOIGdJgARdyCyE3pP2vxlZ3Wye0BZye0eDs5U6YX1yZftZ84sU6tz9DLDkklEt
v8GMwFzqg8LRASVeW3Hg3AOT5+zv2DkNQlaNoXx9JGAbKFf9zZ8bn1bgQTnf+ayt3XxrAZ56ueeq
6YGuhNGZqU5Zrge8Trldu495YliXN2UhczRFys46b8NYbvjyP2SKS9Ccxq7uADZb9zCLPBHPqmaY
GveIRFJcMFJ54cTWELPq5/iy3a11xN9/dWojiG/dbRHCXQ9Jhk5lLArPNBGWXQBCsSwds9pJF9r4
GAPmVetOhuOkyJKMFCFekB4LPYYrLPLzrE1bjiGDERjStDKEY+Zi5nq5HFMOhkHaISZbRh0Aiwf+
TY9OQ0ICTOu1kOJh/U5t0kkZGOx7+1knOXJIyGHOKU/E9Zypv6SPQQ3uXh+kadJvh2cbF33+S8ES
NUxISQbdkdng64dScC8Bf0j7XnHs9n/GgNwvxCqAZSbpasRBgn3RS5bf7ILrbo4Gy7uz7/noahQD
tYb0y7wa2Nv0ZxE8qSD/RR7BaXkvw3+QYERvCjnIx6yJalhIoZDcJV8zU3i6SMSHEalj+cpouaa1
ijwnS1hQdsMHyiHDdp7sYBUGLvz4jzOlDHlcYD9yOEqBP312fkNow4SiBTPS9T+XLGa2uRveApA0
ZiBd1giaH9HLG6cqAIRgteVFsgkDXo7ImWWivIQGL8cCt+V2rf5MsKPxWUPtIaR/SKGabdeyjMX+
33gpkpsylLQazEnONFBqvha6TblwYTFnM3wlJSJFNeWB7GtZ9XkW7S1dDjXiNQ9AYkL4FipaUTyB
xJK2+LoJcckhuhDPsVUjaIb44LBPT37O1NH0cpMJ3GNrHssOiGPlKkg/xkMtWerrYcJ445wu/V0M
mFU+KnBdsGOqNnzEGFiYrdZOS4Nq/HniJALwpTiDKvKLJ94ey5IX5khhzvVgRwADa15uEl04HoHJ
8YXubi7JDxqNwp5NPIekiJnG44bjbk2iQl/8XsD6KOiMrhzpzt0gGxcGFlDOVFlt6aXp9L5JizIT
Tjlekb77IyjSzA2f0mrKmAMuFKnaQMv07y08VuR3AjDafTaW6j0uclTv7YrgcvOIDcYwWbQga73M
cghjNaVpQs642m4G1jp3Mxgqs7MhU9K0PIWS3oS8EgSu7d60dnMm6vZxG/CZhlzqLAluvKWmA7Kv
RAgdd8py7CWCyZTgn6zu3kxp800+S2mp1KQ5uZcFxuDe5+jxvXG6nGeKOgTg7xg6sx34n9F3eCdJ
RPqIIcc8Mq3/6ZXTHfCwr2tlwpi+S877vKqpWd96pShOzUjeWErIlRagElf/Md/peD1F3VRXZ7a3
h9lErwhis8tt6FAkALhqGEUdghiUqhxDsA4lJ+Lv8IZGJWm+iwaWOBRvGBF7KqRiphoycCQ5rlWC
y1dPmg+yFY3tCtLDqaHTGVAuwZexlt6tNe1abkPt71UtV6xCR5DqgKq68IohWKF19xGahIdRL3Bh
bY0URvOUsQ0chXpPgRNVORCHoaeT/raspFuZWx4AGPN38RIk8MHD/I/jDjL7FuaIKaekK1mCIBmo
tVtWS6/H0W48yYssZuapGmMRio9kSWzqtvhkcY5lXRDIHl59QCppHc15rT3HNYYu3qCAblBKmEwW
a9yCy4nO1c1cAZWCkMM0obaTVs47TQ48xDe7Fzrc2BgZOwjCsvUPyNofua8fe9Tj78x2RX89HsZn
DJPV1yzKmS5Zr1uwUjRcwRXLAI8YRiJ7PQTV6ePEBw+YqdgtS/3tOu0yFQCpPfrta2r7MaNfEd3M
ZYbF2CJAZq0kTIt5hh8JDmDXaVSSaz9enCX9fzwdLtwaab0m4B5Q8/zp4KKo/Y44fYxy5YHsBJII
t8CmlmIJT9m+LE0/ziuZPrO4g4Xf/SEo0kgj/HZdmLQk0mILS1ZLLc75MXkFFk6OecxHkqHdKB9p
9KP9gCWReDk7ow1UmPMyWwYMJTFWwfROn4uSxO8Cexbl+B0B6zaTvLUku5UjodbkACUaUYB5qO0x
I8TWHPJfu1eA0pRZBzXcdODsGMkr8Cw4KjXI19yjh4hHfndYgUcYvK7/q8ZNmrZwatzpLg2C4Rzy
2pWM83INfGCFyRDAzWM7oi7uDSgBrt1uuSc8ono/ocyirCeyk9+MFU4o4HTYlcQINNm3lTo/T/iJ
f5S+qXSE/D9VZOua1fZQ8WkmYlreG4WEbFgT34jff1q9aYyW/r1OwVscGJMbkElpxmrF2w6MWfvF
zeH9Mp+GDY+lE2EBN1QjAiW5rsYXnIN3FHHMPMTm3DB5JElsT5IV28dj+LsJYRY13O2HO5O6S7mj
0Vj19a/mb+T94XrNB8Ulh0jeXBa1/lmEr2mlTDfyKSKmzuo8RMUxhdn+vOtvFnmCqurmGss2Ug0z
A80NhAEYmDomRPYjk7Y+3oikvzn3jj5fc4dzP33qf3YjF8xT++0B6XFLZBmJNtLISPU53mhDEeTy
BvlX/byEau+GEE/ARIEhL/N2UyKgRxGY8eWN2qZbZL5oDczWrlC5mJ3ks2HSC3lsAouH+iIhlSJ+
tiebqp58GqKw3lSPQT1vG3lEhFP4yxob1EZpXLAySq+etgor6uGcwMTWwl2fH2fnOf1dEYTE+xJq
FP6pN3dPNc5WqCGX1G4XOQAy3FcNqOHi6IIh8eEstgT/mWfFcPII78qMLDSMIwn0ZAl/dRSxFcsL
/W7lJSkoclyp6sqpRha6zKyCHIoMpXLXIW1vFhV05iktDUqdkrn8owlP4A1tmGpDrOxEFv9ucNta
CoATuLSHjRNZEbnuqzD2t5gXps18F3c7tBTKIwiyXDdmo/14DBOY5NCy189uvuf67/1CMMKQ1zav
7bNSo5stZs2/VuKdydsXdq5szDIhNWkyyTrszFD6/Mv3Lt2orRge9z9sOyjGSRo7kRvf7DSZ1FXY
KH+zW7jFCT/Z98HYrh6fEajEhxYeSjlpud2NdOo7TjFLCpY+D1qwMo57HGOs0mGAPo3GPe0qiC2k
ys1HHYauXDce7LlWkjE8jy/Cxvx4cX9z5oeqRcZFFX1K6xhdIEhFNPFRDEjL6QMJFqbOUK0Waego
S7j7D1NexurNlo+0mx3MxVnQFntXfXfOExdbzqR3LQC5jv1SKm0SNHbGsKM6gsfCJQTbq3d2fJOQ
MvHilcfodU+oUTdDMQvQwvHexsR5UacRkj+fsHs/DimAriN89lr3AX2EyPkHRBZ2JEvkXL/uOXSi
yEEbvJXCVeCJ7c2Yhlqy3XOEGzKceKQghRFioJAOPwwiuw2JBBaYUHukD6GVjcComYMV3dylSO2G
JIlHO6w43uZLrCkBOQ7MkHys2YEdCKMbBIHw84A9BNs9mwc8GhwlaKvn4vBd3oyKxPUB3Gstn1z/
8cJbL0wcWc2dxw9upHbDKQpCQLldCoJmhB2SwuiG8rvZNwqYaY7YPeDx6DE/zK/rKLE6KJgzMtGn
RHP6Lxa2ma4rf5BujYt6Rf30zuHZFP4yP+zgDt7U+LQGkBQB9Ku+e4l1AKvhISsef7zouta5CDuI
r9tg5IvMZFcsKVI/D1UL8kdGYPPCN4pvkjGuzS3QT/DbMU8yXtGUMgK6ZrkP5ZtcycnznT7ZcTHf
OsFUxq9/SRhCSgllBc3ci05IHsyD69SiP/Qh+CaJoKhC4V8MFus5HOrhEg1v0Z7v5ywXBo4lCZmt
cKt/BlbLWPhQSRq0LHXRRT+RMR5oSCOLP0F0CwuSEaOSRf1Nh2XUX1YeIKfRwVrcUuenF8uJe95y
GoWs71zIioiI1aIOD5Q60D3YZgz/XQnoCdGrQNIiI+HVGQxyiMZXRYwN1m1XxUUcRi0jVuMJSjHz
JiCMSt89nnmVasFKyR5LDCj8yURY3FUBsTlP3Xc8lQG+YQUtbdHy278Vd1/e4tmm2vRlVo3ibqWJ
GNHdXrLSMVaSUE8NUhrCLTdzVWchBS3v8uuLHrWFf8mkDQHvCPilkd6ulGknSQ83FjW6cTB4UC68
BbqWseHPj9TjO5InBH05KZxWlT5cx1PNw8fMz6pFfJBJVPbwLPSzdEiH++FnlTdPDrk3dc2z93kc
0z2x9rsvhe434NNMAbvYsOthw2ra5jPxoqdmVtv3ZdmFQuVdD34mX1OpBp1kfuE8xxpGNFDLsIQh
+yF6Mnk+LEhMz+jPk6qbiNaI/Kj6uttR1ah6RX98sjZfsUSdVyR2nLwoLSNtfNOhavpYiEfmaYpF
XLYWfCECbgVOsjeJOBb9nQ4lU2Y2ZhcjojjP/NOuwhPz14Z6Boa/CMkdCMwKcWEVZP9mTbv9DIDE
T6RoHZqP349er/MXizvCkhy9ZUI+WcGHtsDGARUS7+Nm7IJmWJIBjEEtqUIC5TSGb2XMAfI2ZKAo
6hxpoZUYhMu6pktfONhufbrPI6UDSFRcykHLvbcDM2Q/Ztj6QkXf3qvsmZNBMteGSk30UcOzXfXF
LqFjbaTgZU9aJlpE3d5iJxJzE0XbKCUcrDVyUoYFCXiNxibEQWN1ory6mqPAI299U0YUc6hLS7I4
sZ4FuzG+dj2K+q+/RdIf+PDwJQNrSrd4HWFL3b5h3VsTS7jNBwFaZB4v+91k5gokqfA1Svkw2o2E
CjD79FdkLSUY+YnY12Pe0TpdynE6rANqymcFNTFOLH67TiB3DJ8sTys2FSCIVb0Vo5m0fDf//OZH
ZhejmYvm6WZ4U/FqQS2/bzyWUr/CVOWEV8cGuWEwyrs51s1eFpPmNLMzWSPon0m3/ChznqoNEoaW
wNEKydmxRRep0l/iBdhTJc/0aa+v7Yn9bw+gWvepdttTN/eTkwBw+0qZZjIVqqkbZjJra49W6kYK
cIq51vJGAHFwDcb6OorZeARjSZqLuqjxKugDC/X7Ju1PJuF2rZPynfbhqpr0V8mQrCLkMO0XYkck
8hUQZaQ1i9nOSITdYfGvP9ymoEVaViPJBq6uTYH099BLN0cEObifINHmKESSAg55NFW9YqqIAgqx
OjusoFbCrxHtQw8nf0jRkopVMgDPyNvW5b9c82taABFPJZByauiZajElCRyN5jYV8ZnaZ2HV8dah
C/1A75W5+Xp+RwC8m5SrgWYvhoTSxXrrA7WodkQ6W1CocxXSoAcJs8dPNz9umgKG40sjhge40lKu
OMtTpTBMbk4OWbktCgZ7TZ06MUc/m29uqxEnlXR37JWTthMwxDMUn3eR20IBwIMMNxIHONofhuXA
wraZ4lHlSkP+m71SezuudwyacQ3DUmHByFxpjOI7MgyEjn0kJ37b+EscRsTf81ZvhR967IBke7gp
si/Q4EegFLR8Sp2t+uGtnCxlHe6EtviHc3UPWjNJHjjifRuFWqvGIZcB5rrELWuDLwRqQNcIfLd5
HSZ/q3FiUCFwjjdL+YXUHZpuN9rAWNLgy0TP2DmH3qqR66owFhVlJxFCNKBosEeRJjvxJkqWtytA
d2c0nVerbBuw8RaJ7VtVO2PJG249EKHHQIVPVi45n4+I51nXP12JDUnLiEdfk+7KmfcqWQLsD24d
4PRcAfEv84Oh8xxh4cguk7NZcrz7RuJtpT9tX0HGGOLFbS75gLMZ5vLbkHOwexild1trWjPih4sG
F9U7uUeiwI2ToNivllpXyRQLAEJxDr9v8iEfWe6EArlQs8FFuJxsMzRAQn4jmbCbaDsZ0u5LPtTD
iG+fhf9n7irjhjcuWFbOD4wwrKDx/lucR73oYnoeVNq/VA6XbW9gt3cncnGW6FuQK8U53EhqXtj3
/+TpAW1KGNv4qxHh6yS3VRiH27CLJHclMNyburewD7fiVZ8SvDz3w7C3fNxbln7hAbgKtUD1KYmy
dXwAhyyEKGIsGNtDIv6Mlst2y9gkyq2oa5wvnFcadg0oArAes7wPV47OFvqaRPYookp7/Pu5TBTg
LjNP6yM5ZtdGsnPMeXyO6TAKtTHP7QcNN0NN1dt7OBd8IKx2tMPgr7717PQAah0XugSAJDlcf0Ds
N3qz/4HDS6TQVHkeRTW7z8Ai8YXFStLpMT0Fv8F9Xg/i4aPydSMhXFRCXhL6t3Pqk1MszKm4F6jA
Tc8vXE7nRxsdNux2qrMVNd5fj4IBpCYZR+BGFo7flqTYQbtoukDMMZGN3iTD8YJDDVwW4bTg/DOx
TShwQf0q10/vHfuA1MFvOEn1xQp/0OcWc8ho5PGjYGU9ZPZvnoxyBE8z8Yffz0NdeXB5VOBvxlcb
5Qfu3c3Mgg65rbMr2036JzNgoQ87DnTgsMg4/HxQIn9lHqB8vlBjAq1fRbDwT6twS+0kxo58M0wy
3fpDBMG/X3l4Rguv8Pk354U19mCqZjAWnsO1+4D2fii4ERN5EclH/TZ6nFRbgnuYf1ebjw3qovHB
iCaHnQuHYQ9/BdJom9Ls/V7nEh0680El8ompORW0Q3P4cEnZ1UYsAAFU1D96Y3jcOCIf/DPJ724X
8YmvorUPF2etQ/Cv9kubDBZ3NtjX2deo4JxpqqE1JihgXrk3iZN9zqucGHqUZ4S+jEVb01QAQSc9
FmMhBSvUFmpCOStq3bhuOas+gq9z9JQe2AMNxSviv6hUdJ7sdwi0jgRk8GTEiDRp15bo+MwNryo+
4D7bd4tN9dq8dM4uOS8ynuKVOYScbp4CQ4sCofoLywQHR75e9pHwGlQDc2XyyzkpHNRJyEBwarQd
JO0OEIgqUK7WSOabyz6t4BbHEKAZcT3/UsOjAZFuDMUzghfM76K9vSMMeE2XdOEvRR2B4r2gPd+K
1ZPLvh0HgOoKrlDBZyYzB7iy779kwMk7e50b48fYsTYVWZv4QBl8KEBABtkVlF/fSXpuY3M9vT0x
DAh3sLd/pxJ+Bhd9MYQJEF0q4+v0dBoAumRL/jgMnFYuTtd8QrfX1f6Yy/Pj9vaPwPE3mWcBhp/K
OaxPLeC2TaDCIw32UwWBkzvblUM+WXb9PQfIxwCRyP+qg2zmjGjetloMM67GoDGo+rZTm4ukmEr1
EfCytD0QDwTNpFEWLzxbezrIgDHPzRp/TUEFkJyrlogKWdnGwsLHE8z2NGO3LWmn5wP10FF6nbcj
g5ocS75Ddpnmlx/vk2LAtxzZNbejvnjMcduiNq0UPxQUfmRnBN9ZOULoqfuA2dNomvD+6Mwc/LpI
tD8rLqOD1LIfM4CVsLVXYnpEX+V77SpuYjqlJsOeFAec8cBU6Etxoue4XOxbk7NdCK35DTNE8W96
5duOyxNl1Bj7g+vx/YSiJgp3SpDDJHv94V0fyGF4vTJ3QQ/kyDesEgnLPtZ4eO8X7ATRzeC+KI5T
B6DsWKKI+gwZx7yw3FH9KX2Qca2ZZ1ajbSbmQjUKRy0LxPlokUeG1B+iSpfVpGSIXS6Yg+fuku98
414I2/2Eedhp/6Bu2qKFvyThz6/6qE2N9lwYl5/xrPn8MJkm9gPXDLV77vQNXJ84KzZJwEIRv2Yl
j8WcvfNiuYz3wJt5HZBgYHqeAy7jWAb4adUNAXtBffRvUdSwyEtWgWuKBORDZo8q4mpH1gCoaeDK
3pfkf1ri2SOGL5vpuBsOLk9UeSm4hzJCuNVCh78MyoG+Ebmbz85Oyh3kmiqWnYevVbxUn9LL2/Dp
z1hyD/ZsvHJhzXpTbwwnAV6OSndICSS4babzOpuh+SOzujR4WxglPIBet9NiQE44ao/r2CSPfpAQ
6xBiJqCczUzxfblaJuNyIdc+KrSf/eApiQgrP+oi8QlncV0R1xLO0nWBEBbzAgRPCQa6Pas+XHgc
iVoGkwvqk7d78nNo3qJrED6P0A+FkByGNQl5YNdyP85E5rL9XAuwhUiPLk5fxja06mABpwqzQ9OK
Ya0E9kvzkp7ZjsWstQwEuzOgDsC1+aBgahkyf/H1+s950wowUVmZXSqQHTKWUCsK9UK/nDIItRyo
tC54AUdMP+OvH3Ap7dl/Bfgswt6apENVKIs7Y/qtxb+/zr8d+3JJ2NfGAldtZ7gpzcmjRXu0WQnh
jIwDOidxN4yon5qUd4ZiDmZWGmJ8REf0AJFlFJ9ol7x/o+b/LhzUz75OEnrb8B2Jq2FSU72q2p5/
WKBfH/nAcNGzyvA3ZwPad0n4aS6h8D1eVr04JA92be9F2VcxqWmY357KP6yMVz11z7UiZVd0eKfC
5tOHX29gUZUICbmh18nA6o9cfkI1DEkgA3GcaLIDQpEQlUdSgRp1wKmS6uZnDzlYZNnJNAJz0hNP
K325MBQBC43QHTngmcWSrixeYDhzII7SSKC43rxMrZDmQn5l/lfWGNo7ePBuLUoXZV3cIFQsaC7X
Lt0VfTq4ud8vX85GfA+p7KrgZTzkn1PdGr3OF4nHTqoBfsACj4aERzJ3VARo814tqX6vW4wbXNib
OumN1tBZMQ10xLvVxex0Wd3NuLc2ISSeAa7XlXkHrBgC5XkqTrkk4a3N8sxajaMZnLOVn+TSVJCe
5f8pn0izq5ntJMU0Ma6RBjzWxScOng8fMdNVTIz+l+W0ECUowwZ/7gVnm1yESNeQ1RyjgrPEZ11G
VknM4YAi5Q96Fd0gZUf8I/ROwC1GutYS3jNunVXn+U8PKR4aDyhlXdSWAacZ011KIneKLw+UAzNx
+9iIJneyKA1cnDBMSwqM2g3de9bIrfsE3um7NIiprNznZcyb+5Dfv2TUW5kG+eT4T+eJoZmE8fxH
cnkB8lkbLolu901Q1Sh4IWqe3h6dE5t1/aFMIssKXV8Xo43X97lizzFmdjxppCha4MtOgv6W1FQS
syJElU4iO9sdlFwe8NTDZF5cQ37ct7TVDhhPhiVtAiyBMniVHLdc7nfq4ImhCpcjMBVyQ3Dsea/K
1YzZSPz2gvwwGB6IshJ/ZfZPDOQwEbBnF/zk2QSWsismUJC/L0XpX32iXeTUD1Xgyosdkdl4H7ON
Aat3iLpGiZFBpG0ReqdG0ZaVvxscL7Ii2rq67Mw8Myh9uBSAChd1blQqJ2EgVh/oJynHwckm0CqO
DHbnf9aVk4ok2+2fvBNDdK+2sl4yCSPaLKGgudbK7Mb5Cv//AWuzObfFnwcGIQrVoCkzdvFmNXth
cYXIHvBc0N2r2ofOcU97gqp/OxxF6WPUS1vfar0e4jFYsLXriXk/EPeE/GFMn9NFpvF6U0TOvU/U
+RUAmb0Eq6oy/dL8kSxpp9mMAqvtpuvGV3xwiksvBTDW1nh7j71AatwNn4WoV+lmlDdnGtYEK3Hn
gHPRYDBMuTMnQ5PHT0e4D/Qnc99jS+Gb2uSPgzBtWu6JNn4cMhTnX9LjZtD/hvvWlHJ3wzjpMIL2
hhRWXQ8bjxQUowbZUO17xMFuv/UqSSNySxDxXQzz815qk2DqKizvwx/56IcwVrtUqa7YcUcrh2n7
WtxYWXe+/oCryqEh2IVCJEOTHR7NJtVYNKnd1Ttd0bEDv4/xETxVICSLSofeBG/yYSrobE15USg2
8dYcRJ+N/373H5JemYB5ey+y+4Q43r4OOQTqgEzmVL8IYE+X03J5fUo8Nk45+M/ajTAWJcqYgDhl
to6Ycoq0fH6R7cSDHdGl8LDRsTqLYNjB0CNtB1vhksTFGyeUEckrOvAF/0Whj7GUE67+S4W4JrjC
/YfpZO+LKAL06IQOE7AcXV4A9BhMNL2jfTrfc16StLJhefj7acevVB2SN6EkWl7hb+nrxlpM6kUE
zZvQdoNASOWl98DxMj27VpuCMgBgTzjAju2vLtujmzkB/Pb5w3GghXncW7SsWwaShXAtaJxgRejW
G1E/5woV/RP8pJONv3e0zCb/XbnVXYVxGs9LZ+3S0upG6rFP95xDeh0e2PsvBY55IqiGi786CJTb
Ht+HRaLWkrqUYCigWQQQwktIoRxAvpVi2z8JJBFgmV//ugtnqIG23BoOrDhlyGyTbVpo0Ma2cItR
KRYPlFTALcGLmxfuTMLZS+uqREMUutfroCudRQ7hWqS+Y5WrLWSP72E3q8OZNMFDvwAebty7Jzis
MpoXP61g4Gi6IbbhXnuy0XiHkq86VzLDp4kJeSB7fYYF6Qt02tGCd+cXgIAU7lb2Tz8Xwy0D5ReO
JxeMwQOeWgqQRqcZiwMQneboR5TcsA2OOu1Amsh/uLUfswzIeY1IJS/4EMI4iOmVj9+ATEbAh9uq
2XLQNr1LQCEx+dwGUhWwaHjNlFEqMN86Ww6aFN8EC5lxxDnwIeA+M9ChzbTF8wIzCIh+Stt0+tkt
b52SsJDNe1VtHj94/0H3eToV2mvCxlbjx8UQUveCnPZv6n9O45BuSbtCnsOr8ercHV0voCiruwel
PEyxBIU+DQOJBQh11kanjK6wd9Yo+kZ8ZeTWSA4u1Ta+pj35Pp9IDDYH/MI9WDMn82TduHxexcB8
X/qCN5YmVt7jKy1ABGPyBa0/mOrKZyuVJR3eQtBo6TweFMWsWY6W7V4s9+dPX7aJ1XQdnFmHFLGB
2WXcRnSDXrzKS8i4h3E/i7B7ChGcbkF7ePs6PfSi5LEz5rQ6rLZqlVlP8QUTBEYeTFvtmL1MkHZT
WZ/xRLcr7OicU5POtt0EfcsyFQo3oxYMRF6atwKPKwgaqKLAoB77wfpFF229NFd5YcXaPtuLBGlW
6i0zBiJ0RrnP8bvJR66mLcwX9gJ8vSmaiVXs7ljEn16m3HtqOTtRL5PPVS6N/Sk/G0g5LEmMWGj7
nJeJ5MhtKuYVx9/hhMT002PuKVnqRuEShP+CtG+bUZ8M/ajINHSGxxdBzn3Y3XR84TCzrMnqHIwL
7rdST0+Lmyi6zUksgg+/Ef5grPWZcVu1JZuxETXYEnPhT1g8CFubI1il+D0GBz/VBUOA1PZsaamJ
zVjchL4XlveBg0YaDpzn0zmnoPkclh5V0Y28gQrHIXn7MNt3yn3VECr1BT3Kmynr1kRUFxCRsD76
olvmWvo32J9az+aNHgpVvWTdr14gwH9XtgA4r4ODsFwgj8ZdezbZmwfDUVk13wgTyBZX8dc+b3rL
e6J2CWIi99QAgim1CcszIYX80lK0U0kuMBogWQ1tk9Se0qoe5Vw6ZP3X2sbEo/bh3DjM9eQhLpQk
GuFbB7k4mkyig/EmkqmhC235cN+jdbdzbyVzLraxgj8FOuDOc1jOHd2OG0K5dF2XSigVu6/qLXWJ
r2vQjhO2bFpATCt0kd3h8ww5v8qFgAUy5TgI654+DGQiidD+3G4Lqm+f77AXwMT4IreQXfWtsmi8
fmQ3bY/Ut98dA9fp7k7e/uA8P4LXAAdAGy9CMbHHRENZBzhWs7Bf0Z1HqxcH8hzNraTqCne1803+
1DWT/nptLI+uNhlJQlph6M5aqTQ+uuVJ2d1X0Y7qhywpgNLWDfFm8WYAsjMTAhu1is1er94r0oXy
i2SwL8r4NAX0LYfESbjxyEktgxenj/twRvsoYKi8OImmG6Ipk18Iw6QIEfzv/EJn+hM9Itp3mRrx
FrjuTsWWpTwZbDDCqTN6doKn1/pSIrI1qF55LCuM7oVckb+lup6ewfretPYGBc8cKzlAf5Kwn5U5
3nYAZs21C14EbOeq+Tkb+uijOeXGxanAsNtzhpIPXjghfVHAnH/Ezm1LPTUCm0I4IIYC9mQa07Od
yvlfZtlhhzxa2TEeZQvB7u06WsCWH8iu4vTKlQ3n01GDNw7kLDPBVU6YbllPJMDGrMVcN8RbKu3G
d64K3XJ6y2QonLd1ZSg01/d61rPUCaF+EI3GVZMPatPnM2cbly6+lfITsgmALsEm2ffVruAdbQE6
ZSEpsMHa9IxJlMhmAFQtoXa8SoyKWGe7uHBjy8yPwZ9bwk1CHAEcYfqEch9fCXvp5S7hduFrjD9K
s/3HR5aH3Npl8IS3jvtNskgzdbV+go7X+ejxUObRp5o6iNo7WqpFSrB9eEQRLdroZGMAy23y6tR/
JhgK+pHl62xZc8+PXN/0ZKrL826NtgzEwmqWgFzR8nHJxb1w2krAUVcX/pwcDHt6D+qtaVk+xnuq
HVG9uVg/7NvdJeRsZi59NMGsi63S4OnL2NUP8f9lRlqycQnu3XKlAFCFyDzx2cNGLQiTKRmz4DPw
uC5zLJqzR6CpnnGQtaUlTdLan7nlIuMmP4khpeYXiOyKbLj9h6D/XteS8feM1yZKuJz5xaKcVbnY
17DiXGCHohLZHUOWdBXpjoStj+tRRB8ewGXWD0O6iIimkNJeN0fK9fdAIGhkfLiJNkE6ernh1Kq7
bfw1oSXTm/ftTLQK5pjtIM5Kd0WqTApYyS2w75TQKqrlioSaA052qhr4eHOG1QGP4hAkgYiTPnqF
ocddwKgzmTIt3Uh7Wst1LWjy1I9PpEGwM/g51mbCdpcnGdaDI6Oj8x0a8JtfDcy9qWaQaL6eoKHI
bVPoxqGHcf1a/8qrljxPk+fKCoi+Rl+jd9q3s8SgSMJFGLu3EeAntVMPrdrRKZkP7hq5UniYRH+9
52fIQ4+95wM7GeY3cq1X13XW25oAOiTqAbsflS46yeyKswbbLlNfsQfWTaupdv5P/kZzC0pkwbW3
GQ9ENDJdDjT66XMB5nx3nkL3yf4hTW1RtIog0TAiYD9RNGzYQI85oplYn9hjDwIfvHJLM3N9h8np
mOgZVE9F8Rv1AsT4xtaDGq+1sCWeXWWV9wBgISDDsvkKAsJWmeCT+C6+eosPVno7qpDLBUiYAjen
6NKGOg5t2WGKIZkJ1BHcIqHwP5TStg7Vz8CfIKScqC28u8lXHGscoB5c8T8iDMqSf5l5ZmcuszV4
czkjCIU3JdQKpHXh44E8Lp9/kdgAWpZaWk9zS6DhhcZbeSFLYgqDfg1MqlIV0tTN8M4iG19FsysE
/ZuHf6qzhBdr3u04Kx1pixzNBR9Z+cGSWupytKau5Dwhh52kLWnGmLxogR0QvPnAX1TvvMeIiUXl
1Xb46vtMzngHsrFWn8H3RibLbpuh7oAoBAtuJSGDsykQtVCFDqQkhMs5qOMnGihh7VrFSwdtg/AG
9Q5R5ZPSWGez38i8TNFUwMvBHdL07wKrfz2DiknNzLnC0AvPKAiWmuYwjYnJChIdUZNTOfEZDYys
aVNc3+ks1YHZm343jLLPWrn4u6qdIjO/STxrAPT3xcLk2pXtSNc/yVSb7l6cpBYYGFprdvWAsDBu
h/WFe5HEdVT1iBHy4ukyqUJvQLaXVDW4U/7azGciYB6te+Avop74UDk8e14yiIIVf/aQNNcSnTyc
CrRZ+dPm/hDMZdGtP8OO5dKpYbAxW8C5PzlmPh9SdDmlzXM9YhirEhIgamkak7Y0UTtD76yXsJJ4
VNG7+IwA2ZEfggnqRsfUnQgi6y3JBnHY5BWBIxW8lAc/MpH5yoOOSM7XgCChI5sk/HJ2R2FI6plB
QhNAPAeF+gynG24UXCv+wp6gGYc+6ZilJiiLTTXfGFDmHffzTrTmKvthEr8cXrF+lGDZTWVwW2LB
CJBuT66XNYABI28VJOXfkMUUuoI6HV0A0rhzmBO4hLI9oMD/1G+SvFaQ2G+r6Hp481Tdx+r2/MlN
kkni1GyWyDvDbHV4yRAUYQKTWtKp/jy83TgX2RamlwjcDEyRoDdAKWd26wYNff/UoOVzT/tlWnXj
EA2tN1+QQS+zVZAR+vVQdN/sTTxfxMvSwOqhhvDmFSHpblExigybMN0GxnoE8BpWMr+Q+c9LH6cb
jfPOMKPp+R4MMWf+xZkCqc75Pg7U4AzFVxf0uubONfd/bfUhCWrpUX3jV+FzQOsefNEHYJwcBqjD
L4nw4Xpme4nGu3d8jpzGNOoykQ5olQTVNpE3jZGb/8K0izNfw9Xrjjv9y0XcLh1/NVU3wUA9gnsr
2WBp7BQAb4rwPmkcTo4QTnBGYaydC61wJeQuGG5zQORAWLe3fUQh5o+++ymnxvzz4c0DZWuuzcfB
dkXAJT3RddOgplna3BUHcySAIAz2iILT0RcYG6BgbQsByntMQet2HHO0Z/8vfY1Vf78E2d3d+4nf
oK/1I6p4Xa/2pUHL72ORpRUCb9WDXmrUOmnayyBMGOgZCa3Y0UOIkPXID160LdsrtZlEhVagu8AX
MDmYJfB8wmmOe+6y+SSksUFFQuejCZzRFcBGCehknmfqbgRxueZYCC34zRLVAYbXiejD/fa/kVTW
URstOJ+xig1Y0Agzk3kbK1OvpH2QO7JSSdsJR7i5GepSaLmY/p7EC+hvXpaSTztl2zngD8aDYCfw
QvKtqru8BzsFMZ4YHDSgeuRlWAiOeP4UJVCRa0H4DmVC8brM3NFjo4+xFQkg/Z/Nk9cd9rUMR0u7
qg+lqXeFR/MNObXtIgQOKZQVURdFNaM9RMyOi22+GwV5moFGB/SDsq6Lx3EvvDMO4IMxmhPScnSC
eYm14LwVIq0F2nuUHTqZCc1vruVZKsvzOAZrcLS4ELLL/q3oncjiAO9bMbIay+/Y0qxCYjMLvhid
Ece0l1bsIFNIa3fRFwV4bVc27MMzhvfosY2pHR26r6T9NGB+o3k6Kb/H6Lq7L/+k+z6sCqPDDfry
j3PcLtxj+hS4Yztpv24AqlOb606u+5Uf60M09FnHEP+Q9or5h74DMxUj1Hk63CFwLqvmhqti9RpS
7fraO+aR4eorQXdavx13Cgy7r5VLgCqw9PCtVIuoP/AAsAMmICQ9GOQkaM6T1VkccySkpkobSZp0
aVWbbeWaeVjmyzEZliS0kXp0D97oE2KRymcj1T4iLhWU1Ti6XeCq08TNB0P/BPXKw7ZQn/KFBPmU
Zg+op74Xwa7Hcw/9KMT+OVOjfOLP2GwJwp8z2QigQgmZFYdEyV5XyUjak+rYznxThX4BSUEAq5MR
3lQnMtQNrzFYT/tC+Jpz19wa1tz1JlC2R/zHrvoxzyTZVRx+GrRvPGYqZHZ30x4sPodFR6uPLUPj
VApCWvNUCvhckjf7ksLxwTw+ggf6Kdj/YY50gSmwyeTHgLafXlwNvUSYajrMnLcS6vzEfsy4moYL
nzB3cQ3v5fYsX3jCeVltjD+gdlN31bl5iJKOqykp7kvf89avSn0NhYpMrjv4ZFBD+VmQEMcDlXcl
iCSTlurqei4rZvKgCczEmy5bjuGL+QXHm3uBY6ZzRGq+IdBUWN6FYkLL8N7h1SmJ+bwWBsoxgza7
MO2UxvCcfzw9rmm17XVLcoof7qfUenw5YEwOP47vnG0V1TWypd+XmLTZJ+SKtMTMGjBpuoU7wigB
QW8hLH4Fe3ljwAJqwQPF9c6rlcB8Ka6TTuGlakd5U1GoHrE1+sxnuBoBEGCf+tESRmw8REf9Fhrj
ShPt9tRnEdBXmSrSjZwHgFCSJFO7bquxfFejU+voF9wzgU5D58o8d+7Gykh+uAe/0pwswjelUGJk
yKryIu6gvNH6GnIF3LpxbMNUBRjnJV5DDtbc6Hse5/0g5UCTH/GwWsBkhsCZ/xkLX6KsA+T79NLT
NP6PIrxipwm1peCdK07hLessalgNGF64jmDGtaYq2wdY+4vp2VlyPNyM2hRrnyywx9qKH3l+TtBq
/wfXUQM+t5IDsYgITjI543eRYVUbSP51LlF820GE3MDeBD2MeuJbqT4Qj7p57UQqayqCuZ/WFVSx
1cYAffeGONeriDxHjZjEfoXe0FDnTUgNqvKwgsyxQiryEGCYzLihR5+i2g+FXio/+zSMGo80siHH
WInpwB1PKkiDydp6Q94ShrUwML8S08ZQy1AKSdGuAZpx64El7W3LobQLVm2y6wWyEK/DwbE+Dldz
Gi7bNnVdVMbLDV1XnnZpsdgwbVJVLn275NkTBIcI+4HaLfdT5cFE67RmMCjnJzL2jxydAIvpy1qE
eRTnfaldG6DGe4tGuxpDhb5UMjx5pRGxJgjcmnvYTx/uPb6NEMkomkYRc3J8EPH38TYC42Fu5iG2
yCy+yme6FM3qNBUH1w2eyumacG8CS9eFO/zIfGTtAQHzD9zvX5O5nwc2FAMPf10uhyTvZMo/ccU8
0BDZ/rJDXtpEJbTxoZgN6ULGsitKqMk5XQ6abU/ro7OuTxfv+aIHudGFPA9iOFdEeJF+8lZHsANr
OKuVZJSNN9xtX5IEQjWXkxp/uJT7xGnBfY/BxclSnI5mnxlqdbntr3KC/tyiMIlN3kXV5nmSlg3t
3QOA4DCRZgujP5w1VvhVIDlWPjbFccG3OQkmL+Z8W0tBbfUA0lJ/dNGGR1q7xM11V++oglHxBqdc
AGyMG2xYT5nWAgBU4QXWo8PKgm9YbLQQJkoW5ER8oIwne2zHI3PonH9o8UKkr5iQ+y8+ewBTrrKC
vdmksXTRJnXaOuGqHVkzAy1QG7o5W+f2vLKP1as4KnQAGrPOQd7GiRDmByijnxzQHw991AHHSz5R
eZ2w2WuG68RCO3QILIsTywecr5Qvsqbhkj4egPW30bNjA60H2LdaoRsMGUpH0Nm9hx6atCX8Kvn0
UpaHITvBLmfb7qv49equKTz7kZb/gteoCbWDb04diNq7OlZpZzuYNc935GekxG1QRbr2Lqgzw9B1
3ctx2cuuSZnL9rZGfL6K+bFxLbKbd7OWgSyLDZoiMZ/Li9hU78VX1ili7p901JhbNRxQC0O35kEk
D1QkphSWQyrFY9mC73Fj6oq+xn4FkX2nLKnx6s9nWILC9cezV8ZpXM5T6Efn91OqE3mp97A1hRKK
uEkYTY5Y6VgxBGOul/wfUOjXCH33yLN30Z071cKXYWsCGp5Gpa5ruJQvQchIfxZCMKMD6IR+y8bj
wMpZlun7U2xVwwkRipKN2aXHoFL+5Z0VbfRr4ntORkLIf80J91NVWv3OVKEPxzvuDdm/VdX9qCVp
+7l0eUMs1ZNnA0jjC4folPJi1Zak/46gd5KKkbbaQIBjrk5xgmt6n6mt+KLfpvZpu5S3xIaEI6Nx
RcaPC8lkVNsjOFRO5VgroWdVM8OY/eeOX9qJYDDbXJfjt5fjk+OoU5V3Tpt9AqgXJfmxZMa2XvIS
8S2IIiIl4ZljofbNsIv7HbGqKRmkKPLK8LtcFFW4U3Z9xlSLI7wJhlztBvjHyqOGfkdunZGExLpJ
RIaZZuJ2oVTnS9V/RpnjBwK1/doKrGy7uVGbSmmMd7edDwf2wVJTEgVooMBXnm64ejKr+meeQ6Zb
w8fvygHxYq7/bcRz4AWRPAFLLfZz8DwqfNnxaBYIaI251qGlG6nXf0rJlAHbhB7pg3jZy9KCnVQd
75rIPc8Tfb/Srn69SJqyZGP4XL0Y7o+KwC7/Dxm5tAp8OzBS72RszUbQ4hQKkKheAa5tv+SNEaOr
5Z0NUymesNkUfVzSNTtNiLPwFjb3u8oS0eM27oGDvem2E9Chj1m5TgIG5ZvEXPj8tp+E6mW//TnG
QxhQS5tLvB1krq8CV2XLASHRE3G7tNhK/knqGb5engMb3oPHJhc4WdxLy5W8FYiTQarfkE7mlHI+
MtAk0W7SQrUnri6yV4N0vN44F0hld4oCCokDH4TbJj5IDyI0tXybssD2zsml5o8stslcybTHKdTo
lUZMs17OXUsjPBQqg6QYfPcSDHoBBvrX/JPVpnVQ8aISzr1FTclztyvNLHawQ3i2VZTuRWn4SFV3
mhdbb+KNYG0zMTB2lFRCakvyrt8QBP8DdJxJvamzfWXiGpLzOaz/CwCoeSu8PSSVt6q1M6oCkNc1
3gDidqJT5Vje1F+LpaexnoA8NrfUiGxiAWEUobqca3p+QYbEz3HhtqJd+mgGXQrUfeUD86M5vzDg
JZJB+pIq32DsgKZ5KulhdTRJTlNSmgWjge0IrttbyqlyeIuvJuM/3mvJdT/HOYNncXfBnSpDFcju
hJPnTHLjiZ6cRyF7GEkRheiQcWkwh0tj1qhPoqZIoSMmEQY/8CHlUdA0CNSuY9Vcb++fjjvBWqfc
xzgzene5MWvEtmgGy+Un1LRaEgGB3blwk93JvMVoafqyToiJ06tHu9kXyJxwx6m/JViV9OMjU+lt
RQn62effSxPhypShoBrKb0ukxvDxY9wXwyfAozAh0vw+/3ImSIZ7UrSvWJxGnNgrfQPXSxZm7yct
89HwMzhXrgrq3+gn/WmS2e5asRl7SuoKuPcJ8w7+tJiAV1IyZuyE/l46urb/5wPSdePFu/F8lxve
cYKiKxbW29c//7aWp9EWgjEgG367LVXXJkhg5vGFdVtFSkLhqiTO42HjdjCaIy9jRx2WNTyj4rLr
/CbzT+f+esVjg1WTr2jwhQS+VGh8zYALxdvVvkzwijt1HFKkPXUYUBNRHCDU8bxCDLOwmTYw16MU
sI0GcZnfQcTDcYqbR0zef3SVRCPkNUbNlyLqbKzh5OzQbI8S2LgbTyv8HpxVJ2APne4vcJDEgHjN
4UzytOAiuyDnonqS6ZlTZVWID82S0bIC1GCXS8+QRQn0Xgio00C5oqhfY4MlobywC9OmWSr3tEjX
tTCsVN3CXDVvG839P1e82BSZ3QCNUNroBMJZ90ycNE80rvIgvr4Le0nciWM1LRSg6rddHTBW+Mt2
RLOIsYsmpW2MoTnQKlGowRLjQCP1FRYqOrgwoOB4PD+LSohfFWgPTHJ22PXLd2zZuHhKF6jiw8PZ
C2ERGGsgazM7ocamqrN6U4ke/qw6RZiW8R4j+eb16qUWvwsNsEmQjYg+ws0nspUGl3qI5JVtL7a/
W+5GJYVRVX/hCHeDRLm3OGdv8YTzPlxFGfHvCiYSZORcU8H3ilDOCpFJr1RhPvZCUL10e1WwSgmQ
+eUEA6naxw9h23+f6wrYw1WSxvR48QEL3kP9cf5yJhIyiIWCywuxMxI1pGHRwSOuHnr9ATifuplV
mSk/oPM+tWvrhS9s4iay/11ZhP3TLFUZDb2uKxzvo1s9NzbvGRsKHv/OoSLhNQl+rDYI6Z2XJDKP
kJMxfBZ3XYp8yXKLoOxNm/595lPygKexCfxt8O4clhRaglJ9JigFwG6wlNpMI4cOTWssAjbcLsRZ
NPFS/5rQnGyBLp1du9LqeiEZ2EVxyk5n4ZhMvWkVrAaWXBoQC/e2lgx6kOY2rlf9FTBn6JltK/CK
q80GuO2wu6y0sXVaz8hNEHXs8qDx+Yn3sxjsOgcR+OmIFazZGQfEic2sxPorRqeHm/SqJZbjOycE
bksCt6h2Hspw9BHLZ6FlLXWj2toXKadwhXYamtRRses4KfcQtVrUp6xppHDjjna9i8By4wTTNbJ8
9KKffbg7oyTO3duyFhQuDqDqzZBVSLq4tDlYVOno/P7bBO+wcUAdSK2/drGYVU0sEAuEvuMkFttn
PRAndauOsE7G8ba/svujZ0EIYbZWMFqxryWlaDSZ3mVfplFO407sUvVtpc0u/FZWI1OQc9KnpvKr
cT6bHFsCZXmm8o+I262Av9WCIasZZdx9VwZAuMV1nlP9KQ0JSoemrxCF7/jhSHvTixV4ADCjuBpn
/jmSpVtM2yEPjtd4NWN700TUj9rVtgKT/9lBtPMt/i/gcVX0a0bg2uG9Ts5QJZYhhlnPZW0T4rlm
atQScZmv3rbS14i35tQRP24msQOZ5WIsRCBmX+caIPPtxbykEaO34o2n/OFbEKLeEluxNhgu22bT
1ZzW8+Bmzt0n1LCr6MHI1+plbcSsaI2+NeM1HdCXGl6bNCVf10b8QOF8Q16Bw3zuXrXmNHQAptHS
Jm+y27hpPHvnPI60XzP9DRq+oPaGWzu4fkoRkBaeypRxAIZS5/Nlld9DEwC9q+ytyzKEAQTxYsZF
nCltNRWrcklTL1nwdvKMZRl5z7h0dISQRgFPEqrlb/veoxhGCG3krQIa7l2BAtIEVfR0CRkPZ6lo
zB8QScLtUZDAQDztNQuMvuMLNoeyUj22xx7SkAWD7TPC/0cX4S2NtrAUc4MGN2pO7U1+r0yHPv/1
TzcG1HOuL3ihaqqXR3P2mVBaxnC9W6oX8byLrBMaD2+qlJdIiTDrw+GIPI7gV5UKZ3dZvltfcCSC
AZ19DFPtY+8UyfrP6b34tuD7QAVkWI5CHeA4ETWlLp+Zo9JOCsUcE5AyqNz1rtdqiojApDckQ3S9
kr98FKc96NSo5biErJ5BKzQiwjLthn96GNEJQTQF6oB640CsUF7PRiGZ98Q6+MEPTsGiC3gWzxfD
9DFMbeOAJOd9btVJtLzsS2Nj7/roZyA6M+B5ovOIQMQOxAW3INkpsQU8KPFO2h8XE3IVNutQRsv4
CeFAa/bzeRVhONegm2d6wHMRE4HHjl9eR7lbjz+uLD6QokMk7l5nANkSGnZg2jmi3S9/CCEMgWy8
Z7thwfUoQHvvPQuqr+k8Y8cfGAhZVfXdGW9SJMEVe6mQ9pxCgF8Yq0XeJzRblcXcQkJQ6N8NwGEY
0iUwfHag4C3RHayqeeiZq826ygNkx/SJzg4cXoD+NpeurZWFTTCU69I7U1yjT3gacTqIAjc7EWPX
24Dyy3lQrNYm7hpdT/Y8vf5S1LhiHpzJEJj6MTfhp1pa3SWXqaBSOhMcCkg92zsVzr/kYxoEZwU8
i0Z/qYLbyDWOFSOvp8FQ37mwB5rgG7kKXHc7C7IBjwzhK3NLudQ5s7SBxwXm/5CWe44ZLyUottIS
jWEK5l2Z4UsH+QDCk/dfNnRkr9TnDUK1ud2EyfTaJNAGPCuNKCgfy4eUP9WuicfwgIGI3VupFHG2
cLsBRXGajxXHVaGaD1IsxWsx91FvtTuU1GC8z6Z0E4MQsscaXRFv+hen+E/GYKi53MRnIAbyfJV4
vhOQkdLjmngikFx1Wom+L/37ssQy7RwXqBy0kbwJoAPRhKmlQCNKtMb90yFMyyhMAruu9C3i1u2D
eBtfuQyJohA8BCxkVprnz+oMO3ePt9mYOPWXyDm6EYWPIVNq9Bjdsc+10/qBl0rRo8+VcIlHlugg
Ew8olahER38WPq+Tm1lDF9GXuRwxYg7Y+UqaExYW0WAeptQbp6YRlFkZhMaqX6fZrhYVNf6+SQUn
vHCYbrz5rF32COx1tSo09PlXdHkTFdZPxS1g2yoUqWW9KDCHck5xVc0PzdZjblRuT3LaZW1zj4vR
7a5/flmRIx4+hYn3Q8gE3136dohhHKInxG7aZXIRp5PGjTfsExpjf7LN9x+KAkp0WIXmOgrq8eA2
a0igx9QU/HN4G+8MVsPHuzq7YZUf9vUyHCWfRySj96d6c5KNopkNgz4QeJjQj1eWqtIxEcadfwsI
7vum/wRymFjHAS+HQ2ECJ/q+YFmRxFum5eWMo+dWMdEelgBi14H/TmhNmk+sS6Sdp59e5WyJQRS7
4VYSlHjoiB4hp4DIggVJEXnrl2NgTpoY11b27gFe3O1fFcEFZxz+V+8tTmQyN1VYQcFUfkeq2R2+
iChp8kWyal6IylG4HrUT2onbUZ/GzOKANup1m34NwhUNjhXgsi4IqMzZRQcw1mwb4BrNNqDtMJkQ
bjIfSGilZ7v9tFgZEyg+mKwBedSvR1D3UBkacGLMvjrvJqH16ULUngmYDav2midUw+Rxya5JMdBt
jY2zhAcZDnNXE0oqRVsFprtidyM8ARt9tzoNRLYjjXnrjiwg+AJQ0VCkPexfT+/KCUxuUT0IuI7m
3QlTtCgZeZZEwluzh5Hvsl5jntMLgbq3RMwocFLcGCTQlbdRnvJOoilipuLxnCF63wwZw3qL5taz
fdhIINHad15TB93C/5MepJhnpZGfQViSy1HamR0jY1gcGSVgdHNwpIwJiJ4bg7Fq9yisUe/AENYV
VQRfPyUwv0GPdfsuDY6INey2aCQpbD1fI2E5X0iotaMZAlBkEtEtxdcoUMstwZk9EWK8iK4ZGbn1
OAQPY9DUYoM0YUPICyshSMZFWCdl107PXr2dNLxf/Bo2jsEWxwMFEKmWsfRS66GsJraiz8QuzUZw
jXQUhaemXVm78RgVIs1aDytLzQycVPMlbzmF7/p7ifbd6Zf0Vaac0hjvwoV418bBZnDqnDB7nwpV
duxGYlJqRavShATXqYUecKc342y3GccqQSn0ELs8AsP35JTBuR7qu5xpnmn2+VG7Raqwmc+2L44j
B9SPcN4ExIfQ+yWFKLD1WJibEBpdUlgqxAd+o/w1QXJBnt8H3sLcKA36co0TWaD6isdsSksGmoP6
y1AnUJl96a5xSkv+mdD4RHfgsageeSwwj2IIz1qztTHkOcB4RvV8TIBq1I0ML1m20/RocKMDIz2T
s/1feImTktLNy3Ks8PfPTGIzQdZVgUFwp5twM1JhOtdw6ZWJ91dgdAeXmTWMydsB2w8aQC5CRNPQ
RXmRPH0PR7LFHelqjIdhZBkzbjlICT53WppJxb6kDWePUPGB+Uw0cco02/tRQ+f7PhnwSSvL0z6j
FnKTWGzZwOA3vhY9IhP7Yhj9Sci9agTMKDOtKX7mO/ktxZXLv2QmEjXF/wzN1EAuq1f1R9Nlg6z+
OroX1VJn79J7/lorkkljYhJ0UY7ByK1LXCGIbKSUkSGf1wxubMDG19gDLa/8S5hIATGvVJeVC+0O
GeutD7AqJYQgItvbndpKt1IYEHFR5j2FuNp4QiFqCnLlwXlpJFzeICOxH4x6MKBbbP+yqP4aYvC2
ArQDPR89iuMmp5pP9TFqVx1PPWybBh5UpELnZz9LF0SCtBO1bQukrcBPCrC+sKOCal9otdPpG/Sn
nibLEY8784sUo0Rce6mG0LGtyDKs61DT6e/n0Ps3nOh/AawsMC8dOCO/9vIhWRe+qbU5viW2TA+m
xDK3lxe91gZAEUofWC+rkPAJqu9GWOhPO+JRpfNIcCKvUX0ZY1utoMRr7bKlcDWc/18bAs2tpOPE
jisF/ql2VxSAH/H3BzuDWseO/hLMOu8bpsgy9x8e72vN6oZQw2HtFfFgyKpGDR5l+QcqIoe1hjLO
HbcqMzF0OVpH9V7K6Xoy/UECVFKtj5D7ggZx3i3AkqraR3nuKIfjvdGeWyt8S8MkNJ1+nZkvjIFr
qX+JjKZZia45bQlIKUnpr/H3Zwuulr4Cgl1ZG6f7Er5SziFzVvALv6E+5Zb2dFxMj10V81goXKF+
qmc0rkoKvDUVzp7gypnNpSXc8fASHqX3xXy2tyMQ1ECRj05CxR7TjXZ3MuQTnAsgH7JTfP6yrPqm
LUlnhLPy3FV/4F8qJX1QWHiVzRkhKSMHfZqPzz0w5HilgEDqJ82yd5yx/Plm0zZTszvBBoK2KU37
rzow31jzQa2yZYR0ScKikcPsR/xL7QeRqxrGk9kkfGL4LsJk4MR1pvTD8oj/QXNDnh8ShhB9KXzB
bnch0lLod0zl2lb1RE1sEqKoLWEwdIl31t+/ScWjF+5MuSOH1AD+R4NDlfEIaDJq4Og32WawRKMj
37Bbwt9MQfoDem1UNb7Zada3hi4NDOZhpY1Uu2X3VOQzZ/oX2FFhl1mgNfzBjAhj0ZhL9wwkriDQ
DeBF0R5Kdpz62t2v0DK/lvBFrcdz83iVIDrkfsEIGc6uQvnAPtx8D4saRspRz6RD+WSUNWLobz5+
ZJvVvCVPVsDxkP0beQ+QyCuQo5j5tOnqUM+7jBsgSbqC2QS7sLCM/ZCmmR6ceb29sIukpGv+8ZK7
7OuhK+/5Z6YFy7Z8gGcswNolvkNLtyyqyZ/1DQTURZZ7oqyN7Vvhl1uxrfMU1NxkLe5eOmpRVITo
H7msSRH1E0Yx3i5Fk3Y5aIcwgCeDfTHO1W2+OE+Yzw2dJDesh8Kta3ipBuCnV4rFD1eK1TDsy0xP
Et2ebPz8l+s5L4Gd+N2Jni9JFFlDmT9LZqDxFPO6iovZB+QOsPAjTz7jVN6DHglTuJDsHGwAQcWC
iKy9z82yfpammndNqj+LAND427wBWIykjYA/i9qTOs9wZRSxtPPq7VfaHkgPoz1ANpQT9sGg+j+1
lbf1E9hwOvxaH00q3cp5glDXstiiB5BlggwaLa1bh/RYBdafmy8+5nbu+hkfZBQfOl2yKFh7eAmi
4BQibL2n+rfbBOqM6et4BFEb9xABX4r+BdQo2e2hKGs/mRI1RmrxFtBtcNgU7BPSe0Y8AqUrRuIA
WJBL53AG69d+64uIJ62bmODkjQ67oDgkNuH1b7DLxY4QsE4mab4PVorI9PI2C9SQ0dts0yqgbQCT
O13tVc4t4pp/wD8jDCDZOxgmjSJGT2/2oI0o2NUpdanYOnzclYgV2w+lAuUQGCx0z9bVRUep/3+h
0bQ8DNycSH+lBA9b1nP4OCQIxyGXcU9JU84TQgzt22o9cKloxMVJxNwJo972KraO7Tane3Un7QWJ
Isuf+fHQNaNWk1V0idEBqqIDn4j8nJXiNtQZ3iWfsH/ckIjgx1/syChhA/ivltcNBBuDW6gcdxqT
WPY1mIk8h3WYHc8yoJ41cyi7Zjk7CJqqfstQZZC+sx+mj69oGLHEzctHmicMDfI/uZxODqqgrxo0
XTSDbtrnP6DP6FjXTlkNea86nZRSgXi8GMm9mTwQD0VeVtg6aQ7b7Ac5fpHV/c/x4lbkECLa4ZMz
ZGc/GSHP82X9WT41cQ7kna0IYjlHLNF+1gXniLlzqYb+iRFBrBMgXO2X1FGsFdoreeAftFgzV0q8
hZ47WeurMJA9rjSsj+QJCb1ZsF1XPregOaGuyo343mz9sUe0XiUuvDOesFx/GxSA9fD8j2icL9jz
Pc84uzhttDNTvO031BXSK+IiE4LRKQeLSLk1EJ8enwNB0axS1ni7b+bnVFcrGGSvCHST8CIxqAdx
ZBNsfYmN+zQnI+72tTWMy3xKa55yz9ppt3pp55/0+YL7blHuIXgBdnhS/ijX4YPs3D4Cl6cwtVgE
utO0XrMHfBdDS7Ah4W/WWBPqOq8UZoAQClHoSoYPrJy1ITHGGpPdp85O0/yruD15AhSh78j/u+z6
MgASMGVho0721RNanhvbpJ8WMQ8jzQDDYPIazvHAlhiYhVwyJCJuux1LJLPTGEiBu3teaM8FtZyc
ZXeZFOSqH8N4sneTNsMQM8gRwg6R75bKqGBZ0iTs4biFS6SrmWWBaVuqUiUgK59uShfnDs/WVO/r
bCwC7i1EDiwrTsk3Hx+PBxLNMmxlt+4D8YqU1ONB8romzToeP5T3TEPIdKKHvfWLhqoHynxXnEWn
o/5kEt9DziuGsAmlulwdYijgUYNW3qRzpJMfqkdeY5kuLxCBpbO5JftQuyPIVaPlaJ7FfGH/TqpD
hz32KBfZp8RZHJL5RRC4DPhV32HAME37AUwwK4PEo+R3XDDYX7gBKcoHujbeIqL+c/oqU7PefbTq
OXJ6VQhG3Rzf1UhOM5WERu+RWOPAupbjm4VHMukHYD1DJZRXfvinpjk+g+jXPY0Fg061/xWZVWww
W2y4faQpDE6PevSqZcmNOz2YylGW1qsu3Xd7KjRdqBqzoCU7iqP1r/uigt2jurh+JXqfERjdR18W
4BLcthxg7BVgu3zfRwGIHw45aFUdRbQQx7H2RTryXd+GmmF6tZwr7nzzRqhf3Cmhmk9lkjZ92KWv
Enr/x0XmUQrlfTnw3NyExv181z7ZE0F/D+rbCgjOJxKsbQW61ao/URGOhshein1MlV4SZWDyuyQG
TkMTJ6MxviWeaI9z7VJLQzXn4PM2YKea0YVhkhsETgYw7EiL1YP9Bl9YCBAAyKACi8fOkAGCzqT5
Qfei4MZfuXw1bQVyhzZODJAJO0Gggvo8NIE9SI8Fv1vbE+4dLaqXNp2HsLA6KHMexeapW8PdTpkG
eVAJWK86Fzbl8XRNX6xrrIIcp1/PEK3HLl7TzBPwbSxKDZRmiwMgpF+8EHsRKozRj7UnLHJ5j3Ee
QbqXaAwStuNhQtAIAK1Cs9l7EpeYvncMlLiSjVmFewoyrbecx7zGoKOIxaTg7QUB+gpxb4NrqETt
oEsbQBCNS2sBbvY2k9c5hE9HnwfbWj1UnJ9tGUVrxHRqJlHO/W/gDteudK7o8xQOdGihvCZPbwUX
FK3aWqj+QGSOeqEQFcPpV1DD1bZccEpEJEoebHxRUwL3TvRzcrAzUAQ7CxC/1payz4cHQOGp6lEn
RtSi7Lz4MYyYhmw3EFNl74rlzGKeJtwatI/8iWBWPBlpABie3RU9MUYImdQQwTtdKA/xO53NKLWc
DlQNZMUTj+cgULxWC0Lif0mc+4dLDWiVN1XgRbFWDZBJsRG8Zn8qXzlCz28s3yg4y3RBQpB664Na
WVDLf+vuJWzUF7DVTqd0ZZD+PBpXOc10HR1F/sSQxlWCgz7wvlCV2YmKc8bSaHcHzGSv+8j60NXd
4jLwyCGa3mbGzPxoJow5khVNJ8awD3WmE4Q9t2thbDCi5foSbWsA52XOmAWZgFhnpw5rELoaM+rf
VehDSToo4w9G028edjVpPbe+62n3GXNL9vIkrSEG9kNMEF4cjR1GIq8A/d1o0koWf7fZbRzLEv6g
K6S/HcEbR/rdtACTcxtr1psrQqCV7pT+dNNIp97mAR7S61hRD1nOz5wxZL7FY5ThPFSKc9e3XX0i
lKLb7PchLHxL/gnFPP9qlAIXClrcJYHfpug53apwley+eKOs0/wEeyKkJoFQxzmUhzPmcQQfboQ7
Efjeh7zNk+6awvK9Y+Kv9rcyzz3H8NU15RLnRAkCOcq5LqgHbxjYK8bY2j00fIlZcwy9tztcLsEC
r9Aeb1PUs1Pp43qtPm79TN96WU6G7HdBC1rP8HaMcQzCGtaYkC8UCktdYygNqu+Dlu2fbb3INi5o
UrYW1ZHSDpaGd0ofipJee/Sb5SAas3waE4D5kwE9uA9UEfsaBsJKxLGqCLIGaxfB7mJYp6poogqg
6AYVVmlmcoBYKkf4kwxiP/DawoaqelnKxG6p2wXNyEBWkdME3DVgHFOFMW1wbK4/AzwQyqXwCqRS
iNC4WjuNrdCpwlICLx0Fcex+vi6Nv0wlbe7DjCfJJlrdeYfnCc5gsrJead2T+Xmz0WLjL/Ajy8+n
HAoqqq9zTI7yQXXTFNSZNoAii98ENj2o1Mlh+U0kUUR/DfUFMfmYZxfXHCGxw586rpGsRQglTPHb
GK0W1XJkizW7ocJF5byfbeuMWtV+hBaPwUXfZzFbTGbZ6bRm6kDndjMlVdrVpsQo9x21Oz4I6bgs
oA1svLSJ2jg9MQbCpnTEmcLivAL1wwRzR8GVYwW509uExmigEobZwasfRSfPJhWjA5noteR8Doba
nX8JJs0ddJmAuPApsy8ipZ5khcdkxOIwQzK1WAY5XlPvk8bMvO3i3fvEzh8j84rGva9bTkZ/ZSaf
4HVMTFJJ1ec6phkrgfNxZZ6pYfo188qxV5c+HG3tuzGs3PtprP2J5B2w297gMAjOry2YW9xMfJ71
m5M6enHV+LQuT0Fj9cnAIRIR4n9LeEHmS/035+MpJpg5H5WQbWFgVYK3/Tw8Uh8juwagiC4lKBf5
sif+yXd+fUynfAVjF+1hqgWrFD0lA+1PBBgq+3yZrG8eGg8JHH+FS/ybnCyngAgNeDnj9sDBr4cq
VZJBw/vVnhEI8Lj2LMUruDtvk9xjyG/2ufJnsEzijq4gWEsI1n4PCnvl42V90GO0/x+y4UFqi8xI
tq+MRhh9YtbwBMW6zzKM9Cbjs7NS66XUJjfpmvSg5R71CVuUrYbZgx73bsGEMthUFinICkcY6/Ty
kyO8PWA/SCmoAK6g0usPU0M92kIDObD/iGCR9PSAHcP36dzn6tqozuLCAE729xNyGSIT7di+3GDX
njnSXl0HYfn46HrVgD0C2sXlRianL8F2wrjpdYkf8yaBDmwn/lPBOh6Oc7IxbL8ZhUi/1bs8EvhK
tMbTzDsMGjipwAJiFHYWBg8z1P4q0sKqirsjhpsRkZyw1K0yUPg4tfX/OfDTDulJQJu5H0HV2tcL
cSlSpGrnB6DMLxdjm30dmjhrgRZetViwXmuWGDqOhcl/OBusAWl7bDbKOowES2wJXMVaoZsTq/n3
KmrgkEHDgCxft5EWer8LCIDX/eM+eeV1mQR2sf6BslCIvBrGetC8emhCi5WL8kUxTIfE1p7wodin
tZ31kduteTBDRgh6TpHYmMMrF41fBqLFMBY1FImjVzS3VUoN852CdeqC6Iod+psUT7ggC5lTKIPG
6r6N12Mu0AcaEXKZPQbqAZ5Qpb+z6HMWkInYTe4hH0xRX/T5n4EHcyjN6vx2A+2KkhXqIzDYV8ux
LFIKNFiVRdNWl0snlPCSNKA9iXy1whPAbJfUYdfr646bytfNRDeZ+RJwy1761rMfeoJbyjolUP/R
nAub+tixudbRY1WFYs6K7K7YHR6m5jDpR0yObOTFdbpryGSTKYOsQ4p5HKgM/O0GLNKHaeDJUeXc
f2ZvjcKhu4siHBzQ8mJ85u4t3RbMVA9acMDx4f8HA0qnKAgPpo0oRCnhp/wOXgwuYNZ1ca2NPcO4
Cpma7aHjltQBzNoDdw3mzRqPsAUTKNzq/kzckFZx4LlZh/Rqn9glns/GFDiZr4Ddul/8FyQM54Ua
3ayp2Jr4Qc5VL4p/M3sA1yE6T7acN2Eaqcujk7GPt5DnWvmVdDsJIQx7a8r1A3Y3kUVdCGlvfCYa
qiml7jc9SSxfJ+DhtqqoWhqD65r5L5Y5BSyQBLkAtGpo8uubEj/xFIR7e1i2GeOPmTmALzL6xfTf
x7lQKItTnl0wyI8ltdBMMx2fdknVZxIJoRghHMoaEzbxtlnwFgZg6AEXuysFk1+tcbZ89XTyRHXA
URfZZ+hJDs30ocnTYfH/M+fAM69g2sUD2zXApdfKDwcCU/yncX+Pwr3g3nxFK7r0TRBK9ExV+Uc/
bmfoeF9BjT9r13Nt6iyRXu1jmgIjLtOyulOjxbRkBi9RniHWPcyqtMdokiP4ZnqGRm5Pmkw2k8CA
dPzbWEPHWTxF41OJvNSOlqHVYhyfgSYDGmSbf7e882brdhgZgbBjlvN+02Wn13PRXua1axtx/ced
gPeeyRSdyRjT9SUMTx2ymNEcNlDnFYPXt5RbsDL1/0/8TXE+9lwumUnyIjEYOkICaaP9esuhyjD9
dja5Zda6PFqN/1+R1AuscaFL6G7taeXDHGNSGBhnfCdRVeWFWOjcODXTU+l8Wf/vYXmOOcK+lIIB
zLLTi8vbY95mi8SMk10TfT1GOb0F5kwiHJLlu4vYy0aiClf6CKsfbAFFhTV1bOwEV3qxWNyQQnGH
N0aUvZTKN/FCl4wX5NPI1QCLXet9n0B2oYCoHyfdhbpgi/j6aswEjwToKCV3UjK4v06rwz/nTAtb
XPw+rmqo0k1M9dpLfOZzh6jHWCMfsePg1XuvhXwYr0zyePwR7NOjYG3ZttHb+ve70luDv+79P5+O
u2RFvZCrkSX/dpc1EgqDIuUkFlUFCZtc3AoSsYBv2poXm4wEDGHs0iqIqTKe5KqhN/uj10sM/r5X
Zep5rx+cMxim6gCZKmqHRK94kEYm00wYMf9KhwlnWhUNTFDq4HyOfqq997fRJ/2Z4nkImpO+AuMV
sdsPf4N5Ht6nkmJ6T/01ztalCqKDR/D1O8wyZwLZf68EvaH6gqtetz8K5NlcyqyH7OKsTinG8HUk
WKB19BwNdB/pd/RSu2O2vv1q0d7UtG27Q7NCIb4u2189FhIva2dxOLA7CVPDrPweuVwfuIDlAPPr
1auZs8MDTtJ8j2pxS3WAuZpAtxOCdpef0rDZOgKUrJpefeshiACtmZEBzYopHJUCEHrsdVvBX82N
VO1JYd86mudFnVpOVRLTn9LJ2tF1huu8FIP7EE8D+rImamcKN0g8vO26joo6jYn0XYP7sUhQ4nYq
1ba9sMpSP8KibUYh+Vx2oX8M1gHW96c3Al/Y+x66oqJ730/mQf7hcZbkn2nOQM8kVJL6vRYjnAQd
yr0qMIKGRdNlSYfmskI8Wb+l7LHUCRUIhmTmx3s0WBc/NtheJIe29bEuh00ZS3LZoFX/7L0JjQCp
CnM2ri1YwlUory4xGXvTdY+7JdPqv39EcW3GHXAqEG+pUJDT0pH6NwINjtg9wNMoUeFkgnfzDpY1
qjaA989Rx4cDOs37dGOHz8NYj1pC1/VlSFp7CLHpQuqaZ9lQLTEG97GkKPmvktIkiCNhp7TBVYUI
vxVCHHK/0LSoVKFcN2wAQJjT7ejmXYlBMgoaGhXYXb6mwkiAz3LapqR2yUvAquPQMzHRBqPmDB8r
Ta9x/d7RAGdXHDBA14VJb8mJ0pQZCmXDZEC+/f3hVN/NaVE9fr38GBdkoYnSaVEwnh+8KIfAJTzC
UfjTR0Ik7Nn7/R/1km4CWOWTLjfZUGQnapFljgGmviVmJ8tNsTwvNNWsRzRUP1GpYM2IRZZoVsXY
ajVH9suWsFGznfxBWiCQ7ye9ROnhU3FBaw4SpWhkIBFlDZezFBXVdGgjNL8Pltj83Vob4/ZL0a4W
Di7D/bkEBVGxc8Ldb2zFTYtgfE/Tq06AXsXKMu5xzwChHha8Ck28xW2FL2cB3ZSDe7PPwCCtb9Rs
yuqW5JzEIE6PqFwVqKXjWl/4EMDz4SIoHK6pHK2yCLsKSYar55TNy8iQAkkz9NGO7DGAhZRW3LeZ
W63M5eErFMAsFzS63I2zs1vmPBKX5XRVHcHAdax4wNbF4A1u8q5FoH3U5obh20OUqlfl7zQvwY74
ll7x8Z3mRw7zxp71EyKGPlCERzqIViVyn0GSVS3PF9pwrvmRcli2hb+N6Tbvo6xgknxI5L9ZQUlu
Cr7vWHaVo8QCrnTAFNjcufumHKnlJZr5PAl/0UgBCp13UnAoguUdneVgvluti+UNE7Pt2m4inwB5
i/4qa7L1qdCEESo8+TWp9Y62MtNpEDOnPmlAeZvsjzv0Y6ZtsdgE222lg3UKQf40XltH8zWArkpJ
RyKKcpHXsUi9CxS0DCk1nRWUh4wHDrW5uLiWfXIWvh92Zr1EeNKTkySYSpEsVxhLiJd+f1Qd+JXx
WinBz/IFA7Muw99Dxu4R3v1zPk5Z55pARbJuTXZn3bIcpRK3DF9DLw1qR5xlNk3BRLxDGuQbuXd5
dU2x89eFajaXzpzI/w+iVuliK7AWMDGVPr9kG2ehfS+TtxRQAxgA+s762WM/qz70EU54El9GXKyi
zLeISUcYVYdSQMaI1S8RmN7SRmNQd9sJJtiORNubNbrAZNCXHIKaoGz77SvBAZp/DaghorlnvaDV
dpR8l9h1pk3bT1jZwIOgLTkbXETw54aM0gJ0E21uBhTaqdtdS19prCSZpxf6Boc8UzdSe8JqrJti
sjdOftRoZbPxfrUKSaMaYVzUuFsStrvSq5NmzY+IJfRLk5kSWBfbJjOqQPiLcCcLWYESe0p0NFwv
AHuVgIytudFp3o2ACbYziYIYVq2Hv8VttP2tqx8nXgfKDRl9599Q4mU8EPPw0qkrrcvXBZSwjh0d
YGGURSBTaPyn87me7QP09hLEITWN7rDHgUys7xH/PuCjqb7yIa5HJbTKW2Pb3I2FbAHCrYb3kvcE
BhwIQpuMQPySr4ndRgBWgRrhQE6XQ/b0QsKc0K3wM4jNT6li4LnZAYexzs1sohKN/bIWZzm87Nns
DjyE6CE34F7QHEsfHLG/ZewWr1aQFNyBfwwuL3tz1bkA3+nSI7PBUQ6R+KmNtOFjYkW01ZDBIIJV
J8jXty8xV/WwHqTtVBY57Brzqtdsc2uaqiQ3FgWQWGdKT8VdvkryM7ou6eKow5mWsEbkxBKC6CPv
/788TSuB1wW2x+5F1fhXQl4e+NUSdveuZiuKvuYxHUjmAS5AwBunll7HukD2nsWZ68AGVfjyf0Cd
lBiR9WMXa5rxfrfL6eUP2BOzEorHRIDxqKAXzdzOtDMOixgj8hhKdsxFegjGGswcasTKu5qRLBKU
Eph1JiXL1DNb3rGlXkvcm3pIEWvpcXFApWdpfODoGxafWiyAz+hQ2KUF9LeRaR1uDcR0/mqmpRFn
LYMwvceFvr7c/BSzK+1wTMhbVN2zyFeoxmTarz99OEJTpXhBymVYVIoLBiy+1Ga4c/qeBXesiESx
zcWgENaPtJm/8naMzIGqYrRtfOd/0SlSlJnUF/gtt8Jb2kyEmVHskJVqhKTikLl4OdWXEwcBKZe2
jdES74lFMXvCLd+LHWKIYj/OoKY6c0QB8evC1ppCoD51Gh0GZz7yvU2/GYokvEqw3MKcDC5y3i6T
41bIxDVYtE5dbEQHq1RbzjYFvLqbtIaa6FTBrEjBJpB2TpPhYzYRpdwqfRJIo4o4GUW7W9mtc4yw
yfm9zPrBhOKCL7eKjL14fMOGmei/HWxyZ2zeNyCNoBiQHrh8SI5+iJsBG7Y2rzqwanr0qkdrlXWC
n178y7iF7jnTTXKAiIm+4dZA9HuCY6aXuo1M2p8jU16Hmj15xAJ7uuuFmQGmERs0xIYE/Yj9WUr4
sAehDQUbq2kITzjlynVOigYhHfFNZ5GfKXpnraJb5PZy0Nu9Gqd3zYdSIlO+5o58ghh9e+VURMqH
Bi7j8b4a0lc5Pj5yO4V873fusQ356hDG7t21Xp1x4S/+lMHH5KBs84TONm5J1u5IIOnIiDh+loxw
PcspkKhlak1k3lsmLoNa1IoNYzYucP4BtJ0Rahgy4FHjHZjQn0XkBbxN0oJug29gDhKxLaK7Vetj
88XQjSIMGsy+UcF/uHtkYKQOEfkEN17Zcit/MxREAdl8o1oH6wNssBsYP3ajueNrNDGeo+0n2KJd
x3cTNCiTEWO4ztl+5SJmBUivE+/7hxWiE5rsM56GrfM1MNPiYJWPamHUb6sNgODivukyb7Cue44x
tYaJfwg3Yv1vdA4UP1+W5Y/j6CqwtcUugg9BB7qqbYeAKAcUNNQRAI/YiH0T5NRrlduVGffAaRTJ
8HROktdOjwN/91YktYSRqN4ZOV+Nw/3PEaA5dWL+B5ZvPgm+ux9Uiv75XE0YqGvNCvFQgvbi26IN
y1AE+qRlxHMRXZg1jsg9c4Fh+dl6lMFSkeK+PgwplNKZgskiBVvoOmpc+N7+bo7Qj+EnV7Z6uHtU
S1GEcw5YDGBnBNWjKuwphe7gpeeDidw9mbXeITQQT1n+OgP1jkTbTlAr4/3ciuZ0gm2HPo4qAH0A
4q92UHEz289rTCoy56QT2V6Pymbtu9yf01VupZqT7FpGDRYeOn7IyHzkDUimWlv8iAntbFfX2ZPW
yFAR8/fGY7fhT//Vmb7zR7ZlgpS+xDkkH5j4RPWveEmSMQdXOXLSpl26SAYx2jg4jjlp4O3t5EyM
ShOsuxGAi/j2q9AWC2V01vBD58NH9GvDXqGpxYDJUEUZf/S3UXuMtzRFEbzkxAmX6jN4VfgJdF+j
m59dKNYz2Cre+asrEbPAQf0krUIpp2AeBiVXWOq07arbV8OHhQx5moVYhxito/9YqDBkzZ4cLn2g
yTep93xN2V6ckgmjxbbbVhHdjak4ZMEwl2q62/6WmYU5dFNItrR+vIggmRh717rwlFmWX5zg5QTn
DsykcB6eB71XxssRkxXUmB5dQaVAWQZfqnuOya1xh+rmG4xjj6nW+gPcEdoZWDzDUDltFuxZxHGZ
R4IKIqDYUq3KJ/yXdWxQmgkRjo2v6Wg6bE63s2/wYykxnC96MQBgx869A/tg7Y3Y3fSJKSRHIFi5
PWGLqJMd0lsieKHTQtvAFAx45bDp8MXbi4NLzNV3lJG8AuFNNNnHEEiyeDJQolAUz3WvZ1W7Syd3
YcxCWA+L+2SfAa6PU/lsFP+xTU9Y0t+Wjd1tSac1NoHUfSTwr53IcVKSrUinX5ScEYghStqKDQkm
lRuo8Lty8sA/Q4j1AJWfn5wgEIl443aOS0SmZMkYIBGRw7WNCNjpgs7lF1tKSlb+suNUs3LrtUuN
OjDncUX2f3IsuSrjvyr1vZQ+caY0804ybacfvmURuVFOw1/ANi60ol5ehP4VOh7Xk/Tsx9d1pJsB
l621MZjnT+ubfFJ5PtKw6KPwoFjWFfFJ2l0pXjU+w37EE1WYu2ku0uaB9X113834JvH4HZSNCRNv
odeCBuKAO8CvpCc1ctbmtm1qceRUQeDIUIz5DzUyVStT9yLMKyn6zb1kAA3n0BOigjerJqBriBmP
phkstM17yZqLJeTxk7dJzYyKMBnayA0cuuLAOO5oPKeZV50/uW+E+DTQIYvD5X2A/SfAd9Vtb2YN
12deFrYAVC7AW/cHODnRjimHBEKFJQPSEhrpaqukO7Csx5Qr5dD9wK/A1TVlfw0d5Mlp4nFSR1T0
0p01FvuFt88E2lQBcbsX/p/eMC3dEjwDaLAtC19GabTbdjzZaHSt5F4wV3pLLglaUqypyiNMu7Ht
Bh4/IESsI9M69KT8qgFawkyFJWE2yGqSqXO5k+npfD5IY3E9csv6z0TABFog/Ij105T2mU4u0jlo
xkAOLjcn7mOVV4Z2t/vxPv0uS/+eIhB8GL4EGtKFl+6XzibSK8pkhaBS6bd/B0XiXUwRUx237uCd
2rRJ2ftm4czZCbeXXkHc/Inl0hbq4nHJLK2e2CorsUSsfAwTtDR4snLCtbc13GFN/QG8QkbxCmlh
elax1T6pBXbZ+LlRH5Qq0mbGBm3vE28Gomb75fwE7Cl2U7Polg3E4RNFI2FNosnbUXzooKMBRgVv
BpoyxbXhVqbLSYHqdESyq42N7n/uhA1KCBO3Iz7njlFxtuL6dRGw7wcaW3ZbGNHVV0oirLSDGb4R
9Lc/d3SOFi7JTX8YgKr/EAa7JneSwkozPFcOrlEabolIPDOhh1yEPoVdS8mGAzD3W9TeTfjUypdC
aWgZ4SWukAK/P8sC8fFFjImxoN85/5XOude0GiV+IPjlqIX+OdE68V0JTHjZfci3wx1yNxsk6bXn
gvgWy768gUWFjSImcF/OM6ThkAxeESI/iQXWCYa3HFhO8OHFrrU+YfqH9sFFnOyCx7NFO5EZT/Qt
hazMxh0sHAlm5svb0p05p7ae1ayL/+mpSSznmwsyjSKVuANd5Oo7+6i3Yqt3js6dYUaAGAcWxMT6
FrKWFtmmLOGxeSw4FoBBphT7ls2gTUPrsjO2/yVcE+ldcZHa1VZVNwcJ7TddnyTDOUapLgPSO/0d
sggsu1P9ueFUVou/CDoKzzOepuIWjur4WuYDH2X2XKHkOg5ooiLcna/2EUOEMx74fgFzSkXa64Qi
FMDAVye1XzRsyD6c0wN6ZvXQxss0TAGLByUVmKNfaRZrWikaBGvMAHhfYozsXX5ml6kvCv/90AP3
gIVKPBdkuu+rpyklbqe+Zdvx7lFsops3NnpwZ7TW7LTDTV49aTkoiWo44q9nSqVbCR6X+PRXtJC4
ryZntOqNZVDklMhAEKydI8wOdF/Tv3jP/D+7Wdfe+6H9PCSpSdDmhIVLyyUCHB/hFUHlKgh2LPjB
jpqew9x65kHBN3JOgdpY+t2ToD/zU1XHv1Cib3rvf8nb2dn/1nnYw058BMNLq3VUMq+5L0ZeaxzG
71ZpkAo8O0etEWgY0r5gkvG4tDsEADZz6PJDOqnKpGaSw688bDd0OVePQKrFyhJ8JhrAb1R1aC2B
y7vU3ccJwEDJ/BjulxDoUFWv1WICJ+h0267vPqiqhnGHceEa0hoUQgJkcldjDmomCO+J3b4Tu8ea
pPjMCuzNiKNkEJP+57iUdiym+9NCmbbOLzKZLiKMY0RQWx9g8zeigXZtnGf0K+eeAVO9GHKPK3PV
AFb4hJsklm24BjUVG1ZIlKRgzKHcBi13Cp1wB/xTCvmmefPZbZ4wWZJtSSSl3+4AcUut9qtOgoss
JxAobcFfG189oqiORY+W6vg8/ofcBu3BlZ7d4ylifr5+cuEHft4Ux4jtfIZCAREivtgFVZmlIUbd
Oqu9YHQCKMUdjI4SOnWM61zq+jbobso3nf70QSQaRefnfzLxd6+FXPxS0PhIgULSkrzCBPSmD8AC
34cV3fYXkRQzY0VmGaeWNY1964JtKrB48HVyE9XbWmynn99hswbesVHadUL7YWhi3ftWhiWMMDAE
g/a9EQX/Igr77v7gQUmXYM1iKu4Q9qrx49R8KUCxT6zmz4JvPYikfSNVBHuj2k5naJrxmyF9JJ6e
khRYcCjNlkTIFO9EyE74dj/F20NTfgvf2B+/U9ORvqMgnudXGYZlDn9QbssDiEmwlfOKd+dnWDgJ
AAAUBDTm5LPhlNn670ePyOxP5HSbrcPJYLNe4Msc/WXL1nYyfSU/zCkEf4xZ57MgxGHka0s1WaWH
CL2XMUf58LM0sM7/RjrNCYiJLoyQUIlrEXTHIXYJeB34rywVx7l5ZMWqkJDFMQycpnKRDo7WXiNK
XJy6aQFFCBVfZ9E6Cjz7UUfGdV8/zLtcEVsVL9nFEnBwXUXo6/PY3eAXX/jF4q2MczxafXsVFANz
xQoSCvOtZr8IbNvrUlt85yRkbjOsyWzfoDBvFDPL3AnJjPCLFRhHI1RCkErhN5+qb3rgxrOrDISB
tIqtZF0p0OK1VHeUZKEHz93pVe669f8h7/0SKdD5C+ReHnD926cKTNdm3mpHyn52GaG2TAT/xKCZ
M+YCH+SPlj3jS6rVMK7g+5vRSYbU6aWMVFpn1sSvhc0LoqEn8E5t8oxGS1yvMgkK+99fSQ5SF5ne
SPToOwxcv1Urva4MM7ZNdPf0JsHsjU0wBUk9+RE+pfuRv7KMuH6qb0qM3rdOcwXIjCN0yj6DGKxS
nQPjF/LpaQM2IPtxzhr5VbqK7kgus482To0FhQ4meW4H3x8US5zjeUchBPhLLQ8csrWx3zqqTlJv
AIb1UVmYLvxUdOCpUfvFsFuxpYb9fDVUNjgdberGixYY4/LxWnvWP45UKeFWw56+8+e8er8wU2hK
UysKfpbTPPK7bXVjSrMJhfGvlAJd5KQgFLCJompuER3QTX/NQ41yVD3PwvrXvQMQCROuSUmGjtbf
Yh2WEjtunHcOImjkW2I6bwxHwu8lu4a9uQIoZC0Fu6tVM0mAnfM+ZVD6EBPPCZPk4kFirJVIhLXf
qSuSY8LDd5wAttV9+bI9griX3cqAHj6VHfNqeiwy8caXiEcN1MzBKyvM+dE+Pp6n7u7DtKyhMXvb
07/YJfHNZDNJv2SAm2j7MFucG/rLcQbapMMhCJEhECf4KZVvRZM94BPW+dWj3T/8sFAJfO8q74a+
OUO6ebK0RIdWwqN0XCa63S86hFuAnTimpPHn3lg9C84Btp5P4tumdb298dVH3W/tWSeoGcspwj0J
az6JDpq950LTkjJvSUB1WjhBesUkUrntZLhJknSkQ42WiUHmUicxB/7Z0hgxNWQx0OfuXIzcci5s
GsyO8vq6BgRT3OHhWV/AN/6VZGuCGuqAjv9G9D6Z/7cS/ncOyCX8qSjIUbVYmQKwlrvL5N52gFFc
pZZF8wGuTGoGX0tntgq/4toHQePcj/QCmSVbEWClIz1h0ks9BzxJhuHvUEdTZCU8ULPuKi5monP+
TdR9fTSgZzFAhUi1SWVRdoSYkNdU+iGwPnX/5EmvxCAlnSjK4tMSpTdBwjCZPNUshIS961QYjYtu
aw0U03G70YGm+V1sfD/yapw2eq8q1LCb7flcnnf+CNfY01XKmMWnzP4r1m/ZayKnR4RPKmI0zGiO
wPR2owU8+uFyWM8X1P2p5pU5HerMRqBkhzHXLHyQltUBL5g8FUCzgzQy5qH1UJHWzOrRBN2lZwOW
QHNZfRkfBM4DLFMZP0OS8JbCynWmdpfG8hEtH7Tb9O5kuD2hxPV2YihUJUj55wv5WsA4XZGsNay0
N2K6Mfalyv+z0/GDmmHQMoGd+UGXPnFB7iskRtsgwJM7fR/dqb0rtc0dno8W2l/3zr8qJR+6sAEv
2eidRuY9AJbuvsRDgllLysZ5JjbRZY0X4uNuabLll3hkNJCKLf+EBTfcgZlxgPH2mvDjk85CuJr9
Ld2yCuPa6WWBM4HqyZXp2IMFOpC/DCtvukY00oXaxGBw27m/vUbeIN7/Kbu12uPpC+PMdQaC/gRQ
6h8IJTxg2Coy3K7RNHT57fvHg29bFAzGq9TzlZ8ZYeBGF4VT2TM0TD6K1yTsPBhJEXA1J9yRYcpv
tM12qqU9jkSWuP1VGT+b7d76RAvW6n64ukJ8K1ZS+BR5rfMRcByBI5FkNAb+EiiBxMXZMVz3HIUy
dPWSSSjbBHWOEclWy4UVGtgH7uzMTWt8N2yHz+4SJJqqrsQRz/5GwRbflPZ7SfMkwjiqTYto3h8i
xuXOqm8F7Vd3hlnXZ4LLUOyytsVnLEyGWfTHzFCiXqC2NpQHFkqTvmuYIEgArCLTRN+pGuOxJJFJ
YVYMZ3oAdNfogFalLpU1CgHm/jI6rpjdbVH2dg/FBnUFX0Qzkz7xW2v/ElAcznhOmKFW/gjPKH1r
yJ+Q0vN+q+R9jBQ5E/HNqWl9n+HdijH2W8huqCuK2Ofws1+d/Pp00qGf++w3UBeWUHAfO2nLOL4x
2zQZseTOhkxPCYaQwNt0+9Avt/UwuaJ+5KiFzFAf9cbebP7cM68wd+91zCiZfmFhEfhkcmJWz7Rg
N365wp+JZ876Kk5XPhyM96WTJ6L2HSR8t2n7aKmKEZYN0F3I90Qmqdt1ma26VmV6xo+3WIHj9uHc
5xnB2lMP20WZNSgLHKXvb0vZA9v4gOudlVRa4S7Dkn/qGi+v/9PHNk0ZVjckSrEchdoTfRHtQtzB
SJ5ImGVMue3JSUTE7SFkVrZ+I4USF/nSzXHGksKmqEHUcKUdf6LS0hT5J8+TfNsbcc8r8pGkh6ll
udvSd8yb0gIkhmhm3/iLPlcytIk9P4A3RX44xZAonf4X4cBfws/Bl2rXQE2BOpG1lQEBitcDuRiY
Pt9Uv2o4O9uSOMbnNf4OnyJzJZaMBOq+tyg5mmF/FTGAyQn6PI5p6dvdlGmsj4YjebHA8S/peHtM
ZsHi2QUKFKWq/YjJzABJpD6CU1OteP17q/AV45c4WCXBQGlE5rkuTQjRF+T2e+ndZhRpwW0vhiH+
np8eh/Qcpj36kUfZMwgjGZ1A5i5p50Z/PyUpmyLKjl9kEIHgCNbGiCBmQ2uHJimk7HSHVPtmll/+
C/exe27mRwIvT1oxMpb+5dQ5rj8LMibD5hDbzqcBIb1c2K2FkRt7RRoEE06S21Ls5exk+zItR37c
AfajmqIxoIyVvUtNp5RoLYM+OPbwLZFNA++OattPJI2BWTmQ17V3+0CqLiOhVoW+5ONk+HfAQbMl
ycVJD+qXt4es/q6gc3xKS2uWpHhwdWMeXHa73kBP8Ky9AOGGoSAYG+AhURlszBV9DA1hXWK8MLhM
V8PJtV33ICCBQt+dTMnIwCVPhfMFXbPOaEe1kBOsb4tUXCE0mPPE59uTQk3UORcxadierXc+yu8K
U4MG8PCzB5nhQB7AAG1JUOo5zGFU5fRWy6L961nvU4ccLyNhmV8xVS7C4EqFmAWK0Wv+hgnMBzBq
AjXc2EbzeGI1u6pdonbKiYgySBgfBL1Ax3US3DPqeL+6yxGzwkB+la+6yKM8yP83oV+q/WmSrv6k
xPrr/lZ8Xd6MxDdN2r1VaTm78fR039Kxo7YN7TctlcKok95ntjkezYqGOMyrfcMfnEhV3Z4chTf1
IXk6J/wi5dk4KstsqfcKQdxm+cQfBfJsKWyeAwyzwtVOTzR6VC8GESNoLpll2ZnOYfal8G81JT8i
v8Ww1MMsej2HSw577ToDExSi3ype0Ohbdp3D9wGHxWybiIUZ3ySzuvxuRjfLUFEKWz05LA3CHFQG
Yq2CCXwWSKtANY/nGSct8vlRB8z3g3HSLQ5PKi7lzst/199ySPIQFS7Uzu6p00zfrBQMbBGT82GD
NKCf/gGcmLnqCjyWJVQYFBcAa9xHjmlhHMnfYRye7osFW2e0WCso3BOfiu0hoT+LYgVCsKkYJu30
h46xWvtyF2NAy8Afb7xhWhvFKB9iDky+5zc3l0pVyN0WrULFIxWHG6y1QAEYuA3wl/+MxlYopR9t
NdDAXbH6ZBYzRbn3AqZLuB7kDo6egoncE5aThvSdIjnIuPJZ5vQV+aIJxdb2Qa7srguDB5qyGmbg
eUhdfrWLUS34iVb40JQLjz44bbJ55z/iYJbatCjaoR/8GI3dSUPht4HFBb761PLJPGmOa9uECwO0
XnJnP39FkIDKx05iYd6H1XZ1KZVv5IQZueP05fG0G7sfGVEckNy+PggAyk+dOFt1y6R1rKlE7eCa
wW24JR2FmUGw95vmr060VCRJZUXbaq82xSv1czWHQjMHEQND1RQWWWrl6ZSiXav7Gq8SIB/jDBkA
FzWGJ+U4HCgExZmoAxBrAu8aIBva3XR+Dv2lQHnNuH3Atc3biZ/l9z09wMxXo7qQi0IJrTQDwSJs
u+0z4k9QNp2jA/HSoRS8pBphmSQ/ABrybKts8M/xXKcaeIycqrp7qTUbDp0xU32VMp6fVp8oDbu9
Axvh7TCoLbXE1weo7W+G0gJITDPwQLSr+Ge/q4QM0DidOBjQ11VmU0XNcFFkq1LYmdVW8G2Azaxw
JgyErID5Osi9pfheIlZZHpcEoF8gLQjAdX0ShXwe/LxGPGupWZXvcP84tvfpmCN4nFG+IOKET2z/
yKGgpgXqT7VMIquWnRaBp85ZEMQewHD3qEWDxFhcCHsADwGKZjI5eySCoYqU1nrudaBgfLE2cdcV
HvOxg+NHdBFh7AfrQTPuQ3qyZujNxuKeOptr1gFHtlcKwY/umgVnOUm42DTO7U9qIMVD5Nh3K0zT
72KHR/vBFOSk8EMk6N5nGbB9gNF5PyBcehcaZm+ZVQGg9ZZjJL1WWGLW8JCMA9ZbMPoe748wicII
gf8Vr7Jbxq0fQPomZRKUHNKo9Gf7RBOWqQe4Dg+3oM7VU/euzKSgW58zU+bQPwqRCMF5GsU93CTi
WX3yQHduk1zxqnm4EpBQ5oUgFF4JyZZQhv3uA/u4Ds+TILpje5GyNrO7R6+6umMa3h+HRAubuUac
IY3JvqvfEgFoPTFvfSv4N/5ANkY/zGAuKbhKT56PcE3KBHrJ2smWqy6tPvujDsBn4dMVk1ocljAE
KvshHumszatSISKh/sMeF+eTzCk68Mwzb8zO0AwYmWBzs3NByXK4WjOwv9yfTheXLfUcxPXetuHu
nhxc2kHzDfoLDyfnAgd3W6+LviLDOCyovvtgXdI+YgD9nvkQQthSxH2X4e0EC5CQwhBEN/darRTW
+V8Dket+/T/5t+PMJ9CutToZqKmpt9KIuI63GwPnLtwgOv1qGGaqiAPZIrlmQkA9eKND6xusesZx
vSnl39xZB6jRsCqQv67y0GnNyUZY1kq7qU/jkIpUzsNhdE225ODXRcAi4GE8pRCxnZpctrEjuVqF
k6lGCRU6iN5VqonYvWZgam7ukVj8FfUYUWR/q3hwvllyNjdWhuoR2goTBNhpGVzZzIIFrdSOwdyE
ZIvQ5CcbhV5qFvJNPYxK7Vw1t7R5VNQUv6WPrrAH5roV0eJWFXtG2/7WImOENE5k0U7PKqAPqmLb
Lndqb5QpFjtY6oB44Ay15+ZOVQPTd5OSlfKGE2fenhtCk8HtEG2OaqN/CvDisuJqXovx5uLZACZZ
TB1PyWo7GQtOuyivNKtqH8V8vIDaRNnq0911Q3fu0RyVSAiiZ+GOsB/Z0Ip1COQmPvATlxXdXmI2
RY6zvrBjmHFC7fvNIf9JRIR567pKnN85aea816PP9gv13sOLJcwWO5+vcPhfks4Ea5oL16A1K8qx
suqR4enm+i6kNsFhk/NOZrSKpMjicONbKyycoAcUbgSry3Py4Rr2gK5cKQL79lkM/BnZm4vAZS5i
QMKG/NsQuWUP5UTcXPU+ngQGS1K5P23sL8IEUOTBGD2bcF4sdMzXdjWZimF4K0Jm5GwKDqY0/Eqv
lNoxWIK+CBZyM3fR4hAI5If0lI3+BqWUrMBdAwmHm1X6D3LS4Co4C6bgGIQzNC0kP7AM3aGObrl0
0CWF31t6yVAWAuvIC3DCEkyQzJZeP/lr3dtVymHTzmZz0FE8d15ZZAMTtVe4I8qkCK9s8faIGc5b
/r/Qcw+4S7TIsLnonB9FvxvZ4uL+h3h3rPcEevmsR8bHuG8WSw65dJ2U8wQRoWqzhpC62VGIvfhf
qkCZk0ajAbYsFrmwovhGbJ9qHSAmlrdl/XHc5JLjWwOPdAvzPY4Icau4R+v80bYMd4+PwaKyqO1K
yINmlgr7IpwOa1fyEp+UBxEw5BTntG7AaIESW1s/dtWVBhymQWcHzh3Az1dkBQa+JiA14+aIGxwu
b4pmc5vgddEdt6p9UuqLPHk7gFWoHIRdmv4BsoCoGmj/Zis7WhWyolngFcXZ3LvKlRODtfB1C+TG
3LmgkWh/RjZv6t87G7wJXKTiT2mnYhbMUzKOJiTV6yBMy4JT4fznOSPtRTJnctru5sOk589OhFaR
ipwT5KrkLo3RJQ0lZUzL18K07ML3/nBFQAe3UGq6tv9PzCEHQkIp11utsZrVsn9RVoiHyuENSmgG
+klshCoPX90VLtXxvDVNekf/vXGhP4RJ8OJA71hgVuj4syoc8rc3act8gl+5T1dasRcbFv4Fb8fD
U0aRur75aF7sdMnfkfYeG194tqc5S6AwWf4TW5tsqTj5XR9pLcBU/416p9zU066lhgjaF2tC6TRA
DBZ6abJu5+RmqF0/iX2+MeJBT2912YXuwvZs4fzbsUbkj4y6/AOhiwUVDjE5L3x9YRTVI1hbPP6C
voxM0f4FPKS4mGK9i3QVqwiMfzskd13qW+FX1v5v5QLqgQrTVd8r5S0tbWIZHJGqjvg7Prsyhpi4
ahU/xPk3rJb2SnjQTqELXUd9JFkJEKFvLG6e9rZei7uXcVxLcQxgzxEzHwZUIv9peYwUa/c5lYb8
i16JMo2vOcSw19GKMQSQBOfg7pMTHN2nZHeqPCkBMuOxuQ5LGke9hG0XQH+68XqWRy293zTxE9lz
TBGmJYqziKZ4d3/3KmmZy80wMGWksgbFSPRc1o/afZqQ9ruvvv+4xDk8kQ/sTfvFlniFl75PDzjt
605k/dYkz9RlluBgqGf1ZHwmeJk+biwTSKBv8mt7jJu0WD1L4qI6DyEiXb5dnP3xouJs6YiB2c21
iNWVkSWNSfUEvsv9mF+ASOIW4LC/9fBxsmsGmT8NI9QGXOG21Z3HbGTcQNGvmE8C3hNEuIYyjlBj
ZQiBN8RGW2RG3YkhcczaQxROmNzpQ5fNptDWormfwEvlRTq9UN2mJBYMoM7BHf5FOSU+iKtxvE7G
RYxNX1HM3CK3Xfjuc0npqT7cM/LEB2T/kp6EmomJp5RldTLwfQqBB6QbVBSE6jZm81qizDSDwBA5
5WGuwc6ZK+r1au1p12GQPNaSKR8sWOstdrsYskRy8RI7illTv2EFraFIkFqas0md4Wg0q3oGCJg9
TUkmw2lMLNzILyCzMIh+fgNSsrl4fPv5r0ylaA9gCsO1TKPxKUcxlJoHVKpDE66JbrJlT3OQSImR
uERhD1qjRIeLfiqzj+RuXibAw8lgYEd88FJW7BhI1yLqOLp9V9+CLbUXKB5lDr/McLqgU7rWtwOC
lzMSjKBRHcI3EgZouu/giTEqMAPYUTZYp3oUbh2ITplz6hlQ+LMu4EmsDhKwP3W7vlTTkfAOYYN/
W3dmKEE6mGsbh22u614z0lJg7j3tanSBiQuWKjfwmcdvua8vJ/GwT9+CsuCh38m8IkjVxTZ5hHly
/9KCW2WJxy1g9RzYBjKdFB5PwESdr0fShlghYMK06UAoIEqaCYFbyEal8yswISDOhMBC5ZFa5RtI
cWP9hNpmq57MzK+U62LoSClbaWBlOJl9E2tGxjQfqutzD0QzlXODHMEw/zNakp+Wkpm3LuSmBTw3
pdz9rYCDr9Hk1JbEaQWpwT3bdGnBtTPPh3abMz7mk4P6UjdNcd7E+u0f8inYe284bLPQLV+GY3jN
MEXeDownfQ1XMkRmpoKQffYgJu7mFcI2ZKOseywe611mLH1wXbfbRF4Rvc1JdusACIksUjjJVQ6u
D81bYhcsuERI65/XAHDTw/f0FaLZz8yPZs/ISojZ+EyiVPip3SyoXkdH0MlQqoWfG6g6CAbk7fHt
RAs1/0TmZ6RRHMohe9F9KMfJ8fuR+uzzPZbPWMpQTUdbs0tlfDuihKxaV2BwlkbFqiy8b/ixfIay
+CplNKaTo+hKR8G/HWXBZOmhsP3gSNhTQWZenBPys3Agjhs1LMZDRXD/fw3WU29agKKawsyQMIfB
uwdJAfELyr9Vn2B/Gj8amIrnv7/EwG87MQdATVlKpaT2rC7q2/QeqaY6t2g5ZcxHrz6jaqFV7L3h
rJ2h8jHm/bZ0aqatN9gOw8qs4yHbmsflUgJ61YYqgALbn4mqODhJOYS65WqHi4DTLpLz199Mpc3z
3K524zLps1h8jvwiCP7RXJn+BrDwCd7pn7FudWSphApdX7xwLT4A/TdEXehYAkeyaHCEyQaHCzKU
uFRtvb5byGhLgddPAPqfkxp0W1XXg2tSvl0KsXB4LGz1Ntg1VEZf7OMzmfnfkx3VtY9VvgmOrOLy
ZDlyRwQXcc51/QxMGyQMRnrH1m8HgkSM2WcG/LjIsAHx4LJQx7ntDhpaTI77MAnwRTfuneyBp0yI
yPCBontI6UWpyjiLIQFMdB4ObzcP5Z4VrWCL65280gn1QslWdDQMQ/dLsXzJ1+39J+gCLp4zK+fp
ACsWezJ914Of6n/eX7GtdzBAh16Wg4TUV0NHvvV/K4OlYIHah0uTwKoiYlDMSTGOlQvIm9NzbYKI
aQJj0WtlsL2y6ThcYiDwSAxYXaPPVlZP1Gs2bcG5GwlxOL8c3INKRK7GfF1pVISY4mT6M6Z7we07
KK3v21I95izwctIw9TrE6+//LJz45mD/YU+gQvwa9EQ21OLhQ/y6A/zBTkEsG1d+nQcjV/6nnaiW
35PndDIM1oqS/FRY6W/cSNmV3SnkCjtWHwvwBoL/k2sNq5ACCKsTKwJFWnE0hPNfC/kytLOu7R7y
Aha0lwXn5ArAzZUc9+NpJAinPLIBNGR9fuqB1qFpv2484l9jKgRIadsLsP6z/NXzupbjFRTQkiAb
NPogcioNU+TDDqSaOVytH2G7T9jMOBStGtJFjNBX41Y5dHAc2pFdVBk/9ai332N7xeYXnSLvwiMX
Q7eThNG0530F+1RZgcQ9a0nEQk3EaVOel8gNteoAV/49OvoXds61NXCbs+H8un9odrn2y51CBOck
ZHDik+Mr2A/+f/lOyYDiI/Ldat+fmlHGunhctk7UWn8JlOQaDNIUKr+cVNgddn/NAT4l0QejYvPL
abpNVHmXE7RowZdNqeo/g2Tn6PHoCcnF3SGyqU/i+RqBQJ06SjHfjvyJvism3mdRmBQjudvKJSwK
8pW1QLtkuOsxPu8kimutOP7Uy6AWLV/9aXaaVBNoJylCpB6UxVQBQuF91+DWESBt3jEWYm/Z2HKj
HmkAsZj/eHBEVKOGyaE5jhi2e1Ehl/SYRKR0570Nr6SpqD5Yw1LQDnSL0WdHnPbtJwA2Y53dR/eR
t54+1TIcVtkcbSheANdf594+niONnw4HIO19Tibtoz92D++KXHXwxfWC/7xGZxAWO4cHimtbvPpQ
+TZGve7o5qEiin/NoatuHrUsjNWLoeI+pk64n73fJjLqtOpeASAcPw97UNTYC/nSMZFbjSoH62Bz
XZ/8h48DcMFS0MdZW9FQ9br413fAfLzWccMCooCBs6ZPUJebbCSlVK3c8aCPxEiM9MhJsixUjVgS
0XMdzwV9JiNsANZ6dngeTZc52BuOatDvfOaQbTWoUpKNIciXRvqxguC0D5RXt0GeQmVaCaD6/wHr
QVEvQbkpQw9bihrHRFFjERS0XQlAgdWstMey0WnaDuhTNEaXClRl8Lx5+z+dkuVK+3VojFEEQfVv
1obGXs2uY0BpkeSDCagm3fKsNCocOekXFINZEHhGmz5MSt0vQa8Ky/oVxne7CLi1K9q5BTHZRP62
kIFXzdnIaP3DTxsK1VemeWVnk/bCijwBA9sDoBQdoHdKrHo+7uod50NxfENjo/ZCIwWvcXMUjCH/
ntqW5oVX5vf9UQ==
`protect end_protected

