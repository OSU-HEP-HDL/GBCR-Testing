

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p7OtZBpltt/h9CD5IsJBmAQ+bQJxazkQVbRBjNJ7LWO+cgudo/XA7alKhPL+qAE8nYmt8n/nhFV7
1FHJnU9EmQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o0V8lbvMs2u7Pr48iEK+soyjigqgrrzx5HsGK4k7Ph8gI81XWNRtIljFPpaeGwucYu/H+gPVGgh4
LxNZUBJhgeC8kZr5P0UJ497gR4WHGLQSo0hvtVYHYDlrxnVk2S/+il/2gMAwvI5YF/lKiRUCJMb0
2mL6cpx+2git922rE9I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hIqrLT0Q92Qul/GeORaSvJHHAIqLk6EmPwtSD3Sw8K7TFMN/pzvjFhA6g78oxGwtYju17YRUOAPP
BxWjMZac0YPGSx1A1AySaj/jWf8/sND51mJS4hxixMPKgd+iJln4gROFDpToYNAZ0eBhqGsKoRPf
Exo4YtwLGOksTW6jkb5XyScrMy9eg1uc2W3HXgQfQg9hr9gpWWe4xqhKUCFXFb9eiIDe3eaUQ22t
Qgz9S0YooH+uhgkKhXgOsKoG8s8RO9q+oyyLd0ANkoAdDySOy1H2+qKDhuJHoo8oHgkWp+t8x1nO
sbVK5ZibMfLbKeRbGwFkFsj+EKfWfOy4ck2AmA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O+omGGx7WVLIBeJijOGvFCJZ1IO2vxCm1x3fAW3H6+gw883MkRTmRZO0ddVzk3pvzQaBPeJUDRsY
1XbF7OM1C/khYSkVv9TjyhihrgNNT2rgkTkWtfQNoOMnsmtYkK2fHBBMyNXzHPZRBh+2VgTZHxjv
olfJ+wvlLAdf8BqZKWo1gutmRCut9sBqwVpKtMbEKFGRBnt2pETIJcWkewW45hEmUxoPlXpgWrRg
sESpeoKuutTTWJor2paEV2RoktNIWs/+x82raY47L1AIZ3uy3vEVemolA7/fyBhQXHdXuWEXntN5
bzesBXIrWmoZpCMSf+IISz8dywoKgC/dpdCKGQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pc9IPtPXrLLm2VmqSrmdhsB2/sqloTepqxhS9rXzXINDRuCWOADiBYd/5aw6fJ/PtHP6hvfQmgPM
pe5Rbb9vXhfZlTdZe6IYAV6ajOneMnpE0SRKlyLpgkbpQbwWF8Ta9x699vjybNfWF62AYBS3D7DQ
b0t7dD7uNK3C2oBkpBFbB3y/rTrUlQxN4AZtlp8BUDmTdKIOwvLfH64R9omltAgRoa9eT5fKR+NB
hJulrR0XnMdnz4MTDv9F/TNStcRrNIf5MM0b3o9Lm2heOPvkpoBOr22fj5c2jTQHuYFT3gyiU8GP
rFykj34Hi9/EcnhfJs9E3mtp1Tszf4e89AyXHw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rp2qWT1ngiwszVInFfAgNDsqirvFBRH0fhGMVLdTcJjuZF6cagj0r5deSp/lHSGQXbQ6hn2NE/pT
sVS4xwCY2B03TkdpZqI4G+dZXB8686b5iwRUQ7S4WwcHb3WXRb4Df1OHJ6dgH8h0dIOxvwXXNlqh
PKzd3cQ77q4ZzFc8bvI=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JmHrUUSZT8PLNYfmwBtqUH6qJ1p97BdaA2q40RVMw79ZG2/5JMAd6P3xNNzdIISzZU+jzu0NYPxL
Z/zfPbolJrCwAck6UGljZ/OOpPHLUDGkBAu8BIP536kFNfmsl2/w8PHTByudSnwDI/YKiNqfsxGP
M6Sq3+TkXml3dJEoLhHWDNi1mL1f4wADZ5vEh09j4ryxXNWZ0T1vCwLDq6JQfC0fF5S+fWguWeoy
y4GDwuB3WNo6v4nkxnIBm5jk34GhklMVorbQQ90znGRfAejdTRlBiH1jH/CASbqnXiNzj4+1wJ6K
83Kv1+Hi6TU2vQtu3O5wYTXjTMpJrASuG6iNvA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
5QigutWVzZ75WW1fsVEiUpdGotpSyssVZGh3VadKZVAb402OiwpapaNL618YyNlQA0ygjr30ANCN
FQ0PX7qx6tw5js4RumxEochXs7ajtqKH/HYoJiKdprO+EwGDUyB6cIfcaJm2QMgrt6L95B2bJrOz
+PYP0YPWNv3NTCQ0EPxON7ujYs/6mioWbCUESojvGfORc18eXxTuFxvpyrDRB0m92lHVnQnLdDm0
T7Xvfp2xhjrtkrJWN3HYz9crVDl6QyBHhhrYlHiTmRMctmP91y4Zvrw59eTKkfSo4IC1BfKrBp3k
S951CNhOf/XU9KAbdPGDcr4bQALYnw1421jw4BpdXegXFBfMSVD1v8xlmsWyKb5EU4KI4NiWeEtr
L0cie1OMo8dCWvOLlxxB/l3USS28KtM0UGLoBS1XF6foqTnpliF2sBiduCZAWrN04o8bWvYm+x6f
0G81F1DrAxJ44P2rGLvcLpMFXaE/8ryIFSUsTHxGkjVf7wWB5ghsPHbeHdLUEOTBLSQ+O8JUhRFo
xOxKdcSALYoR+zxQSTk7chYvK0/BYyg6gvJzLv1gEfikdnXQ/2Oz6uSky3p+4G0Uv9cFejZV3naz
KwH+1pU2zDoecgeYwDeQ20yTorvD9gkWPGLHP81JRG6L45xCP8Gaf/RLz7huzRtKYLyq0xlvwcJW
2EbCEFArHMzKk1JLHHIsFUCNb2HPKOv/eVYJOkENXvFgc4bLDYh6fX57QybYon7oOfyeNJ3LNWSI
17ftGIUXm79qPZWdrfSpn/RooiRgVlkjOhWNS2Q8LbhWT8mS3bmlgBt62olI24r+3Xudgy8PRkCA
RjV2jqiSheU1HiwQNUsOJY2+1Xrdw/6xJagDdH+Lb5FRuoyI+MuQKQVsoRTb53d4Y+ZR1Hy0jpsP
iZzeU+zmkT01IusQiPfCX5Hj0zt6KfQg2N6IGMIA1Gm5ztv5c1eMC/zQP99O/NPa6qxXSgIQkYEo
Nm0FZxEAEp+zSnr9/FHfuNULEkHXQJ2aL1+2qhumMDv3V8DVMP8cbeb6FVxqLarDbAOsCtqhcJuA
JesaS2MvSExbecb33x9ILMPeuVMRa249rJKVkaXG8E95xbDvkknpWFdp+Pi1kjEZetPEPYVqyUE9
TDR66vwvvgZxLptit5kwr++X1NE2rz1MMhYR0U67ObzAqn9jzJ/4pzQ7XdI3BKIJ/Kk3h9z7kwhO
AYAGIRctTslQxqyvhCJkAKlhJ6wUfVAM0Bw2LkmI23/Sd+mxXw0EM/36j0gxqlDXilSyo1XRhv/Q
Vso9Nfn1A72diON+XX9c2LhKXurdeHTO1+BfqdyCKSJnDpr03KWHW1M0jecoqyR2niw4MNULRqhF
WMN/ZXE+1Qs/k2B6DJ0HbZvN9u2Lpx4PGVpZZoI3ZOoKohvNpyrqZ/0L580KoK9KoZOHrWxQ1ope
6iUrmP5Xm2PDpB6w6v13d9RmMTrBB9VcZCxJmwANsEDhKlv4QDj8mscrgrQG0j7kX1n7Xe1VQ3A+
hhowPE/WwDeGUvSX6Q9VCsJOZkRitazS3c2+hZuUppUA3NcXzsb7jcsdzzb48FcasgXuUuW41BgZ
7EHTsWafiuzOVSGfawSmrkWZ+S60NRO8jZ68XLi7s1xcYX9YEq2ECMA2UK6LzsjUqtB4yoql7zwI
g3w4p/l3a53Dduu+dOkhiQDxQsFCNlzFANP64YdLPDGGMoWr54B8nqykxmjMVIS5p6zC9/8pQILn
76TtcoN7AzO9xzph5e5vyBnBaUAyxH7v578LF0dpyoyeac1G5QNtn1egBB2Tp2mbEt89VSl8RvJ+
/YiHvw/Vf2/9Ro4l+9zkq+dWuWBr15wFbzFV2HvRQqKkYDQCR6fdwpHYY/bxO5/bj0WZCt5N15Z7
Pqir/y4+/zmxTCnt5LJRDvEXOhKTFWmG5owzojturaS54dIRLKnOUNVteeOFZeRqpbAF9Hn8unPQ
bcKBBnpapT026i/jJ5VpEu5NNna56qin779CgzH8MqZ9kM8X8QSn1dxKV3xZUBSH8awzwu7uvoZE
tN98jmjCf9jhAAt5MRZxtpuOfL2Ne64zW2f+VbWFaAtBaWgZtPBxSuK3AnpYcWl4F53bKewGg9Z3
0bWwMMZqteIvx1/gn6Z+3elxNUGsUhHV4VVfCc/FADqWwnjXdYrNPoPRjrw1tFAJHHtG2by0en8G
KDmIX0x8fonFgtmn/sn9OTZS5XAQ2KWEk/bwwW1ZJzjcfCTekKqEd3WqBZWL0BKEmdgDv6Wv4QK7
xL3uVgsz6+Wh249PhVSdtXLK97x4BAmNI8Wwj91ATSfxmX3HdD3zlK/jXlKXJ/4n7fAbXKdlqbdk
qYlu0Ja0EOgaj/RWMOvl3WZGA836VDm/WqRKXCByjo7kZAbeJuZ7tHosRrzRIJCAKAW1EUEfAoIC
p9AA2wtCh+/meJWHnDKuD19JXum4Xk7/bnSRHYveKhSFFS3QlYfL3JRl36R+JfS2Y6mzZ3ZdaFre
zmzQeXRXJB9wnWHtNGBYrAsZlbZqhz3zGxHoUWy0PaJtq78GrV2FROpHTqjIwPz/R5Dt7if3XBim
uz2fq40e5cnXQ4fmmbHVPbfm0tui6UWCfN/isThxOKxldI3rx9yFVgZpA2yZpLElTxNHpfXWGgnU
VFPV3A84LKZEKw1vFFQuftDs68u9RP6Q/2Kj4sC8KWPvFnkORXBp0Ei+4Kl7B1rQ5pDKXuf5d6KI
P5AXtgdSWka9741pw96PbV8p5y5Ok94XO2Vhyx2XKxBsxcP0X6rUILJOLYv/RulN4o9baojeF2A4
el9R3Dg+z+3W3ri8ma53aVC+K0WM1sYo4dSL2UBZLz6vTSR+39mMz9fw6bxMW4BifNFpXRkFehx0
okjLazsadLmcYdCu/lNmTk5HwWxbckbYITC3G84+AHBOBuYiEBOxckzLqEi9r1lUS49DlKr08Rlk
7vUnA6+RGuOwX4RVoElbT4QWCjG+FZ6B+m8gUW5aTv+ADcu7VV42KuyLSdwkg+H9PZMmcJ08s0gr
xlThMFyO+R/IMvo5MoFP3LawkHkHEUgIGnP4QBjbT6JkKSSP2X+xjzntIAL6wViD2WhrA44oar29
wAcLy0zjltJ5G/Yi+EMTWPKXyx4P6v7UvKHrw+etUAscpUogX2UA5yE0AeTMjwmRm9VMaw+9ENFX
o8IErg78kBtq60aGeR+v4thOYa+O7IKZpGFXzNlaXLivERYe7QjhfK65dRErqQspkkscmf/b+gYZ
fPzXNrrCC2ExfnS47u2CQ0ll5zfcRJu0gjY3wUwGTfcy7NhBGgyfYOwFHJ2eF6GlLbd32+aYaiGK
lYi6t8H5sqGaGe5Lp95bsoYGi4F/Yi1+zAKuBfRXUKt/Meyf/Ev2x6VkfdrWqYJYKJ5tmoRKaqaw
wrKDhCtrB6hGepWpL90Bq3PjfsZUMeuCAvhiblgnxBZ5014def4ucJzE1SIZNrij88TCgFfwk7lE
oi++ACG7CcgZV/A6+Gf0X2NFwerQzkdXRD0V3QZdQiUKRnrmdxLx1LAQERFsLfte/lZI0Kt5Rp6Y
69EglcMdapfmBXX5HflspzLqj54605aBqqrbstCGzGGlIc8cnx8g7rqRohrpGo34gRFJjbUgY/AH
pPOqQCRd4OLOufk1LN19jM+mGWxuG0OD+fpKPvF+ITJzq51MdGRbtR5DxBJt4mCJu4Y/e0rwAYw7
pCjX/W1pR7v692ZCqT8Q6Ar6IEAxk84TpGeAEeH8rwcTK2Qc2+ImkRMDoYAaqKjCJN+ddIJks8S1
oAgN7aztaOkSUIgtmMe2QVRqC/YybSZnERY+VE9ui8620WrmM7E6+Of1sHoL8ydBAsfXlZwi4IgH
56xV4dIvnTmqYWw3ZZ7slISrCn1Eqz50obvUET9XKHvZTnvpGY+gfuACT1ekIgWkOWSsmkcNndku
AakFtMUakHFPN/l30UP5tuWH0secOJXsiemI1cVlOpMC5CXohMlU7RatGWYMutwxo1TayGosss/j
REv77+KOr/Ibd4H5n4PqYwAcJPUOG3SOUCumyRFmuKXuU3zyr4ABOH4LIHhiRZhKOO04NzRhjNvf
Ibp/GNi9d+aPxL958juL0b9Rq6l51ImlVjPjeauHQ4lYIh1nJXYGQ2wY9Pdn+NNPTMSvbcP5j6Yn
1tHtUwk5ebzfqqasJE4KbC7oOT0rOCBzT58CTX7XjBsLCQbTEmg81Qxe6sb5FXEjUqCe1ItbruQM
IhX09G5rSLh32QImvQ2i65zp5plWcHLujY9IKqPTwRDnRs4fCxMyxGL0CMSxmDuimQ8E1MkaiuBp
i7OrF+STM5qT/3YHgaMdjXrLMRBwk55/LuMOHRukFZBL86qXlaZ1+ELtkat2a5z6NTttaMzqXZD0
mvKmEdEexeTRjJtqh9j/2gYCxgD+8gFXiOqsK9hG+hGR3vanSP97d0RIeK7Nzj7w4W7LNCR6022g
gdDO427ccn+Vc3OACq+tZIW2foIhgsFeFp8qo6KF2yMjDbfqAux6mvx7NAcHM6d2U9it5XwAZaVg
5uXiufU5yRLQiasv1NLtVb9wsbR7Vb1jwZmaOsf6xJr0BIoMaiD7l1VA6TC+q6M/XFedlVP0KAMH
Y58cVgoYM11vG2Cltng7SttnyR6qsUfHQIIIlFZJLfUn8D7ErlNgHSVVPDB8Trdo3K7h6xy4Sz5n
92WFMlCPEcbs2L7/Bt4FIAXyFwZ7r6efY1fIKoivqKHQCtvstEI1sLv6rpkRPQPVeH4D1/WHUvwc
enWPhbqDw2TwqBjFlzFVhaTZ88z4T8ntgzmpjoFYOanMGNt58XVdXJtqx30YpalYiYq4+5kZhplm
7K53PjgKuizYy0g52hf5v0jDyWSLPhnhEwW4fI/oiUAqp6XHcW1dBD2j2y0msKf1lPk7nW/5HWoQ
0+omniwPMVyvHd6CaN9qpusRLMsYEj48wfMhcDFP2/zjgWPM+JTxzRwSqrE+k/eMLYwASdpvdxcB
9mGWA6y1PynIxJ38r8aON7/aCqtHMMsDZSI1qGAueXifJRQ0yIFWjKu+5Hy9ZoPswb6Ez6/kBRAC
fY4/kUZNG/QK5l2CB3AZQl/pCCb94JkV+e996dgw/+CjgpsDzPCthkFs9J1zZJ5m2EpVQkf4+5Sx
E4/vNx5co9Oj1wbRP9ivYj/ZDj0fUrVe3zd8OShKjghBgOpqYaxhrrApgCkDGZkUt2MMFY2B2ERl
KDc0Je6MwcF0vu9QXA6rI8tt2wwD49CMdDCN6Ot4yXyQdJXeV8NWPZSYBVONVlXQb00JZrt5mM5G
e0bKCQSP4yccuo1GYJmYiw+XEJAnLAVYOZyH4k4hzxp5fptcV2PD4UNE87QfW2Zppx8KqFjbjDvx
ELz4Sc/NlPlJz7VAjiZzCFicGxhDIu3U3AhEVf5eAUgGAb2WWp/ThF3/49zye9T0DTkYiR3nYxIh
c5d/BFcbUn2e+erq3Mv0V4narIeYYU745/TwmaJXUIEiXHmqWYnIK4rQ4Z4EfInNsrThg4y28c9U
f+KgGFJtTWeugbVpECcfYYPrmG4MRs9Yem8rSGd01C6B6pY/aga2Qyge0M+WJmssnAf88g81Fyfu
8nOgCLgFdCigTjc5Cz0qv9sGOWtxVG0lyX9oR5mlBLlQ9IDBlTiHVFBUgRcJcjGXdfd99OZ+4RuQ
6E6BxlTbin3CuTtFQOzHxeIoa6BSNdO2VbQ/5M9D59Awtxo096JrMcyD8dDbuzYQDnNMpy+3qXRQ
71lxY/95/qU1JGBpYyQc8yTsuWMaWwx47GvhupYGXxIIfOhNo99bfrkNkfM2wnKSUcnGRCIi8aju
+IPpwKyAFU4pSlR4dIQOJZytlNClNwF8qlPxebetkgHPHu3e/vWsn3qGKvp8XhfbBB9EzTwtUR00
FOdsNjeJXtWE1B+SXqxSksNEDSjCQFXNUKT1EXNldicQkIHtfwC0x0JF3XBOKYHkZA0VuOVl3rXl
JEA2A+Wks5tEQII3TzE030Vza3tzrUwaN8kzIkxA5FVnCQzW//WHSJPH4JUwLdtnHy99hsZz2gZQ
hg2W1oOUP+xm6oGqX5PQqMHx9tFV0BCS1Lx2WKuHk829HLsbqJSlWd2qkyHtuvM7bKudyDyxqFbP
UYC4DftYzkiQ0RJFtS/kVPI5fSudBKJijK9evDCneu5GMwNn0x0R+YPrmzivIUZi6U4iZGpj6tuW
U8bfA005lSX9+aMFLffancaJJULR7syM5gK9GqG1a/c7wmv86B545xZWvRf55iVzx+2sXo5wfuN7
XUWNy6SOwqLG+hsy9f2FZJdj53t3qMNZlTVtb+7F+C5JV6x4eCs978oTOTDiUzCbu06oglfYGH5o
GD6MzXHLk3C6LQFy/lHLAtIBX71/4JUg+3/t30ZoxCDOf+ItpaIiwvjdWXUSdyf5K8f5oiHBu2+o
JIOMJSv8P3u7k9ZMSsu7K/8pUh+khmZlXMji7AlWNreCu0hpwkR4sLHaDznGQc4mhr07oK0+UZeT
g/fcVxG6FQvF4MFYsjijq4yppOaoaYcxGSIG2o+v/z/q5Ty2d1+3MigRaIaZQ2a1aRiqUHE/hzGg
ToE91sEx99HuETIzI0FcRy4EY2mAH5luftPqyoDamKP2EUfsYlVhmvCebMqsoBgHUbGOJISEWV88
6q2WDV9I3IZ6EEwH8OgUVn66DlOmXWg3aRVgQBwKdbxWEKAGfLJE4R5X+1ukPNeYwEUQWPO86hIr
bLfGyjsB/n0Ofyz+4KpR/f7ZrpI39lszU3qwLbm4doRvTCLAP2WWxFPc03pYUs+ILxHM+HutOpYP
nGeVOBVIoWJTTblCZbJGzm8BfgPwMujU0Y3SBcfync/YTiG+8JIY6tZ5m0z/vGM9mlZnUVp70wtc
jJ1v/fcZRGsSSFAfzA1BquZZc6jAYsjs9bAYg37qokle2xbm8QPsXhjxywOwvHdJPlGh8gZ27/uV
powLe+hn+PtoyL6QSxwpKpSK7cNF3gwlxBSDWFhlZ4qnNmdhNPvyDqr7ZV9ulIwEDdNbNWxCS9+Y
/sCiL47GSlpQYmn+MshSFcYDytY1TyHP9Sisl8tqaXAK3jU+Lv/QjrmqhWGTLp0woyRk9wXAbAs0
zrBVIdLPmT2/cAcgzQf0In2gqNacTKsB8M9AKRNhtj1qDBaVV9XWKFCecC0cgdSp7jgNjSaAHr/F
Z0yCqskZTDMWNv1bS9lnrizEyz0G6AjeEYFRYddF3URKd2bvLKXmbVtO6qTNJu4dM9NTqKGrDg8o
3ZjcbJtAGBJrPjjWax7aYqNZ+cdMIHl6sl2pwaXiS/cj+IxDyr8nXDEZfkCrguNdxXbtueH7SgrX
RQ/ul25nn5zwd4404n8UiZsUAqy43FzAS2R7C858o+tT0FhVEIFdgxmtOYJO69mddfpP8DtkIceK
mlewdB5p9tSnpH487ihju/OVvBMLGWvcbWBQw0EOyN/gSlzw5zSoR5WzGVqIUlG/1nkKJH4CTrNh
8yQc3XxdAQPLXhcBxKpzBTWktNl+WCwAhhYLW3pgctgYAMMxNx8Y/Ahw+fsva+fB7xLpeBY5/Jff
U2W2JT+aTGlWGCEkKCLhXJb9xf7bntEVlsRGM2tcoBdwTXPsVhBGc7lYp5SCcQKvB8+bzniLymsi
3hHKXBfZGzPyMoH8fPcJmaL6A4yCHs4jl2S5T1y758SdtEnPKkHgsSI/ifOnoWlDdjwFhadBMxFc
MHicg4JxUS0wMRikFkZvki+gct7KhLk4qct0bW8OOqu6lLaW7lNGchZy6pZDnv4kLq/OVlxgvIU3
vtNTXsNa/ta/5Ggws/K4HTgIt9A/c95Ndg7AudxvwZu1SV3jV6upM64VcwMXLmOYVdE880ibRWzD
FkCbsP3y03anJcPJTpL1Izx+4F9ywe33JITni9Q7cWjHU+Xs2r6yPd4+Nx1J76R6U5O6fOEz3X6g
FTeZbD1UDIBotsTrRwYMZorHEbV8qE/TboSVZZlOlUJq4cblubARwYHsHh6uxinzYVHgCKPZ3Tb1
qtj4YZi+bT9S8qGwSTFvRrLRZZ+dIIWtZqiqUrNW6dL4p7rkKE3bWQKMoWDtNNtDB65mlC1IqFSv
bQKQFQStAuuYfY36y70V6AssnfvrEKctdEO9m9/tFNKg0zTl+4HV7Iu8wq8MnQvTj9eCIZuMpwJc
85TJEIoqU6LfwEsuKPhe2+Gxj/4tY0QXGZ9oPKT+tVpQnR1iF1QPN4gA6QvdpAfUk+C103CL1Dfg
oHu8GdtEE2xEtzKeAikfYyzAlef6I1L8UVmGGpJ22t5dmEBddpulelVyQNP2GyLT7O+apaXxjk2+
pSHGYz355omkky3lZlaQ3XNRPfyPW3X8qNedOskIltZfMLw3D07iiLvlsCH9cp5A/ln1qjDTIAT1
dAGKiW3LgxLYLQ5WoXfR7itfbcfZkYl6eWdeinQqwxk/Jtds/fLn8VWb5RMhS6rICBwc1OGUp5aq
vart/lSs0vR8FB3PKe5scGTJeaYtuJchmpWU+3KxxRPexxeSUK3in5i4Yf6JusrRnJz+X72btbcX
k2SH5GMm1zm24ajboqQMKZIC4w05Kzj/lkGedNGglK2PaHp00zTNadv7Mxo0+2oOMCrJhueSei8K
saYeIH2WzxMMcBLZCU9pK1v3leweC042fiIKgkpvR5Ed8XnltoqfvN5IrhENsBvmbJCIOZwdyOO+
hS6Yi7x1Q6+ZI0W1sby5GgtAFXHTViZESw7PnSX/TJI6xbPJfYcDOtXWT/U3g0w3/Wfj2ifC/NNu
Aab52d4dcrU7QutuLll+i/rqyekQemukYmKCclw9YwQO8JTS2sEy4qrSzbclH+pw4xepsNhrv2d2
rL4YBTgz8psgF8+9yFYVPiDLxzj2smzb/ICVTEw/RNtYm/28NkqMXO5HSSMfRbkgrQ7xuyl7w/7l
0FYpeT1QYEcTpruwngotAZZjXN6tUahG9EAOmgx/Y6WEfTLzOc3iski31hdCaD2GaoBT502P0O2S
u82ccolDKB8DidFY7oLZVWHCOw6MLFWfFW/9y72/A2q5GhuvtvadSxKyfuyGepywu/iFtivkuPz4
PxbC6rbsiBhcPoB+DhMn6Zi84hgUHCrwUkoPLX1aiPyYZzFmTOzDCvSdlnIClt4t7I3d7ACU9xPB
W8Cq5vBLo90zXwlRROU9opyXVPrb1epG8KnJpuvoZT44NCV6HxtzIKjKW8hQJl4HiGoq4DijdHL+
OEegQcaUgpEUsq6/QWrdcRL8d7rBUJI0qYtQdU/nnR0SCwCnxNova9Ys34+zHRPfgOdwh7U6Aq4F
f/3zA61+7hpbGyT9OPJfajZNRdeTi4I8zj7jRTQaUMZcGeXYlIl6JP0vSt2mLl+pEU8ZwZcV+mhw
RMJM8EVtYCB08HO0vrn7lzbX+YwtnQDEYujNmL0naL1pCH9z3i8e46tsM+ZT4ML5KxSBKsHW+59R
hdz5AV0z49YFbx+f6pCOTTHjABvlH3x4H1WlFjJR48b64zZPbml4HKwc0mUGXdNLNXUavTo7aS/4
5ZhqtH7H19jNoBmKDHJ4gjGE/M5E3hZ4PxleIr+qnEF3bZpJTf8LsVqjnEF2nEdzlveef/igK/TI
AS+JJzcdU+pcPhpOAga8iCEhwt7OSaYPwuYnjdxMh9Nw3+uMyRN7aGarcIab5hCxxiXwgJ+ESiFN
6pdHLSF1MpSCgkJbnn3vsauBShMCmTqrtaI6Px2glJkEnNUb15YHgr8pOtv6zbgqtNlQSh6bsS3i
M66wDVTsZKKcrFnfhom9OlFWRgwtDMViFL1RHZOiYN8ZIr2P/FY6knzbD9EAF1zdpRfTosgPvhW6
g2Q5mlxZczo5rrIBA71P1X/0WmNL6F/eaIyxbU/CpY/ugoiqodXnGjOehOJHhJs86jOU2ZIRhS8G
lzGcEB6aVOLjKGHBlpGPJ2fjY9O74SRCp3kYTNrwoDcWRfSmi3fbLv1YBHqXgao440QwsWaQasDw
Jes9C7t1P4lueMp21vvIkyTJxEfws9fh+daisE4X0u1Ti5+kKZSqZere8jWd2zvEfzIxIux8/0LR
RsAeClijbgb6/oTi/KHlDLFAx+GZPJB/xtBXtEGmpjlabrisquP11IsrWT/N+qO+Mo//0bcvSQes
yU8k02xCNtJoz+rwJPjeMoIZhTE2LOHKgD0xMK/lFdBF813vFGisNebwomQ7am43SFyLhXoj+uy2
Q9hxI2H7ToiLvgvUIAJxUj6ZDVqbIZgQPJRryoe9bnnEpf8F65103zAGKtj2cG0pa7ESccVDNkyC
KudnmqMdvXIlA2JCF26VUm4feB6foZAGDd4TO3TqL82ZY+k57w+MovoKaipIFhSqaJkHoXh6UrPQ
rR1hFGDiM/l2C+yOoNe0yjijL7ITHDSvx00RC9uewIvP7NHJbwIakJMH64MW245doJg5X/fL5YQf
w+5n3SLJqLD16eiKnhAN+DJUo2HNkL5Iz5t0N4VAp0ueL5vlGwXRukmtmBWCfqZzHHRrYhMtuMjU
usVufDlwAsQZgxiNq8DUB1Kxsqot7bSDoG5x00P2EtCZVnmWEQDIyG5HoiuRv0Em4eYW+a/TX6OQ
T837SPWYwUvaGL83nTLxlhzGxAMzNQvNMI4uSfxQXMBfO/LSCefElyF9lZGbqHgiA9ijKw543/3w
etzUurO18ekVf1fTekVYk7FnmOD6ICECv0Iphe+wwp38xpIPJtNOBZsIxL2d0D9vyigOMxY/Nj7H
qxWZ8rjN2ABbrJjmORlY15k/fVRH7dCBnZhc0uAIJqPoeMyMyrdKrD65Kt6iJ7D2jIkpSdwq1zMA
Qrsv+8Zv+hYHjDQEHbpW3mEjhPldSxBkGwgyPrj0GJpn3wC3uumbeGg4RLMeUI/drIZBnruAengZ
YFsCoI5Yv+jb776OMsk+4ZMH3yCAnmRdDaHtcgRPrtskSaSb/r8guQVfTEZ2K97VAj3SiKkPAncd
dHeItu0SHEcO+gBgA30GVnwK4+p1o/dz5yzfzXbCONNsAXl3MGEunC5GaVQ0MX8pF9wgu92KjvVB
FgMYMNtEnQpC0b+BL9nznCTluQqQuGcMF7pLdlqyrEgnFVK0DZYpvbwW13eX24lpZqxnsAlyPVq1
VwINJk4CJued/rZcpTFqEHUf6Or4A+YiOjhp5Yudf8yaez+iYYlCoFq1oeMkZlfGxhdlRI+2oB22
NJoS/gtTIfBAjHxBX8sFgtgBxkbdQPjHH5+c+MYr0GhC+Wz7pJAdZZ/R0chEyzA/Hyc81ZrRxmTK
Au65agLOFcY/Qrh3w/cFG3flbkZA1lsYLiY8sfModoBRVxgG0f8TzVyYb7DMvhXGfhwvuMYa6zZU
uLnoXAtpsxGxexs/zj/04SRsi50ZV9hXNzDs1dwPwpqCaIRD+X0xynpm7U7dk/oyN+lIk57fUXZ/
2jmVpFv3M2d/v82C4TtpC1AXV93snvwJfiPOT2w+KIRa3XRMcWNvg3kNLuBkFzo7+zMkzEqeJSch
POrZ+OvXD1hXJBXRXInZvWlytqkCc5IPG6Dhj2VNHIuNCY0d9T7F7lB98VVAlteiE5+Ej0H3ivWj
UTX56WaBqw8h2+KsmWLG3SW4lRttAJuN6q34bDtpvT8BjqJu+rPhzs3L7vq+6KswotU6fcgu2dl/
esgQy6jh9yCjj0n/ISty5vo8OuFa+dvj6/19jDx8/BnF3jCEOSbMew03Qf4gwS2juylLVDdiS7oG
TuSHdAK9cR5KuplSEpEPIPdjrpR4dh2P0m7ARwZbxl27QwOdfnm/PzqJfXjoplQ4fCr/i6gFm1+5
AGiaF8GuhmP0eLinrtUFQh29Z5kp0oJBCRmWgxsCk/XRkwR4pbMpCqwsgGR68TxS8GVgerM02O0C
ZJBanQIbFO5BUmj/0pOO2Z3SWwCg6ND/b7KtROZQEOUItoAfxU3dqT8qwMTpPGDVSi6ynHjDPl+e
H76h9LLgWmBC+1hCLlX86lYv5KpIIyglayJco0MIYlerNzMbp4J15NBqY9eOTNPuJfbrIEM6R9lE
pIrdVm2kw4HLDxe9XEujqCgCeT0dutkQSttf1AHZ9Mox3MLcLulZ05swM/LgMZNUFSvH1n3yTkoY
TP049XA9D9WkIwbQSvG2ShPyuCwFRf73Y8VMrNR/HIKWsLmlpdP+ow7afmGgUvtfx4Emjoxvz5jC
hHyFO8d26t/0g434JZRCewH46gzuXQJOIFduDtYugNie24Ds3HYR1U13XJQlWt4Nua6c/tyUWpwB
31ZJldiTfnOYsB9GZbMlLRiGTbvCBY1tC5uZIMJhZKR4b+e0OJwsolzygfkQKee6/QAKVZhsh3fp
oBhsc1eHm+yYvMOmoBj6/wc1WEaofZY7LVmocuavWzvOy6Zikkss8tGuI/WY61zeyB7SRsJ+0Qxi
ljQ/CcG7G71bGrmtgmrqKV7OifZZZGengnJTknDgRqwNl0pqeHv1O2H03N3WOOh0eV7v6cKEtZRo
4tJdUDjqPJbgLezA1JILmHWs16XbAHzwQwGmLEQ/QzY83m8Z/jRharvVFXYZpQcdjVGY2WW5Y9rp
pjVSUx0+KCOLNw16kQF0YY7EcIAqo/HQ2nxSii2jm4W6tTl5liHxwq/1eYXkT5+yapfuC1m8ET6N
zmk66QSzhppxPLrh/NgBq8cbg8e6UaMOu4jbnfVnlsXdpzuBuVyuJXwKqAq8DX/AsIn6z6ldIhpJ
wh1HkW1QyKraPADtHI71bauSwpoBRPunaP/9JWMQ+qiKHT2xYriwmLL1pLewyxBHkfQxgmeu1KJx
BPQo9YFk4cF33V+tV9V3EM0E+fUk0z3rXzCrXGfz9kTMyA5tQeeYYLu4e0KkQP6DqWhDx84/ETid
TS1LEQTjif3abzI4jhMdYQO37mhtbQZSkGXVsgfzru8zudXqWaW8GrzdsF4YGODHisNabRK8xyp8
xlmzfGcXZCIW+uA+t7lJ7/WMDC0q2gy5dIVjLNRpU6RKmsrys2+GkZWh/MXoZpJHD5HtE55ONKhD
TDzbD0YPO1gruUGeh4kMsQvUnLHHmgOOjsXBvNcizJpCAusU7jA3bxxQcRmGgRoi26DEP3C9flzL
Q3U3jCPUp4RVel3gMvoyLkxle1r3wzEm0zYXTkOCmLAKK6QzewEA+vxeaCKWuEbnGzL0gy4yZz0s
xiIgKM70ZEpD6VF7OVVL+UreDhGspCTzbVsz6IqKpQPAX22lk7RDSzuSaGvHpt3VAVaI2jUQ5jzT
eixnanJKJ3HGJvoEIGUY2NAdKTo7WlEKATXcWR3hc6xp9ZzE/O9KkHD0KUjiMQAF1IVR7qYstRhL
Bq+EnwDbk/bJJCMmX2tbtdl3bMMunti8hQN/c3Xf2N0aUt2uBqZjPJ6cGON/uvUaJIyTf3cWfdF6
tXR7bWTgm13xOlllpHncVkGRKRgH1/+4wliVwgiR+AbzDo/GtRlYWUjQDrQ93INuMMw4lRww0k7z
hMqVYZrCd53YpxelMewSmiz7n/Dtu+sYxrQk3qe1FVoGOrsHoWWkNs9ukGN0+xEcjKhC6cUPxjP8
zbRUkSey4YmpGR028kYB/Oix5eEMAoJB7uKapm7RbpEGLdN3ZE0s5sulCwkuTeUDF3q6mWcyIKAs
1JZc3xVHGeS6LgFT4vjXActF8Gz4LC7k4Wg1+MKKHPkXGgB9lDPkRM9ecUakZmkLUxm1dOxFxdEq
EyWaMSx+j+xeA8+mtSFle5gm0s+h4sIBH5/hhNqhpZME0WmkVS1SGNGevgEKc3XMqWX1H3FRzweE
a6BhtxnH7X558d7/CmzGgehZ0j7ulDTAfHIRbdMbr3SlAgWxTHLe647IjJKhMOaAuFM8e40ljzHY
x5d1A3ryCwAA5GvsW0rYNuARkjBfT6HVv2G6U0cJxZJH6VfAZyOtf3ekH54NkpDsiWpT8mfJkunf
OsGXhX+8Owx0gaXZhBC6/YU7aHuomvDBlsPJX6l4MFnd2jUBo9WddGqleQT7iNh8KUmHvlPcBtnc
ybT6/oVMGbV9U/FyKmLjNC71xhojPxk1qRpS7ybnaesxwn8/u1ZBY5/TayXSop1H8w/pTqAuTKbB
JvNIKAxk2U0FUCMgiBIOqbA/9/oKOctC5HEc+lcOMe6F1TSmKJkRVvuRjjhMdW4x1sT/WWp39g+q
T4+dNdu3oHkpgF8HVaIxKQ8wJVjcvKw+2IUVbiqqvwr9FfwTRlydSXY3RfyahUX6+rlLuuKsajxA
kV0ydPiLwuBpAecp4Ii0UDIt7YI8JwWchV5e9xHGu00LNUHeSBPoxSGOyK7ved3mX4uTpgFwpp7z
kX5abhX/efgu/enjGyD42fHJIJBGU/dzbA5daarIHHjIcEKM4jZxu+mF+ogOlhw9PlKN6PPBhcqJ
g++DV15gvPD1Y8q+ODO0ekmA+Rsb0onXb//Q/7iCr6yXRrAPZspfgXmoMGFeB9NSKn8p9NeCITXj
8oTky87KhhTiiCWaSWeIpZWfmRkq1UdrT+QLYhCAoEnjNxVp7kEaHzygZP4CI1wkcxRt+Dc+YQCs
OL+n7HZG6u/0yEaMaeIXvTXxovd+Z2XJv2JIPuk/ab5JpNI7Irib4Kv4HW9CbCmUml4BHiupVKX/
0PLcuSTCPtxZGUOMUeNo5RT77TRepMnRgJ7Yf4NvrcJJJPep6vgEzobqF/xZjIr/ESvLP5b3pFwd
4WCMw0FuAcQMymYG41br1kHD5+zBqvYuaNfYkUa+pYvy20B0rE8KHxrsWFG757HdvE5+Far+PYxU
9qmqoPLFgB3mVWEyKIYsomRnyGUNm5ws++L0aZ1lVopDTq05Sa9Ib8XY3Ca0FcEUYNR6U/Hc10R+
t9YDdnnj6RMy7Nr12VAD1fLIh7BwB5F9ccfzCBiQTK/7HlHKpBVp6OuiVsXarfsDAdhDgFg1Z9WY
aIwgPuDk0uJk46ZXTuUFETCJRUZ9TsV6Js1sLCf/3uuZjJacH0yglrw7WOveVx0YX9fdkqE52NOz
kRQe6kssek3q8d+V27pSNebZ9l180Y6jAcNYknUfpwOk7HkUhOXsSEZ0BO2EmejA9CEv1iSgppg6
dScdNPPtSl0Vw1qIC19NYNZ9+gsJW7qAkwTxhNtj9cXt1krwzXDnnoBdnqKbHE2/YSTVqundm3fI
XoQjNq3INcq9TNBY2t8JSq6bktK960NJpJqca0D/1yJiNY8W+eHwjEEZrs6RgbH8A3HtwYU3jaFc
RyWhsMc4S9LQB0i4nUFU7drzMUg95T27yNl3h4zunQfk71dE+0CzCOJBdlnfRrR8R1MzRs1/2al9
8PJ1ZeC+oxnM9rqFNWTrnF3WDiw/ay3Omxvfe+2HF2i8R1lJS2YFXkrWnuk+yD+Ur1Z5+lSp630s
pmn5ApX9h4lA9Ux2w0Rx0HS01hkZ0xlT2AEM/1SBYgCdT/l+weW0nSVjGzAjQyyatJeF0v0uTAQS
dLMrefxZ+ptLnPsb8VHrIfkoxTOUYKaZItkJvt56U/O96tYQKE5xydAsrsfiz5SamWzdhVOFfuh/
q1NZ92ussO5MrB6TWtppZz7EpgW9qyVpGt+mrb77Yb29l2DMTVhSRSvBs0eMBYBBZpBn5QOUKOfq
C99ytvkc+B0/z0Tqy37T49lBWe9x1uv/evgZDkj2x6W1B+x9Eb8IFUDLQzzoA/tNP36tlBxULgIP
Ao7L6GpWe6IOklKaBwuXdI2eqNJXCSIR4iKa1qQyJ81a1NTFnEQSzNsdUR1vCUjprckMLosEKbBC
BUusWat83rceXY6ENt21xksdzDoP5GrkLJt4Emptim8cTrhh2TrYhelZX5PqSRwMO1jH71VjyBzB
a5ymt7QFTh1TliUHjkTlP9xMcF1i4XJHm0QNDKs7a+4HtDKBupjU7kCBSpIj9JMV3nkUH+WYOPIw
dkIQ2Cv+k2e9v8dQjZpjUmsVr3PmP9YgEIGuINAnJkd4H5rIbc7cRk66IO7Q4Sx38sHQXI9CiKYy
4tJWO81rvAIDAbI9hSt1y/Vwd2f+9Ib1ETpcQYHkacET+nu0GXWdzpxg7DPIZfZWJQXHdrlZRHnY
/2Vlq90JweYFXjeTOruLief9SO7//vTpMWwBHqaQVRwYw/tLsWgEUeNshgubPFtc1Rjs2nJL+nmF
13mzzxR9rgTA+XxMTQlJXDTjIz9MRBBurJqKKTZ8yh187MiPsI97tf4DrlJh3M/UFsvqqah6Of4z
vkc346yHmqw9xX6QqZbZkvEbtfxgVaUFIENajODUE5taQKS3G3fjFWbdWQVsa6ylynuevEmyoyHg
trx+zZo3VHEHY4zGDuwPV0/ySsrEHVf/MuTCFs13AVNCrYgmTyXQqOg5PdJsZGIFrrYP7FhBMrMS
dqlBNMqDj5IDKoOlPInj+qa47TcHd2r/62+E02XI8M4W5nHgzIe34V3S3jr01GX67dOQ2KReqaMV
vPmXWoCUaA5i3qgPEpfGXL0rNwodQLUUWhpRvrri5T4RXvkC/9GlAhVe4SUPzxhAl/QG12aCTB59
HCfma+glCuaiQds1RTqbaNhIVUawMzJTFY/RlOo7SndYDfCg3nsWW+xEbVTYxHV2QU4YowAeHyCq
jug9HyAklt/VrqbKax2JytqY1qe4BRl60gGt7A9BqNOI2UsTBMAjj+YyEZxwjXfGT9CaN4OGKCZ4
IFqruqgn/qBhbMaCdeMcyY9sOGhg0tw+ujkyT/i3TWehfck8VZhwwDRgQPpxBjSUjR44rfgxD7wd
eXj8qE48KCpm8eyJrgyMTm186+GPlhceewEuqitqwigNNcyJOT0qujwRNbCKIjehjr1ORWH5mz30
0/0uyoCSKlANs63cwzOjwzv+f6bhjvLMgI0Dsm3tmTRLr9y53mhCUihsopjilxeYH7G8TPbjetNF
lDto6B2P0FBHlVkjCyyig6BlHUrDpsqZojmY/kbWtsLfPhBJUbg0vIIDLgNHwinfnyljNWAU6sc+
7yXo1IR1DfPtMi7OKwBqkYWiTkR404QqtIUqNBjcQ5NCftaS3paUpGm/q1aSdTqNYbeVY1fDTS38
bJjHh3LMA5UvVkGcbiaP2FSTgPCpzZmQYkCBsOx/BhbDJTVdvoetu+ukXYgF8Yrg782R9cizbCTL
iUnyeaz291W97fK80w5B4Gia6N4mETSdkGUxlDln63/++JbjmQp5l6A9snpnwh0BJl8/r4KiEPOg
cGdx7g/usjRrKYEL0i//oWxujm24uCYMNsSUzOm7C/tpwvtrFVe+dOeZWGK42/PeeQKO5cjvZ9XY
C9TQEl1UigSbnNm81cG80na2hFfzmwS7x/fP/BaEslr3O0+9LWSJFjRvkJkEfZAjOUs1Y2I6XIRZ
u+N8CJbb+XqxkYRQbI5Cjc9Nouipb9xK5YvH4bOtCdJSAbiY4fAF2c9vJHIiWF0Xf1q73ZYjyCro
MJ4+5yyZMz3bPNvc+BmJw8hPdj13CheNZcIrKj5GGcS/Wmu9Nem/Mvj250prxjlQe3sAxMcVTqaC
P4/65ynSv9op2klISfQYdOhYLuqTzb/qKrwtrCZ6UmjRh+rid8r7Z7n149FikmpC09JzRDuD1ITO
aBnyyKLp5ORT3wRmIOCt0vWDnde3ao6aTGbZ/0myUmvqyVcxIRr/taQ3bk8Pb2OrljYzY2aB9nVi
NL7qlbV8ZRCYzbqMFQnLgig/t6HxLvptinoOFdkO2amn4cBBWDMEtOYnEzY+r2JbrLLRbB0B2FAU
R2w6PTdGGEdWGVaFs8rm/Li8EMXf1gLRclgH84LT82l+fdaCoV0zmTtdr+8aiD+WwXMNpenY8w3T
Q+8DyEnqIjl3T4JecmSilDsLCsNBmkczYf/cF+U6n9vjpQ2Aa6d9cVGdZUoXwuzREoyYrTlswEjc
nQwJZYZE2GaQd7qk5h64GZduu0pA32rABflu+3pbGN8Xr6g/VCpRkoc61K2DrUhGTP+T5WuEZ/OD
BeqF7S3vDhxKAJVFu5udlb4kOnsr2Ww5028ZviQz9pgIoBDWkYhvQHq28G4wz4rIrexqE5j0U+I8
ksX8ulfH6hGMhVY2aOPOmY7x1cwLzHMVKYmDlcdHb3avtPG2JEw4/ZgCPp682vEdcUjyDNFwrq1s
vMl6TmvcNtGwwsWm2VT+q2nEaUFJIFte3Dzwyz/HwS5xC797ggSLqh0zlp2EhOlTq8H6yu2YqASz
G/ECBtFp8aO/vmgMFN6627rec/DghixI1g+eIw41fLRj7mbdjmKDMk8FEon7JM2NnVD5Ljz+eG7v
LOEy5n2arPbZmh1X58dagw1NRKAkdFuvOWHsqIRY2vZHtodhEv+VAAlh983bbomOMpLcat+oqrt+
KUpboX9+jH0cJjsGRyQIjvdeZvaqKeVt2bbUvrcfcQteZG7eS063F8V+C0hL7qJedZfu++uFaqVT
sGkh+B4lzuoZJH9NKLwjTZSCol0NxWTyEHljkwwfLnZwknAoH9eY4T4gd6UouCFByVka2xWLAMB3
3KNwPsdIR8zmNZ3EvaHWnQoj3GAoZJdwJAUA5fumEs8jXsW3xoGM1f+QLUG3eomjkvhQG0jmuHLX
tJW4/fyOz9iWNOYpMwRVQLL/+XPTA/T1MlN6oa3gwOYQSk0fMYojxKwaF3NktDFNoPR7uHjaFHFj
pmsostOUU4s/1G+K1j9LRbZdf3MUQNkq1OiB9ywhCnY2eYMmFe+8FjIKwhz8NGpBh3iVZoe5nJzg
jHfrLRvOAyH61JzkCb4s01CXbGyGwA+xuDNHjedEq486jiQeWozZIFjaKui8TQ4H20zSebA3zYWU
OQ7WqH3GexH3RIjhrZTWPWwVNdCgzrQsA/HkmzRARqWX7oeqFH2YPwrOUTNCdIV6jPoi0S04dEOs
HyJkzeqY7R9kWAKy9btAYfwlRsohn+hLztHw7SvPZZlZlTn7XKLPx91OFHU2NfbF+0D9HWDShd6J
pG+9zv2oVCFKc6N9UsHmMxAHQJ1HxsxzxaZ5yOuxsrOh4ALJd2OPrVi7eQEOc6RsVvBjSiyWEhGn
uBL068vv4u4nzz9/PHjKvty12Xu+Mn7VxpjB9WpKT/s+zIIEVr36t7uOkL+Kxh8K11LYinteFiaD
eeFYaM5YFeIOCEqgnTXpbqLAwynm1xmxrpdqsqqr9DMEuFUDX3XL4ghyp8Ws4ur9V64hihmWfAud
SAaiP+0l+FHFI7/sTTQsMCTBzP2G6OLJNK1LkiOBeWhcyGan1eRpn+tKzmTlbsR+drJt5DRJn7s+
2q5L3ACOAdy/6zPkpMvW0iCl0eF7ktF93uLLOox97HfjsUL3fcgjZmMBClK32WzhVzBpn/feH3EK
PGvqCZiQuXCpnEICpf9omfS5DmT1+t+jU3EBSEP2ae/UPsMSWcgu3NuN9AyLLlgfio+4+RaeqMWj
xFtInUo0/ancgXrRRhChDjrwy490IaLgAFy0SaSxh4EGNs94eDKXSmG48sJvUSJ+xLyoYlBGzmHU
lJuU/UtX+vZDD8forzVi01p8VWCv+D4rkBB9AlEMrIaQHOOqKos4Q5ESejp277FU8z+gpjeSRHaV
gu3qiqLj1n02Zi4ycP30fc+5ljb1u4VLndQGoUza55TuMLnltRzrI3eDqK0QMrvOsUa6YIgh3Az+
ifpRYNHOibdixCgxXsyoeE2RLXD78qB0ekkzGT6fWaAObYYXhp2a6eZob2dJV6QxPcMxU/bIBLfn
WmjnJLPGYmpaUg/EuBlDQZzH27xGkv++ziJvohSjnpgknH4SazfpWMwPqIYLdr7Co0gUjzif+6rv
cHJeeBgSdJH/XqVqmaOKCuf/E1hdNJ2qHhQ/4eJwnkhYczI+t4iwMjNVg8eOw4kj4RAYUYSq/T5B
K0S/7mInXB7jiGPv7yu7xYe92NYTGj9K0MU/VLw5umTWWI4ZBh0smCZ9NnLppLPSmVkrU741pzJm
3U8q6x7PSorMs2vAea1GCX+Ekubl4Z2bO8NdYaEGy9IzFgXEESx2myRF3yQSohxdFh1nJlnKwr7u
L0J5jXmGWbIpEH3c52RD6RUv572p+jGNolVwesvXBpQWRrZ1r7VplDNBdEJ3BxXKlhZfU1xaN2QR
ebuPrQCn5xkCK/ijaPw8/Cq5uHf6ayCV/JFS9ooSyLtBfcMzbaIiOHPXXw1J3cVFsAPq6j8hE2zd
6kF7eZg5+kf+hWamrDjb2A/hKSswcet2Zjf1X0a0MUMpabW47kPSwrxUmo97Rh2huAILIgC1WG0G
bBsTPDpixPlpXjC7JLpQm45pt6DMLKWASQImwBlWwZ6LCID7ERYny0oAY4ZQu3LPRyctLdbb4gGt
f0IqQLf5n1HmEGRuJfObwaOsxAHOom7AC3NSpqrXlWi0antdZtTgOE1GhV6ZF4HI5vBF0Iw8n9ka
hVcSEHqWyw8njusC3hQzMybFCdDNB0LkifONr8QZZpbjiXZwYry6gdLMmm6bTGIz8qYbPDDgTARH
j2803TZfc/Ino6/xoW2m+N4WPNl0gO3SJ4Z4ebNFHjcqCCj7+HF6SJLVyX4cX/TQ4cCwoQT4LWwY
cSm8HkwiyOmCFoz5oe05zogMBVCgrdMlqVgaEFPl2OR0k6eRL51cwzLeShd6W5VoUSLqkDI6qdV/
ZBDhkfAUnP5VeG6Idlc/vMJxgYQ6kSv5TDh7+VGmB3AYoesFuGH9iT6/iGsvVRj/vyogw9Y0l+CH
2lHF91S8cK5zbTEJzCmXk2hQ2GBubjvETgMhUuhdA9eIci5SCfTF5HlqiGgx8barf5VduUlHPG+m
6TfoVSE0HwOZdHxNOF6rkiJflqlQOkckNhUG5mlk5SRo/A0gA/WhC/TPTQc0+8x8ObW1UdjgG/k2
DfkEKtaROFFNX6mOWa/nJc0pfzQvUdDRttK9HEnrReBVTHD9LW0lRJjX9DKReqpZMBIf7Rd0pRhB
3WM8fGwSn6IT2qnYcmSh9SLt0Fh6xvIXOL/imqY6Tz1UK92dyj1G8oi3aqfJC9c393M9Hs2WJZZS
wTB4NsXj/FtZUvCI7EKvzA82FLHQyIJgJ5T0NSV7v0KndPR4mXUjB+Hk1yfdlXYlAcJ6YWOmEce/
OBfAuIwTJQ5n75us0FjbMj/GbZ+Il41P+nZ/h0NYadRIcy3iuXtCq4O1lA2dCxhmLXv2l6i8gr6u
iu8N9LFein8CTc9JzRdM3qFxUu35CTprYR4VqNVT1CYAFGc53QYb/Vh6Eukri5/L2PV6Q6pcX27C
GUFN7qhkE4ByqwadVTQECAQg1Vr9h6ADK1zK6v2hBtqwLLC7EzqIfc6MAYjlVW2RqlvwoeUQ72Co
vHITww/tH6mR2fIvAdnM+wQK93wu40vThLimZqUrdRLEojH3HhyK/pHCld40PM0WEjt4WLLcNwct
JoUU5JdI/3xcaaPXIcFimWUSih+0KVTHMu0G3azV5kL9CRW4HojfOuspILOqnGIJgHYV11r6gzdb
52V5w6GvnvHhWkpfvMJW70NjRER2vFEuDdLzz42arnGsogzRuEgvhXaFoY+UpjT2wYszgXTzwvpr
+EbJO2mbi0ZHskTLA70gj/XVuqvieaY+YxDTgvvFJtolRgWCiyv7sPMRSQ01pcguV6KohivL+mpQ
R+ZYmtVEk9BtOhQWEKCOoBrJtDz2prPckyHgSHZxKDXOHFn/NvRsjHWdD6vpWbGrWCI7cALNGpz/
eaw/epD7VMim4hngEFL/AYw8bqzWnlObwOgQizylqAF6nPDSdAUMjXCWIRAYtB75RO/RBhtjfIDa
5/KJJtDH9Z8l+2XUOrTY5mIJRn2QsiEaKolQxxskMZq3SjfxlndZdeo3n/8BuZJ+t42I7ylJ+tWY
hldCeW+n28g3yCizGn5kQYa/a9/y/KmSEA/y1AtbTTRYSwKmExMAZmKJiMDZGEgxP8jPzx8or7E1
sWcXzKAQ4WJqPOv6BV8nOVAQm7pi5VUnDsOVNKEvFpETYztIxuq17s83Dq/ggwplnu2GbKXxBzeg
THgS5ZAf3r36CwlKBi8n9kLvIxNNaMfZcHwJFzovL5ssbJtZVwtF4SqRy3w/QSRRFAQWpL55GUQg
StSrr217JyVQ3ywnZrNjzOGQIVh7t6QabrWhO8VWPei7NT3PPjr9Pwz3rDzmTyk8XvDe+ahBWU40
oLVW7zid5vx1E+Ca71PpIEw+SxpYhXTmzMPMM7kXAZZkJrLEpYY+jIiD05cBldtGPVuBINQgE653
1mFWwp9vhMezWGKj77tZ7D+avglpzeoOQ8uVlsa1hiCbSvj7/DtTlOHaZZYUpnho2pdV6cOn5SRX
5er986yeN9F8mOTMyhbBu0bub9xmO6PHl4emZZekwe/CIza3oKB3zat7nZmS6dCWalHYpuQ8B3oC
zIaJheGcuGB0nSD6jwHnYWqGQmwXSwFWZ7xPr+t0OCzBXiV8eFusv73jiLx5HmkfcHXLcpeW1uHR
izYJJgliSOE8kfcxA9Phtjpnd8CiD0N20GfhVfczCpdM5z5dF7NPMhPg0fJ8hgErPg2DqZ7Tuqu7
PFK/Lqn/jpidVprPavN4rOyCqhUi9Da5BqfK/fcV3DHMOmz0rb/J1+Q1OMiR0RWQ+Cj2oCDqDLfm
BTwJYprMobYbBNk9ubVAcZrgFbcAKcqJosdNsDXHDUGaHq3yzUKJ+arELYhXO7jOAbE4Nx0fmisT
13Ww9hkHpD/YbRCrtF/4xUwVqOVmlNKggqlXEL/FPx9IzZ+IY0+/+NmiN36MTSYVW04WVqdv4bl8
PgSGUbSFu/bjqTf2+zyp2mS3FfDqjMLT0Y670+L9q/daMH3q19qnKbu7GJs37Ca3RUEY4wIdLwk1
W+DiJ3I3X6O8AvQgyLw68A14Avgu0Flv3S26ySxPAK+PIMD6VRYChwd+6tGfTTTK94smew91SJbP
9SXtUIU9vC9KjFTJTyu1KIaJrB+I8pB0oieb/SS6qeizCgJYldvnFRLytiXOyJ7fy1uvNxz90yAF
4CQ2qkoSpnhDEUGsvSXNoGhzNJTTub+H/7fa1nPsoWJOB7PLvMzFjWgQt2ELy/Y9g5tz84QOTYMG
1Aqa+DxTIkfoU+4LMhSMZruOvZCG6GUsIZAmOgxryjb11CQX8VTzCJRuZqQyBCKB3nDVXgTBAxfp
whJN6xW8WoCCa5TyUaTH/2jf/k26TF+wNhOhQue14VIkutlCZF3vYGwAW3LKoVJbvSLcP/1ZEuyO
Jhsjkw4MRKU+9eWROLuofOtYPX0UxAFIj89e0gIqINofREATf/ZboVNVanKGWsIUOkpcTBJU73Ir
p9ZCNjlkFCpjLbArRCalGA9dUzTIqWW0AkP6Q8S7RjkNDvRmmlQP3asa/Ufsy0Qhi4vMoByhUfI7
kCU1qZMEsZ6kKLrzgpiR9//2yH1ilQfoK0RnV5NTMUHUMNYdrNrBYrcRuxk6Oow9tRS+js6h//wB
xVL0rI2P/1/9aXm4nN6DxtJ4bD/q4xKZc0JyguziQeMlp3jIxfhzYs6BIQtPx07I2Vmi/X0t/n/p
1jtjzB70BAW/Z9VVnuPkzUyMTyXnLZDq9TN/WOihtnOMaI3iIurcEIbCGt1wYhELpCLWOJaH7KXn
x80p1Uee7NmC0zuWQa0HDKLUBVnUxJSOyBj408ycOvY98h/ChDd1Te+uIqYDqQSmMDqSiYi1fvij
0kvKM2uMk2A2U2jqCvctPeEnqEV6v4XrJSKo9mnIWvi1nO30cj+USc2JOqpOkD100uNwKw7k4TCB
FncDWx9nXytAvccBF6PIGKsNTcgT/2CffOYBM9011jFP0g2WLB7/tiS4miwuPTBoo3RIy1BpJW0x
z49vtAb0wrBWaD9F8KopOBzBT3OTNU3vPpbMCOcbXudO1tJjkTkhlorHN08BHjWklKW5rEW8Nujx
SyUM/PFK9Ak3WJV42LjZnLmuNOVHidnqZKbSPz5YPsMRsM62ayEOcQ1mTTkqOFZdhaRjKdnlnl/Y
zzxrvHPXR+ZdBJ+v+s7p064PE9ScoxdgfGaFE0eEvSowb2AioVrWbp/EMEI1YptnKU917+rzRq86
vvcxqeOmzWMMNPOVy5lftV2XlmQpA+oleV9raVWtsYoSVKkkf+nayMMuatsKtiIIMh8AbI8/vd2f
BbevHcbHRbJDyk/tV23tASWRmDqHX/cWalZtyzXflUuiWLA/d+MIhGNqBdW2yKugiir7jUM3Gh9Q
Zs0Evkfnp2xRANOkRJZ8m5R0o9GkcjMcRfR8YplrBOkhhcxbT/9Yc5ss/V3eqUddR/oxwpexG5gh
bO40LbTJBOFqmGzKJeuFzTqMCoXXVjlIJMyK5HFHX8l0vc64UWlMG8w9oaMolg4uSB93UaMNEVzb
3L5u6yHdUIYR0rQYGCp/bv6SkqUsLmHFm6mjU1gYxwuWJaOThOzG7iNzSWZ9Ym9G0GXOFpaFI954
9EKsC5qygPNGeHVj6pkS/pVlTtlkPK2JIcihfmZl25bhuLzscQzkb7SZTllG1YCNlrinfGam/q2T
x7a2nVdbvb/Ci3U/+CE7+M+A+gj4mzoDWclePfzy3n9CiUnViBiPvTMkjAX0UosGwqrG+Lb1NJOp
Pz5BQoc09+kI9ZywX1FwlHbwEZC4K5BjcbhiE2GbYOWvunkX5LtGNJZ0zHe7lCSPuKPvrMm796dY
zdfNakPn1k3+EvIEuZ0ckSkNFu8vboYylZsh+KEiCcqUuqaWmua7TOPcoG1RAs8pp02xsC7qSdrz
WGml/V2jpvN5Ts01fVXGIpEx/KIVppK1r5G7nX6B39pMz6hsfndrmAv7v8wgFgkdcoHMP6AHqlRt
ncAQrKhm+vL1OWMsZrtEaiM+UmYGVs8gnM/JwV7024dVNtIqVc0x+Tgl2MpdR2ZVm2QXR69nnpV6
8rzN2DvW9HK7Ttt1FWI4syS2uDhuczFf+NOs6awgwajpsWIv083j7Mm6+wl6eiyitz6i3oWA67tO
gaK2JN/4JcDEteTDtxa7JeNrnepTpkUEO+khGuhj1RiLsLz+oIlqRgAZiD20u1ZgyQQvxcZbTv1m
5tt3LgL8txfJNcZfZ2vmHtVazt0NmiUJzI+xLFGkGyyn4KIC1GPzck54TpB2Az/+hZaLxvrJlX/O
GWy9Q3qdUScZD0EVyW+Q6E7aUOIXYG9TGxSuXKfWJOA6e7UYnqCIIljqtePwJwJUB6lHSrPuSGMX
T7mfUEZ3AOGk9ODW0LG1U4WjulUKUZV5pN/nkgj92YJUwkJQz7x+BjW88wOuJVT4zTny48W73FWW
BlH6wRsQlSbTS4OCZsJEoRr2zEGceY08Nr7y2SRu7P2wl4jtaJvKbuP88eZgX79Yvwe9n5QdTJQg
0OVE6CfdQMt+znm+11s6E0/5ProF0C1ESOJz846io+wL1mCfMuCd8ItxUAn8LoGZ889mhzWZ2PdI
E34Zv8qWEViPGzFk/PU078pSp/LrBCc5+vg3xwZe/i51uHcYcyh8zNhlOCVcyOrRdUL+6gnkfusL
Seutbhhc7bU/a+4ZxEfSkDv9K3p1kZ0y67wl5Sn9FmKi6PViwSuaSaHqa6frl/lEha9wnB/DN6G/
FhVFvfC5UgVqT2hTdFlseIUlthgm0vaUlquD/vqa47VoLz5vGJvQ9o21O6DOGWZlPt6NkO1OKUP4
HV9yNZe3rCqqYiGoGQWJRs8S0jZULfDAPMof0p4x9x20mYZ2z6ni2gYTV0A9hcI2X8QLiznDEPPP
GhAbHM+3UpeiQQPo9PX3H3IuAqtB+KbdyvHRNyXHe7AyYvFva2aAUBDhI0BaIAfqxlUILy63GUyD
k0HF3tDHWJAb6mpl4DzH7J9taa9NBUPVuCq4BlESpR515HO1XwGdXR/+NiCi1U7rj0nt9HluBJrX
9sptMSg1zm63itWPIn1j6CrGZXZgt1GMBIa9PeMF0Ld5kHcGhUN/PBosoiVroX2IfKwyjym71Q0D
zgioYXuoEPWo3Roou8vqSjSzla9p3W2Jhw55ZrvkePrVNyYVPBPtkWtYkvSdeeuzcZzl9xw/YPN1
vgdoVwsHBTV+AQTXmmyX/XuzimcR+LmGR187RwB1gMeUxtOzPojf/9gAsitCxfpO3Pru7xHZWYcS
QViX1HLFNmH12xVtrJKEFqse6zrPosoIzMX0S7/dCjVlBtSEfvJvzHCF9p6AwksAAM7zGFcyIb31
E+49lVGLHW9wkTeQBL8q2z0qYY9aFgMhbSDK69GJWMeCoDWA2VQ9Afrhlf5rwPA0UyLbV0jWmE1Z
F92dZUfkZX/6/vEGFmffwlh5CnKYyxkcDMQ4lEB6lLRxZqX7T9v2QjNbPF8oPPyA8SAW6q+9d0Ao
z93zWrfxZtgjEWBV/kGVZXeiwDdZXxrY2dCg6/c2RHfgtXYF5tOzjEEcqAa9/cE9j7s35flvd6oz
RGKUs1yPdZpTPb2b+5StWzYiEbBxRo62pFjqTdqUmCHOjqp+q/1jv1ZBfhwmk1kqsdhUgYx67lhc
5snI0QNr1whZ0krd5iwD6iM3dfqhsSIRnZGtw9jrDRnBhAllIXQpjnNAImSQLRbhcmY4UHr5lwI6
qY7ugkHKTPY5AvwAFrwzTxSKTwWrq95Ja8qDFKLbARQnEunytyzxnc6gDRhbgbEZKHkJRGDVU9P5
JoaVaiyPljuWRRGX0VTqksM+0ZaidGZ9jrwb36x1JYMkzo3o1ekWuRJRfPkwr9O0sIHRSTTb1IVr
lwAv5Kf3DFedF7Sfzor9TlZrcAvqzApq39dgqPCeH9sUTHyCey4APItoqxm8vlYkjKgo3uMdICr6
jfTkHpsGUw==
`protect end_protected

